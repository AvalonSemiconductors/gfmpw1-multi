* NGSPICE file created from multiplexer.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt multiplexer ay8913_do[0] ay8913_do[10] ay8913_do[11] ay8913_do[12] ay8913_do[13]
+ ay8913_do[14] ay8913_do[15] ay8913_do[16] ay8913_do[17] ay8913_do[18] ay8913_do[19]
+ ay8913_do[1] ay8913_do[20] ay8913_do[21] ay8913_do[22] ay8913_do[23] ay8913_do[24]
+ ay8913_do[25] ay8913_do[26] ay8913_do[27] ay8913_do[2] ay8913_do[3] ay8913_do[4]
+ ay8913_do[5] ay8913_do[6] ay8913_do[7] ay8913_do[8] ay8913_do[9] blinker_do[0] blinker_do[1]
+ blinker_do[2] custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] hellorld_do io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[10] io_oeb[11]
+ io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[30] io_out[31]
+ io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] mc14500_do[0] mc14500_do[10] mc14500_do[11] mc14500_do[12]
+ mc14500_do[13] mc14500_do[14] mc14500_do[15] mc14500_do[16] mc14500_do[17] mc14500_do[18]
+ mc14500_do[19] mc14500_do[1] mc14500_do[20] mc14500_do[21] mc14500_do[22] mc14500_do[23]
+ mc14500_do[24] mc14500_do[25] mc14500_do[26] mc14500_do[27] mc14500_do[28] mc14500_do[29]
+ mc14500_do[2] mc14500_do[30] mc14500_do[3] mc14500_do[4] mc14500_do[5] mc14500_do[6]
+ mc14500_do[7] mc14500_do[8] mc14500_do[9] mc14500_sram_addr[0] mc14500_sram_addr[1]
+ mc14500_sram_addr[2] mc14500_sram_addr[3] mc14500_sram_addr[4] mc14500_sram_addr[5]
+ mc14500_sram_gwe mc14500_sram_in[0] mc14500_sram_in[1] mc14500_sram_in[2] mc14500_sram_in[3]
+ mc14500_sram_in[4] mc14500_sram_in[5] mc14500_sram_in[6] mc14500_sram_in[7] qcpu_do[0]
+ qcpu_do[10] qcpu_do[11] qcpu_do[12] qcpu_do[13] qcpu_do[14] qcpu_do[15] qcpu_do[16]
+ qcpu_do[17] qcpu_do[18] qcpu_do[19] qcpu_do[1] qcpu_do[20] qcpu_do[21] qcpu_do[22]
+ qcpu_do[23] qcpu_do[24] qcpu_do[25] qcpu_do[26] qcpu_do[27] qcpu_do[28] qcpu_do[29]
+ qcpu_do[2] qcpu_do[30] qcpu_do[31] qcpu_do[32] qcpu_do[3] qcpu_do[4] qcpu_do[5]
+ qcpu_do[6] qcpu_do[7] qcpu_do[8] qcpu_do[9] qcpu_oeb[0] qcpu_oeb[10] qcpu_oeb[11]
+ qcpu_oeb[12] qcpu_oeb[13] qcpu_oeb[14] qcpu_oeb[15] qcpu_oeb[16] qcpu_oeb[17] qcpu_oeb[18]
+ qcpu_oeb[19] qcpu_oeb[1] qcpu_oeb[20] qcpu_oeb[21] qcpu_oeb[22] qcpu_oeb[23] qcpu_oeb[24]
+ qcpu_oeb[25] qcpu_oeb[26] qcpu_oeb[27] qcpu_oeb[28] qcpu_oeb[29] qcpu_oeb[2] qcpu_oeb[30]
+ qcpu_oeb[31] qcpu_oeb[32] qcpu_oeb[3] qcpu_oeb[4] qcpu_oeb[5] qcpu_oeb[6] qcpu_oeb[7]
+ qcpu_oeb[8] qcpu_oeb[9] qcpu_sram_addr[0] qcpu_sram_addr[1] qcpu_sram_addr[2] qcpu_sram_addr[3]
+ qcpu_sram_addr[4] qcpu_sram_addr[5] qcpu_sram_gwe qcpu_sram_in[0] qcpu_sram_in[1]
+ qcpu_sram_in[2] qcpu_sram_in[3] qcpu_sram_in[4] qcpu_sram_in[5] qcpu_sram_in[6]
+ qcpu_sram_in[7] qcpu_sram_out[0] qcpu_sram_out[1] qcpu_sram_out[2] qcpu_sram_out[3]
+ qcpu_sram_out[4] qcpu_sram_out[5] qcpu_sram_out[6] qcpu_sram_out[7] rst_ay8913 rst_blinker
+ rst_hellorld rst_mc14500 rst_qcpu rst_sid rst_sn76489 sid_do[0] sid_do[10] sid_do[11]
+ sid_do[12] sid_do[13] sid_do[14] sid_do[15] sid_do[16] sid_do[17] sid_do[18] sid_do[19]
+ sid_do[1] sid_do[20] sid_do[2] sid_do[3] sid_do[4] sid_do[5] sid_do[6] sid_do[7]
+ sid_do[8] sid_do[9] sid_oeb sn76489_do[0] sn76489_do[10] sn76489_do[11] sn76489_do[12]
+ sn76489_do[13] sn76489_do[14] sn76489_do[15] sn76489_do[16] sn76489_do[17] sn76489_do[18]
+ sn76489_do[19] sn76489_do[1] sn76489_do[20] sn76489_do[21] sn76489_do[22] sn76489_do[23]
+ sn76489_do[24] sn76489_do[25] sn76489_do[26] sn76489_do[27] sn76489_do[2] sn76489_do[3]
+ sn76489_do[4] sn76489_do[5] sn76489_do[6] sn76489_do[7] sn76489_do[8] sn76489_do[9]
+ vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_stb_i wbs_we_i io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[1] io_oeb[0] irq[2]
+ irq[1] irq[0] io_out[4]
XANTENNA__3140__A1 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3155_ net264 _2604_ _2605_ _2606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3086_ _2541_ _2544_ _2545_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4640__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input108_I qcpu_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3988_ dffram.data\[60\]\[2\] dffram.data\[61\]\[2\] _0868_ _0935_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5727_ _2194_ _2230_ _2232_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input73_I mc14500_sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5658_ dffram.data\[41\]\[2\] _2183_ _2186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5589_ dffram.data\[43\]\[2\] _2136_ _2141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4609_ _1476_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5932__C _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5504__I _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__A1 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__B2 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output327_I net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3024__I _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5959__A1 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4056__S _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4234__I1 dffram.data\[39\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4698__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_60_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4870__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _1685_ _1715_ _1719_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3911_ dffram.data\[12\]\[1\] dffram.data\[13\]\[1\] _0740_ _0859_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4891_ _1665_ _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6630_ _0587_ clknet_leaf_45_wb_clk_i dffram.data\[60\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3842_ _0770_ _0788_ _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_74_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6561_ _0518_ clknet_leaf_152_wb_clk_i wb_counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_17_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3773_ _0718_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5512_ _1508_ _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3728__A3 design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ _0449_ clknet_leaf_144_wb_clk_i net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5443_ _2034_ _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4689__A1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput401 net401 wbs_dat_o[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ dffram.data\[47\]\[5\] _1993_ _1995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4325_ _1255_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4256_ _1188_ _1197_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4187_ dffram.data\[44\]\[5\] dffram.data\[45\]\[5\] _1022_ _1131_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3207_ _2555_ _2650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3138_ _2578_ _2591_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3069_ _2502_ _2528_ _2529_ _2530_ _2531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_93_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_35_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_137_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output277_I net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3742__I3 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4852__A1 _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A2 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold81_I wbs_dat_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__B _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A2 _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__I0 _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _1034_ _1041_ _1047_ _1054_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5090_ _1803_ _1804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4041_ _0981_ _0982_ _0984_ _0985_ _0854_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_88_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5992_ _2414_ _2416_ _2408_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _1701_ _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6613_ _0570_ clknet_leaf_1_wb_clk_i dffram.data\[32\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4874_ _1627_ _1657_ _1661_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3825_ _0707_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5020__A1 _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ _0702_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6544_ _0501_ clknet_leaf_131_wb_clk_i net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6475_ _0432_ clknet_leaf_61_wb_clk_i dffram.data\[62\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3687_ _0622_ _0619_ _0633_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5426_ _2013_ _2027_ _2030_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input175_I sid_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _1484_ _1080_ _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput275 net275 custom_settings[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput264 net264 custom_settings[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput286 net286 custom_settings[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4308_ _1248_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5288_ dffram.data\[48\]\[0\] _1937_ _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput297 net297 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4239_ dffram.data\[44\]\[6\] dffram.data\[45\]\[6\] _1022_ _1182_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input36_I mc14500_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__C2 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__I _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__A1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3212__I _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5250__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3610_ _2942_ _2949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ _1441_ _1460_ _1461_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3541_ dffram.data\[32\]\[4\] _2903_ _2904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3472_ dffram.data\[35\]\[5\] _2856_ _2858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6260_ _0217_ clknet_leaf_126_wb_clk_i dffram.data\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3316__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5211_ _1821_ _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6191_ _0148_ clknet_leaf_163_wb_clk_i dffram.data\[25\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5142_ dffram.data\[52\]\[6\] _1839_ _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5069__A1 dffram.data\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5073_ dffram.data\[39\]\[2\] _1790_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4024_ _0823_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2390_ _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4926_ _1564_ _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _1650_ _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3993__S _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3808_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4788_ dffram.data\[63\]\[3\] _1599_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6527_ _0484_ clknet_leaf_141_wb_clk_i net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3555__A1 _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3739_ _0687_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _0415_ clknet_leaf_63_wb_clk_i dffram.data\[38\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _0346_ clknet_leaf_88_wb_clk_i dffram.data\[41\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5409_ _1648_ _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_50_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_117_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4440__C1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5535__A2 _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3546__A1 _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3936__I3 _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__I _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5422__I _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3077__A3 _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _2210_ _2249_ _2252_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ dffram.data\[11\]\[4\] _2208_ _2209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4711_ _1458_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _1474_ _1497_ _1501_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4573_ net234 _1312_ _0642_ net154 _0645_ net73 _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XTAP_TAPCELL_ROW_96_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6312_ _0269_ clknet_leaf_105_wb_clk_i dffram.data\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3524_ dffram.data\[33\]\[6\] _2890_ _2893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3455_ _2335_ _2841_ _2846_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6243_ _0200_ clknet_leaf_125_wb_clk_i dffram.data\[50\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4498__C1 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3386_ _2793_ _2796_ _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6174_ _0131_ clknet_leaf_157_wb_clk_i dffram.data\[53\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5125_ _1830_ _1700_ _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_127_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input138_I qcpu_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _1775_ _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4007_ _0774_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3787__I _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5958_ _2390_ _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4909_ _1547_ _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5889_ _2337_ _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__A1 _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4489__C1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold41 net500 net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold30 net498 net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_max_cap403_I _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold74 wbs_dat_i[10] net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold52 _2456_ net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A2 _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold96 wbs_dat_i[0] net514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold85 wbs_dat_i[28] net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_129_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5205__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6022__B _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3240_ net278 _2672_ _2673_ _2678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5692__A1 _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3171_ _2571_ _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_109_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5812_ dffram.data\[15\]\[6\] _2285_ _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _2214_ _2236_ _2241_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _1956_ _2195_ _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ _1490_ _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4556_ _1430_ _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3507_ _2847_ _2167_ _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_40_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ net187 _1381_ _1375_ net38 _1376_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3438_ dffram.data\[36\]\[0\] _2836_ _2837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6226_ _0183_ clknet_leaf_124_wb_clk_i dffram.data\[51\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input255_I wbs_stb_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3369_ wb_counter\[18\] wb_counter\[19\] wb_counter\[20\] _2767_ _2782_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6157_ _0114_ clknet_leaf_174_wb_clk_i dffram.data\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _1803_ _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6088_ _0045_ clknet_leaf_38_wb_clk_i dffram.data\[37\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5039_ dffram.data\[49\]\[5\] _1770_ _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5910__A2 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput120 qcpu_oeb[16] net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_132_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_132_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_133_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput153 qcpu_sram_in[0] net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput131 qcpu_oeb[26] net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput142 qcpu_oeb[6] net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5426__A1 _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput164 sid_do[12] net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput175 sid_do[3] net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput186 sn76489_do[12] net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput197 sn76489_do[22] net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_19_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4088__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _0650_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_93_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5147__I _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_172_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ dffram.data\[20\]\[2\] _2001_ _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4341_ net145 _1272_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4986__I _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4272_ dffram.data\[8\]\[7\] dffram.data\[9\]\[7\] _0827_ _1214_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5665__A1 _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6011_ _2428_ _2429_ _2430_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3223_ _2481_ _2663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3154_ _2556_ _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5610__I _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3691__A3 design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3085_ net400 net470 _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3818__I2 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3987_ dffram.data\[58\]\[2\] dffram.data\[59\]\[2\] _0757_ _0934_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5726_ dffram.data\[40\]\[0\] _2231_ _2232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4162__S _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_99_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5657_ _2138_ _2182_ _2185_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input66_I mc14500_sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5588_ _2070_ _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4608_ net252 _1311_ _0641_ net160 _0644_ net79 _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_4539_ net52 _1414_ _1357_ net19 _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6209_ _0166_ clknet_leaf_167_wb_clk_i dffram.data\[24\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5408__A1 _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5895__A1 _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4698__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3910_ dffram.data\[10\]\[1\] dffram.data\[11\]\[1\] _0737_ _0858_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _1665_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3772_ _0719_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6560_ _0517_ clknet_leaf_152_wb_clk_i wb_counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5511_ _2088_ _2078_ _2089_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3728__A4 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4138__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6491_ _0448_ clknet_leaf_145_wb_clk_i net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5442_ _2007_ _2035_ _2040_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput402 net402 wbs_dat_o[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5605__I _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ _1945_ _1992_ _1994_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4324_ _1256_ _1261_ net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_50_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5638__A1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4255_ _1190_ _1191_ _1193_ _1195_ _1196_ _0714_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4186_ dffram.data\[42\]\[5\] dffram.data\[43\]\[5\] _0954_ _1130_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3206_ _2581_ _2649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4157__S _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3137_ net375 _2587_ _2579_ _2590_ _2591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_2_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input120_I qcpu_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input218_I wbs_adr_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3068_ _2506_ wb_counter\[5\] _2488_ _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3795__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5709_ dffram.data\[16\]\[2\] _2218_ _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A1 _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5515__I _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4152__I1 _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5801__A1 _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4368__A1 _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold74_I wbs_dat_i[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3966__I1 _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3040__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__A1 _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_75_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4040_ _0689_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5991_ net231 _2415_ _2416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4942_ _1701_ _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_119_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6612_ _0569_ clknet_leaf_30_wb_clk_i dffram.data\[33\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4873_ dffram.data\[56\]\[6\] _1658_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3824_ dffram.data\[48\]\[0\] dffram.data\[49\]\[0\] _0772_ _0773_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3755_ dffram.data\[16\]\[0\] dffram.data\[17\]\[0\] _0703_ _0704_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6543_ _0500_ clknet_leaf_130_wb_clk_i net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6474_ _0431_ clknet_leaf_24_wb_clk_i dffram.data\[62\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3686_ design_select\[4\] design_select\[3\] _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_132_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5859__A1 _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5425_ dffram.data\[0\]\[5\] _2028_ _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4531__A1 _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ _1953_ _1977_ _1982_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input168_I sid_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput276 net276 custom_settings[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput265 net265 custom_settings[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4307_ _0685_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5287_ _1935_ _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput287 net287 custom_settings[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput298 net298 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4134__I1 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ dffram.data\[42\]\[6\] dffram.data\[43\]\[6\] _0775_ _1181_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input29_I blinker_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ dffram.data\[60\]\[5\] dffram.data\[61\]\[5\] _0737_ _1113_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_143_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4598__B2 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4598__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__I _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4522__A1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4522__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3089__A1 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4589__A1 dffram.data\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3013__A1 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4260__S _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3540_ _2895_ _2903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_54_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3471_ _2327_ _2855_ _2857_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5210_ _1884_ _1885_ _1887_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4513__A1 _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _0147_ clknet_leaf_156_wb_clk_i dffram.data\[25\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5141_ _1822_ _1838_ _1841_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5072_ _1746_ _1789_ _1792_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4023_ _0963_ _0965_ _0966_ _0967_ _0968_ _0837_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_95_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ net261 _2400_ _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _1695_ _1690_ _1696_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ _1647_ _1649_ _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _0664_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__S _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4787_ _1548_ _1598_ _1602_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6526_ _0483_ clknet_leaf_141_wb_clk_i net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3738_ _0684_ _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _0414_ clknet_leaf_61_wb_clk_i dffram.data\[38\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3669_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6388_ _0345_ clknet_leaf_97_wb_clk_i dffram.data\[41\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5408_ _2017_ _2010_ _2018_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4504__B2 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5339_ dffram.data\[21\]\[0\] _1972_ _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4409__I _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output302_I net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_157_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_157_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4440__C2 _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__I _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5703__I _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3223__I _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5690_ _2196_ _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ _1548_ _1541_ _1549_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__A1 _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ dffram.data\[31\]\[6\] _1498_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_62_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4572_ _1441_ _1444_ _1446_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6311_ _0268_ clknet_leaf_128_wb_clk_i dffram.data\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3523_ _2876_ _2889_ _2892_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3454_ dffram.data\[36\]\[7\] _2842_ _2846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ _0199_ clknet_leaf_124_wb_clk_i dffram.data\[50\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3385_ wb_counter\[22\] _2788_ _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6173_ _0130_ clknet_leaf_157_wb_clk_i dffram.data\[53\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5124_ _1663_ _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_127_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5055_ _1750_ _1776_ _1781_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4006_ dffram.data\[40\]\[2\] dffram.data\[41\]\[2\] _0807_ _0953_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3473__A1 _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input200_I sn76489_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4273__I0 dffram.data\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5957_ _2359_ _2390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3225__A1 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_80_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4908_ _1683_ _1680_ _1684_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5888_ _2337_ _2338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input96_I qcpu_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ dffram.data\[57\]\[2\] _1636_ _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3528__A2 _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6509_ _0466_ clknet_leaf_120_wb_clk_i design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_140_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5951__C _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5150__A1 _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold31 net508 net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold20 net477 net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4139__I _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold64 wbs_dat_i[4] net482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold53 wbs_adr_i[7] net471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 net506 net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5453__A2 _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold86 wbs_dat_i[26] net504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold75 wbs_dat_i[11] net493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold97 wbs_adr_i[20] net515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4075__S _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_119_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3854__I3 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_162_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_54_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_128_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5433__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A1 _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _2601_ _2618_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_109_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_137_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3888__I _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5811_ _2270_ _2284_ _2287_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5742_ dffram.data\[40\]\[7\] _2237_ _2241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ _1582_ _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4624_ _1486_ _1489_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _1429_ _0749_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3506_ _2880_ _2873_ _2881_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _1320_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3437_ _2834_ _2836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6225_ _0182_ clknet_leaf_118_wb_clk_i dffram.data\[51\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input150_I qcpu_sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3368_ _2775_ _2780_ _2781_ _2764_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6156_ _0113_ clknet_leaf_173_wb_clk_i dffram.data\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5107_ _1816_ _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6087_ _0044_ clknet_leaf_34_wb_clk_i dffram.data\[37\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3299_ _2723_ _2719_ _2724_ _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input11_I ay8913_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5038_ _1752_ _1769_ _1771_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3997__A2 _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3749__A2 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3038__I _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__I _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5123__A1 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A2 _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput110 qcpu_do[7] net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput154 qcpu_sram_in[1] net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput132 qcpu_oeb[27] net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput121 qcpu_oeb[17] net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput143 qcpu_oeb[7] net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput165 sid_do[13] net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput176 sid_do[4] net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput187 sn76489_do[13] net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_172_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_172_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput198 sn76489_do[23] net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_101_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3501__I _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4937__A1 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4004__I3 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ _1257_ _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _1199_ _1212_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6010_ _2395_ _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ _2646_ _2662_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input3_I ay8913_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3153_ _2581_ _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3691__A4 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3084_ _2473_ wb_counter\[7\] _2542_ _2543_ _2353_ _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_134_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_102_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4928__A1 _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3986_ dffram.data\[56\]\[2\] dffram.data\[57\]\[2\] _0865_ _0933_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ _2229_ _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5338__I _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5656_ dffram.data\[41\]\[1\] _2183_ _2185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input198_I sn76489_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _1462_ _1474_ _1475_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5587_ _2138_ _2135_ _2139_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4538_ net201 _1356_ _1342_ net98 _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4469_ _1340_ _1367_ _1368_ net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_input59_I mc14500_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A1 _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6208_ _0165_ clknet_leaf_165_wb_clk_i dffram.data\[24\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6139_ _0096_ clknet_leaf_17_wb_clk_i dffram.data\[55\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4417__I _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4919__A1 _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3840_ _0718_ _0748_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_55_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__I _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3771_ net220 _0675_ _0685_ net150 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_13_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5510_ dffram.data\[45\]\[7\] _2079_ _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6490_ _0447_ clknet_leaf_145_wb_clk_i net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_140_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__A1 _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5441_ dffram.data\[46\]\[3\] _2036_ _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5372_ dffram.data\[47\]\[4\] _1993_ _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ net139 _1258_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3649__A1 _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4254_ _0679_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4185_ dffram.data\[40\]\[5\] dffram.data\[41\]\[5\] _0772_ _1129_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4310__A2 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3205_ _2641_ wb_counter\[24\] _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3136_ _2588_ _2589_ _2590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3067_ net284 _2520_ _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input113_I qcpu_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4173__S _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4216__I3 _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5708_ _2200_ _2217_ _2220_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ dffram.data\[2\]\[2\] dffram.data\[3\]\[2\] _0849_ _0916_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5068__I _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5639_ dffram.data\[17\]\[3\] _2170_ _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4129__A2 _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output332_I net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5565__A1 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4610__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2390_ _2415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _1687_ _1702_ _1707_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4872_ _1625_ _1657_ _1660_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3823_ _0771_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6611_ _0568_ clknet_leaf_2_wb_clk_i dffram.data\[33\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3754_ _0702_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6542_ _0499_ clknet_leaf_130_wb_clk_i net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6473_ _0430_ clknet_leaf_39_wb_clk_i dffram.data\[62\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3685_ _0631_ _0638_ net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_99_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__I _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5859__A2 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _2009_ _2027_ _2029_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5355_ dffram.data\[21\]\[7\] _1978_ _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput277 net277 custom_settings[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput266 net266 custom_settings[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4306_ _1247_ net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5286_ _1935_ _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput288 net288 custom_settings[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput299 net299 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4237_ dffram.data\[40\]\[6\] dffram.data\[41\]\[6\] _0772_ _1180_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4134__I2 _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ dffram.data\[58\]\[5\] dffram.data\[59\]\[5\] _0998_ _1112_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4099_ dffram.data\[4\]\[4\] dffram.data\[5\]\[4\] _0983_ _1044_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3119_ net259 _2553_ _2557_ _2575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5795__A1 _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4070__I1 dffram.data\[39\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output282_I net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__S _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3089__A2 _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3884__I1 dffram.data\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_100_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4605__I _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ dffram.data\[35\]\[4\] _2856_ _2857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5710__A1 _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5140_ dffram.data\[52\]\[5\] _1839_ _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5171__I _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5071_ dffram.data\[39\]\[1\] _1790_ _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4022_ _0764_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6018__A2 _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _2401_ _2402_ _2396_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4924_ dffram.data\[54\]\[6\] _1691_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4515__I _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3252__A2 _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5529__A1 _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4855_ _1648_ _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_63_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4786_ dffram.data\[63\]\[2\] _1599_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3806_ dffram.data\[56\]\[0\] dffram.data\[57\]\[0\] _0754_ _0755_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6525_ _0482_ clknet_leaf_142_wb_clk_i net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ net218 _0675_ _0685_ net148 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__4250__I _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input180_I sid_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _0413_ clknet_leaf_62_wb_clk_i dffram.data\[38\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3668_ design_select\[4\] design_select\[3\] _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5701__A1 _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ _2104_ _2195_ _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6387_ _0344_ clknet_leaf_70_wb_clk_i dffram.data\[17\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5407_ dffram.data\[20\]\[7\] _2011_ _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5338_ _1970_ _1972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input41_I mc14500_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5269_ _1878_ _1922_ _1925_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__B2 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__A1 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_126_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_152_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5940__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3951__B1 _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3504__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4640_ _1470_ _1497_ _1500_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2993__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4290__S0 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6310_ _0267_ clknet_leaf_128_wb_clk_i dffram.data\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4571_ dffram.data\[5\]\[0\] _1445_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3522_ dffram.data\[33\]\[5\] _2890_ _2892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3453_ _2333_ _2841_ _2845_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6241_ _0198_ clknet_leaf_125_wb_clk_i dffram.data\[50\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__B2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__A1 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6172_ _0129_ clknet_leaf_162_wb_clk_i dffram.data\[53\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5123_ _1828_ _1818_ _1829_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3384_ _2794_ _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_127_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5998__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5054_ dffram.data\[25\]\[3\] _1777_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4005_ _0886_ _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__A1 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4245__I _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5956_ net288 _2386_ _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5887_ _1647_ _2033_ _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4907_ dffram.data\[54\]\[1\] _1681_ _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4838_ _1615_ _1635_ _1638_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input89_I qcpu_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4769_ _1584_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_60_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _0465_ clknet_leaf_161_wb_clk_i design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_31_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6439_ _0396_ clknet_leaf_49_wb_clk_i dffram.data\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4489__A1 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__B2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3161__A1 net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold32 net486 net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 wbs_adr_i[23] net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5989__A1 net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold43 net509 net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 wbs_dat_i[12] net494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold87 wbs_dat_i[23] net505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5714__I _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_91_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3234__I _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4266__S _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_122_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5810_ dffram.data\[15\]\[5\] _2285_ _2287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ _2212_ _2236_ _2240_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5672_ _2060_ _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__S0 _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4623_ _1488_ _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_143_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4554_ _1188_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3505_ dffram.data\[34\]\[7\] _2874_ _2881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3391__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4485_ _1377_ _1380_ net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6224_ _0181_ clknet_leaf_119_wb_clk_i dffram.data\[51\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3436_ _2834_ _2835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6155_ _0112_ clknet_leaf_16_wb_clk_i dffram.data\[28\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3367_ net235 _2773_ _2781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3144__I _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6086_ _0043_ clknet_leaf_34_wb_clk_i dffram.data\[37\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input143_I qcpu_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _1463_ _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5037_ dffram.data\[49\]\[4\] _1770_ _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4176__S _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3298_ wb_counter\[8\] _2724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2983__I net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__I net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _2376_ _2377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output362_I net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__I _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput111 qcpu_do[8] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput100 qcpu_do[28] net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput133 qcpu_oeb[28] net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput122 qcpu_oeb[18] net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput144 qcpu_oeb[8] net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput155 qcpu_sram_in[2] net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput166 sid_do[14] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput177 sid_do[5] net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4086__S _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput199 sn76489_do[24] net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput188 sn76489_do[14] net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__A1 _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold97_I wbs_adr_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_141_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_141_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4613__I net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3229__I _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5444__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4270_ _1207_ _1208_ _1210_ _1211_ _1196_ _0786_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3221_ net389 _2654_ _2647_ _2661_ _2662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3152_ _2596_ wb_counter\[16\] _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3083_ _2384_ net213 _2482_ _2543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__I _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3985_ _0907_ _0914_ _0920_ _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_58_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5724_ _2229_ _2230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5655_ _2132_ _2182_ _2184_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ dffram.data\[5\]\[6\] _1466_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5586_ dffram.data\[43\]\[1\] _2136_ _2139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4537_ _1418_ _1419_ net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ net209 _1345_ _1277_ net111 net63 _1352_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_68_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3419_ wb_counter\[30\] _2822_ _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6207_ _0164_ clknet_leaf_162_wb_clk_i dffram.data\[24\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4399_ net136 _1250_ _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6138_ _0095_ clknet_leaf_16_wb_clk_i dffram.data\[55\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4864__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4616__A1 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6069_ _0026_ clknet_leaf_11_wb_clk_i dffram.data\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3355__A1 _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5264__I _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3107__A1 _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_86_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5032__A1 _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3770_ net69 _0683_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5440_ _2005_ _2035_ _2039_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5371_ _1985_ _1993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4322_ _1256_ _1260_ net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4253_ dffram.data\[30\]\[7\] dffram.data\[31\]\[7\] _1194_ _1195_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4846__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3204_ _2549_ _2647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4184_ _0700_ _1127_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3135_ net261 _2582_ _2583_ _2589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3066_ _1110_ _1135_ _2503_ _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_2_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input106_I qcpu_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5023__A1 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ dffram.data\[0\]\[2\] dffram.data\[1\]\[2\] _0662_ _0915_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5707_ dffram.data\[16\]\[1\] _2218_ _2220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _0700_ _0846_ _0723_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_73_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input71_I mc14500_sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _2140_ _2169_ _2173_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5569_ _2119_ _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4152__I3 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output325_I net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3332__I _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5262__A1 _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__C1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5014__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3966__I3 _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4128__I0 _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4828__A1 _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3500__A1 _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ dffram.data\[28\]\[3\] _1703_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4871_ dffram.data\[56\]\[5\] _1658_ _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3822_ _0707_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6610_ _0567_ clknet_leaf_3_wb_clk_i dffram.data\[33\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3567__A1 _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _0498_ clknet_leaf_130_wb_clk_i net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3753_ _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6472_ _0429_ clknet_leaf_38_wb_clk_i dffram.data\[62\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3684_ _0636_ _0637_ _0626_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_132_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5423_ dffram.data\[0\]\[4\] _2028_ _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5354_ _1951_ _1977_ _1981_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4305_ _1221_ _1246_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xoutput267 net267 custom_settings[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5632__I _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput278 net278 custom_settings[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4819__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5285_ _1830_ _1649_ _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput289 net289 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4236_ _0700_ _1178_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4167_ dffram.data\[56\]\[5\] dffram.data\[57\]\[5\] _0799_ _1111_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3118_ _2572_ _2573_ _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4098_ dffram.data\[2\]\[4\] dffram.data\[3\]\[4\] _0849_ _1043_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_143_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5795__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3049_ net282 _2479_ _2513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_142_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3558__A1 dffram.data\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__I _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output275_I net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3730__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3011__B _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3549__A1 _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4269__S _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _1741_ _1789_ _1791_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4021_ dffram.data\[30\]\[3\] dffram.data\[31\]\[3\] _0904_ _0967_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5226__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3700__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ net226 _2391_ _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4923_ _1561_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4854_ _1631_ _1507_ _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4785_ _1545_ _1598_ _1601_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3805_ _0753_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3736_ _0677_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6524_ _0481_ clknet_leaf_139_wb_clk_i net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6455_ _0412_ clknet_leaf_64_wb_clk_i dffram.data\[38\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input173_I sid_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3667_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_31_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3598_ _2940_ _2933_ _2941_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6386_ _0343_ clknet_4_12_0_wb_clk_i dffram.data\[17\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5406_ _1827_ _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5337_ _1970_ _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5268_ dffram.data\[22\]\[1\] _1923_ _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4107__I3 _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I mc14500_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ dffram.data\[56\]\[6\] dffram.data\[57\]\[6\] _0799_ _1162_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5199_ _1878_ _1875_ _1879_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__C1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_166_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_166_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3721__S _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ _1440_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4290__S1 _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3521_ _2872_ _2889_ _2891_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmax_cap403 _1447_ net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3452_ dffram.data\[36\]\[6\] _2842_ _2845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _0197_ clknet_leaf_123_wb_clk_i dffram.data\[50\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5695__A1 _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__I _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6171_ _0128_ clknet_leaf_169_wb_clk_i dffram.data\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3383_ _2787_ _2786_ _2793_ _2782_ _2794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_5122_ dffram.data\[24\]\[7\] _1819_ _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5053_ _1748_ _1776_ _1780_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4004_ _0945_ _0947_ _0948_ _0950_ _0801_ _0802_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_140_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5955_ _2387_ _2388_ _2381_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_36_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5886_ _2335_ _2328_ _2336_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4906_ _1544_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4837_ dffram.data\[57\]\[1\] _1636_ _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _1551_ _1585_ _1590_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4699_ _1540_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3719_ _0664_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6507_ _0464_ clknet_leaf_122_wb_clk_i net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _0395_ clknet_leaf_49_wb_clk_i dffram.data\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _0326_ clknet_leaf_100_wb_clk_i dffram.data\[43\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold22 _2356_ net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold11 _2829_ net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 net503 net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 net496 net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 wbs_adr_i[6] net473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3839__I2 _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold66 wbs_dat_i[2] net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold77 wbs_dat_i[25] net495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold88 wbs_dat_i[29] net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4436__I _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_91_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5601__A1 _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5740_ dffram.data\[40\]\[6\] _2237_ _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4282__S _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5671_ _2152_ _2188_ _2193_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4622_ _1487_ _1437_ _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4263__S1 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4553_ _0639_ _1428_ net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ net164 _1348_ _1378_ net83 net4 _1379_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_3504_ _1477_ _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3435_ _1568_ _2118_ _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6223_ _0180_ clknet_leaf_123_wb_clk_i dffram.data\[51\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6154_ _0111_ clknet_leaf_14_wb_clk_i dffram.data\[28\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3366_ wb_counter\[20\] _2779_ _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6085_ _0042_ clknet_leaf_34_wb_clk_i dffram.data\[37\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3297_ wb_counter\[7\] _2723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5105_ _1814_ _1804_ _1815_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input136_I qcpu_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _1762_ _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5938_ _2359_ _2376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5869_ _2323_ _2318_ _2324_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5659__A1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4182__I1 dffram.data\[39\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput101 qcpu_do[29] net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput134 qcpu_oeb[29] net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput123 qcpu_oeb[19] net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput145 qcpu_oeb[9] net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 qcpu_do[9] net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput156 qcpu_sram_in[3] net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput167 sid_do[15] net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput178 sid_do[6] net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput189 sn76489_do[15] net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3996__I1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5725__I _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_120_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3220_ _2659_ _2660_ _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3151_ _2550_ _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4076__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__A1 _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3082_ net362 _2477_ _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_38_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3984_ _0921_ _0930_ _0750_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _2133_ _2019_ _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_84_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ dffram.data\[41\]\[0\] _2183_ _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _1473_ _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5585_ _2067_ _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4536_ net51 _1414_ _1357_ net18 _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4467_ net180 _1348_ _1350_ net27 _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4398_ _1302_ _1309_ net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4313__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _0163_ clknet_leaf_156_wb_clk_i dffram.data\[24\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3418_ wb_counter\[28\] wb_counter\[29\] _2816_ _2822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _0094_ clknet_leaf_16_wb_clk_i dffram.data\[55\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3349_ wb_counter\[16\] wb_counter\[17\] _2766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5370__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5813__A1 _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_77_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4616__A2 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6068_ _0025_ clknet_leaf_11_wb_clk_i dffram.data\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5019_ dffram.data\[53\]\[6\] _1754_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3052__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_95_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__A2 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5455__I _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A1 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ _1985_ _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ net135 _1258_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _0777_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3203_ _2363_ _2646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4183_ _1123_ _1124_ _1125_ _1126_ _0765_ _0766_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_59_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3134_ _2572_ wb_counter\[13\] _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3065_ _2511_ _2527_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3967_ _0908_ _0913_ _0723_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_132_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _2194_ _2217_ _2219_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3898_ _0841_ _0842_ _0844_ _0845_ _0713_ _0715_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_66_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5637_ dffram.data\[17\]\[2\] _2170_ _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__A1 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _2119_ _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input64_I mc14500_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4519_ net196 _1402_ _1403_ net93 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5499_ _2077_ _2078_ _2080_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output318_I net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_171_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5275__I _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3959__S0 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _1621_ _1657_ _1659_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3821_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4764__A1 _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6540_ _0497_ clknet_leaf_131_wb_clk_i net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3752_ _0659_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _0428_ clknet_leaf_42_wb_clk_i dffram.data\[62\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3683_ _0621_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4303__B _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5422_ _2020_ _2028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4516__B2 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ dffram.data\[21\]\[6\] _1978_ _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _1227_ _1233_ _1239_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput257 net257 custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput268 net268 custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5284_ _1801_ _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput279 net279 custom_settings[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4529__I _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4235_ _1174_ _1175_ _1176_ _1177_ _0765_ _0766_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_52_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4166_ _1091_ _1097_ _1103_ _1109_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3117_ wb_counter\[11\] _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4097_ dffram.data\[0\]\[4\] dffram.data\[1\]\[4\] _0980_ _1042_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input216_I wbs_adr_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3048_ _0996_ _1027_ _2503_ _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_26_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__A1 _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4999_ dffram.data\[53\]\[0\] _1744_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__A1 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A1 _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output268_I net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4294__I0 dffram.data\[36\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__A1 _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__I _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3549__A2 _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold72_I wbs_dat_i[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_88_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3518__I _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_17_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_12_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4020_ dffram.data\[28\]\[3\] dffram.data\[29\]\[3\] _0831_ _0966_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ net260 _2400_ _2401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4922_ _1693_ _1690_ _1694_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_32_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4853_ _1503_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4812__I _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__I net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4784_ dffram.data\[63\]\[1\] _1599_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3804_ _0664_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3735_ net67 _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _0480_ clknet_leaf_141_wb_clk_i net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _0411_ clknet_leaf_62_wb_clk_i dffram.data\[38\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3960__A2 _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _2015_ _2010_ _2016_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3666_ design_select\[2\] _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_70_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__A1 _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3597_ dffram.data\[60\]\[7\] _2934_ _2941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6385_ _0342_ clknet_leaf_86_wb_clk_i dffram.data\[17\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _1858_ _1439_ _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input166_I sid_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _1873_ _1922_ _1924_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _1142_ _1148_ _1154_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_input27_I ay8913_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ dffram.data\[50\]\[1\] _1876_ _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4149_ dffram.data\[18\]\[5\] dffram.data\[19\]\[5\] _0972_ _1093_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_50_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4425__C2 _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4728__A1 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3467__A1 _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_135_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_135_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3801__I _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__A1 net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3520_ dffram.data\[33\]\[4\] _2890_ _2891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap404 _1442_ net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_96_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3451_ _2331_ _2841_ _2844_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3382_ wb_counter\[23\] _2793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_23_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6170_ _0127_ clknet_leaf_171_wb_clk_i dffram.data\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5121_ _1827_ _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3912__S _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5052_ dffram.data\[25\]\[2\] _1777_ _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4003_ dffram.data\[38\]\[2\] dffram.data\[39\]\[2\] _0949_ _0950_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3711__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A1 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5954_ net253 _2377_ _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3630__A1 _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5885_ dffram.data\[14\]\[7\] _2329_ _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _1678_ _1680_ _1682_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4836_ _1610_ _1635_ _1637_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4767_ dffram.data\[59\]\[3\] _1586_ _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6506_ _0463_ clknet_leaf_133_wb_clk_i net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_113_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4698_ _1431_ _1509_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3718_ dffram.data\[26\]\[0\] dffram.data\[27\]\[0\] _0666_ _0667_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3649_ _2928_ _2969_ _2973_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6437_ _0394_ clknet_leaf_50_wb_clk_i dffram.data\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5135__A1 _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2997__I _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ _0325_ clknet_leaf_96_wb_clk_i dffram.data\[43\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ _1934_ _1958_ _1960_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3697__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6299_ _0256_ clknet_leaf_111_wb_clk_i dffram.data\[47\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold12 net484 net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold23 net432 net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3449__A1 _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold45 net487 net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold34 net493 net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold56 wbs_dat_i[5] net474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3621__I _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3839__I3 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold89 wbs_dat_i[18] net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold78 wbs_dat_i[21] net496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output300_I net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4452__I _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ dffram.data\[41\]\[7\] _2189_ _2193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5365__A1 _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _0682_ _1089_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ net105 _1250_ _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4483_ _0650_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3503_ _2878_ _2873_ _2879_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5193__I _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _0179_ clknet_leaf_123_wb_clk_i dffram.data\[51\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3434_ _2833_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_115_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6153_ _0110_ clknet_leaf_13_wb_clk_i dffram.data\[28\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3365_ _2614_ wb_counter\[19\] _2768_ _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5921__I _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6084_ _0041_ clknet_leaf_34_wb_clk_i dffram.data\[37\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3296_ _2708_ _2720_ _2722_ _2718_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5104_ dffram.data\[24\]\[3\] _1805_ _1815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _1762_ _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input129_I qcpu_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3603__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5937_ net283 _2372_ _2375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ dffram.data\[14\]\[2\] _2319_ _2324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input94_I qcpu_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5799_ _2255_ _2278_ _2280_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5356__A1 _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _1621_ _1622_ _1624_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output348_I net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput102 qcpu_do[2] net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_hold5_I net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput135 qcpu_oeb[2] net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput124 qcpu_oeb[1] net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 qcpu_oeb[0] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 qcpu_sram_in[4] net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4447__I _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput168 sid_do[16] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput146 qcpu_sram_addr[0] net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput179 sid_do[7] net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_129_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A2 _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_150_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_150_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3150_ _2546_ _2601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3081_ _2370_ _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_124_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4293__S _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _2214_ _2223_ _2228_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3983_ _0922_ _0924_ _0925_ _0927_ _0928_ _0929_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_102_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3061__A2 _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5653_ _2181_ _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5584_ _2132_ _2135_ _2137_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4604_ _1472_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_135_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4535_ net200 _1356_ _1342_ net97 _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3436__I _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4561__A2 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4466_ _1336_ _1365_ _1366_ net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4397_ net134 _1250_ _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4313__A2 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _0162_ clknet_leaf_156_wb_clk_i dffram.data\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3417_ _2765_ _2820_ _2821_ _2806_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6136_ _0093_ clknet_leaf_168_wb_clk_i dffram.data\[55\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ _2690_ _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6067_ _0024_ clknet_leaf_20_wb_clk_i dffram.data\[58\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3171__I _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3279_ wb_counter\[0\] wb_counter\[1\] wb_counter\[2\] wb_counter\[3\] _2709_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA_clkbuf_leaf_161_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _1561_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_138_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5577__A1 _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5098__I _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5329__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output298_I net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__A2 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3043__A2 _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _1256_ _1259_ net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4251_ dffram.data\[28\]\[7\] dffram.data\[29\]\[7\] _1192_ _1193_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4288__S _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3202_ _2624_ _2645_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input1_I ay8913_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4182_ dffram.data\[38\]\[5\] dffram.data\[39\]\[5\] _0949_ _1126_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3133_ _2561_ _2587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3064_ net397 _2518_ _2524_ _2526_ _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3966_ _0909_ _0910_ _0911_ _0912_ _0713_ _0715_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_85_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ dffram.data\[16\]\[0\] _2218_ _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5636_ _2138_ _2169_ _2172_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3897_ dffram.data\[22\]\[1\] dffram.data\[23\]\[1\] _0711_ _0845_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input196_I sn76489_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5567_ _2074_ _2120_ _2125_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5731__A1 _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ dffram.data\[45\]\[4\] _2079_ _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4518_ _1404_ _1405_ net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_57_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input57_I mc14500_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _1347_ _1351_ _1353_ net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_106_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _0076_ clknet_leaf_0_wb_clk_i dffram.data\[57\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4725__I _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__B2 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__A1 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A1 _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3959__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3804__I _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3025__B _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4635__I _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4461__B2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__A1 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3820_ _0698_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_119_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3751_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5961__A1 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6470_ _0427_ clknet_leaf_42_wb_clk_i dffram.data\[62\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3682_ design_select\[1\] _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_82_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5421_ _2020_ _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _1949_ _1977_ _1980_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4303_ _1188_ _1244_ _0818_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput258 net258 custom_settings[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5283_ _1892_ _1928_ _1933_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput269 net269 custom_settings[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ dffram.data\[38\]\[6\] dffram.data\[39\]\[6\] _0762_ _1177_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4165_ _0921_ _1108_ _1053_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_52_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3116_ _2571_ _2572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4096_ _0908_ _1039_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_143_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input111_I qcpu_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3047_ _1481_ _2511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3255__A2 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input209_I sn76489_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ _1742_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3949_ _0893_ _0894_ _0895_ _0896_ _0815_ _0816_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_34_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ _2154_ _2161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6599_ _0556_ clknet_leaf_32_wb_clk_i dffram.data\[34\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6000__I _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output330_I net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5286__I _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5943__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_114_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3182__A1 net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4434__A1 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _2399_ _2400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4921_ dffram.data\[54\]\[5\] _1691_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _1629_ _1641_ _1646_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2996__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3803_ _0697_ _0724_ _0732_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_90_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4783_ _1539_ _1598_ _1600_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5934__A1 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ _0673_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _0479_ clknet_4_10_0_wb_clk_i net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6453_ _0410_ clknet_leaf_63_wb_clk_i dffram.data\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3665_ design_select\[0\] _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5404_ dffram.data\[20\]\[6\] _2011_ _2016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6384_ _0341_ clknet_leaf_85_wb_clk_i dffram.data\[17\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3596_ _1477_ _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3173__A1 net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5335_ _1953_ _1964_ _1969_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input159_I qcpu_sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5266_ dffram.data\[22\]\[0\] _1923_ _1924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4217_ _0806_ _1159_ _1053_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5197_ _1807_ _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4148_ dffram.data\[16\]\[5\] dffram.data\[17\]\[5\] _0742_ _1092_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4079_ _1020_ _1021_ _1023_ _1024_ _0815_ _0816_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__4425__A1 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4425__B2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4284__S0 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A1 net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output280_I net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_175_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_175_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_104_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3529__I _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__A1 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3450_ dffram.data\[36\]\[5\] _2842_ _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3155__A1 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3381_ _2690_ _2792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5120_ _1476_ _1827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _1746_ _1776_ _1779_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_127_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4002_ _0761_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_140_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4823__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ net287 _2386_ _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ _1477_ _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_105_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4904_ dffram.data\[54\]\[0\] _1681_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ dffram.data\[57\]\[0\] _1636_ _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _1548_ _1585_ _1589_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3717_ _0665_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6505_ _0462_ clknet_leaf_129_wb_clk_i net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ _1538_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3648_ dffram.data\[9\]\[2\] _2970_ _2973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6436_ _0393_ clknet_leaf_50_wb_clk_i dffram.data\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3579_ _1454_ _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6367_ _0324_ clknet_leaf_95_wb_clk_i dffram.data\[43\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3146__A1 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ dffram.data\[8\]\[0\] _1959_ _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6298_ _0255_ clknet_leaf_70_wb_clk_i dffram.data\[47\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold13 _2369_ net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5249_ dffram.data\[7\]\[2\] _1910_ _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold24 net499 net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 net511 net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold35 net492 net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 wbs_dat_i[27] net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold68 wbs_dat_i[31] net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_97_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5071__A1 dffram.data\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4885__A1 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__I _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _1485_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _1427_ net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_143_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5474__I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_72_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__B1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__C2 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4482_ _1276_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3502_ dffram.data\[34\]\[6\] _2874_ _2879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6221_ _0178_ clknet_leaf_123_wb_clk_i dffram.data\[51\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3433_ net370 _2541_ _2831_ _2832_ _2833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_122_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4876__A1 _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _0109_ clknet_leaf_13_wb_clk_i dffram.data\[28\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5103_ _1813_ _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3364_ _2775_ _2777_ _2778_ _2764_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6083_ _0040_ clknet_leaf_67_wb_clk_i dffram.data\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3722__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3295_ net252 _2721_ _2722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4628__A1 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _1750_ _1763_ _1768_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_151_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3300__A1 _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__A1 _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5936_ _2373_ net424 _2364_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5867_ _1454_ _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5798_ dffram.data\[15\]\[0\] _2279_ _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4818_ dffram.data\[6\]\[4\] _1623_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3367__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input87_I qcpu_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4749_ _1554_ _1576_ _1578_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _0376_ clknet_leaf_85_wb_clk_i dffram.data\[40\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3119__A1 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3632__I _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput136 qcpu_oeb[30] net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput125 qcpu_oeb[20] net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput114 qcpu_oeb[10] net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput103 qcpu_do[30] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput158 qcpu_sram_in[5] net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput169 sid_do[17] net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput147 qcpu_sram_addr[1] net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5292__A1 _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__A2 _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5559__I _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5044__A1 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3996__I3 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3358__A1 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3807__I _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3028__B _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__I0 _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ _2511_ _2540_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5283__A1 _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3982_ _0745_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5721_ dffram.data\[16\]\[7\] _2224_ _2228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5652_ _2181_ _2182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ net251 _1311_ _1457_ net159 _0644_ net78 _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_5583_ dffram.data\[43\]\[0\] _2136_ _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4534_ _1416_ _1417_ net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_135_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4561__A3 _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4465_ net208 _1322_ _1361_ net26 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4164__I3 _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4396_ _1303_ _1308_ net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3416_ net244 _2814_ _2821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6204_ _0161_ clknet_leaf_162_wb_clk_i dffram.data\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3521__A1 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _2752_ _2762_ _2763_ _2764_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6135_ _0092_ clknet_leaf_170_wb_clk_i dffram.data\[55\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input141_I qcpu_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ _0023_ clknet_leaf_20_wb_clk_i dffram.data\[58\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5017_ _1756_ _1753_ _1757_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3278_ _2707_ _2708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ net420 _2360_ _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4458__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_106_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__C1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5017__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4193__I _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold95_I wbs_dat_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_143_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4250_ _0777_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4181_ dffram.data\[36\]\[5\] dffram.data\[37\]\[5\] _0759_ _1125_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3503__A1 _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ net386 _2632_ _2625_ _2644_ _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3132_ _2578_ _2586_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A1 _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__C1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3063_ _0647_ _2525_ _2499_ _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3965_ dffram.data\[22\]\[2\] dffram.data\[23\]\[2\] _0711_ _0912_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5927__I net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _2216_ _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3896_ dffram.data\[20\]\[1\] dffram.data\[21\]\[1\] _0843_ _0844_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5635_ dffram.data\[17\]\[1\] _2170_ _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3447__I _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5566_ dffram.data\[44\]\[3\] _2121_ _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input189_I sn76489_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5497_ _2063_ _2079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5662__I _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4517_ net173 _1396_ _1359_ net46 net13 _1318_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_57_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4448_ net204 _1345_ _1277_ net106 net58 _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4379_ _1296_ _1298_ net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_95_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _0075_ clknet_leaf_0_wb_clk_i dffram.data\[57\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6049_ _0006_ clknet_leaf_19_wb_clk_i dffram.data\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3357__I _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_129_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4128__I3 _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3306__B _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5238__A1 _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold10_I wbs_adr_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4916__I _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3750_ _0698_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5410__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3681_ _0632_ _0630_ _0635_ net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_55_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5420_ _2007_ _2021_ _2026_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5482__I _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__S _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3724__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ dffram.data\[21\]\[5\] _1978_ _1980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4302_ _1240_ _1241_ _1242_ _1243_ _0834_ _0882_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_5282_ dffram.data\[22\]\[7\] _1929_ _1933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput259 net259 custom_settings[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5477__A1 _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ dffram.data\[36\]\[6\] dffram.data\[37\]\[6\] _0759_ _1176_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3931__S _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4164_ _1104_ _1105_ _1106_ _1107_ _0928_ _0929_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4095_ _0722_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3115_ _2471_ _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3046_ _1482_ _2510_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input104_I qcpu_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1742_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3948_ dffram.data\[46\]\[1\] dffram.data\[47\]\[1\] _0813_ _0896_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3879_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5618_ _2142_ _2155_ _2160_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ _0555_ clknet_leaf_32_wb_clk_i dffram.data\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5549_ _2077_ _2112_ _2114_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output323_I net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__I _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6386__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__A1 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3087__I _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3815__I _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A1 _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4646__I _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_26_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3550__I _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4920_ _1558_ _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ dffram.data\[57\]\[7\] _1642_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3802_ _0733_ _0747_ _0750_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4782_ dffram.data\[63\]\[0\] _1599_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3733_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6521_ _0478_ clknet_leaf_139_wb_clk_i net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3664_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6452_ _0409_ clknet_leaf_64_wb_clk_i dffram.data\[38\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5698__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _1824_ _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3595_ _2938_ _2933_ _2939_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6383_ _0340_ clknet_leaf_88_wb_clk_i dffram.data\[17\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5334_ dffram.data\[8\]\[7\] _1965_ _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5265_ _1921_ _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4216_ _1155_ _1156_ _1157_ _1158_ _0713_ _0715_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5196_ _1873_ _1875_ _1877_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4147_ _0696_ _1090_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5622__A1 _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4078_ dffram.data\[46\]\[3\] dffram.data\[47\]\[3\] _0957_ _1024_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3029_ net268 _2479_ _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4284__S1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output273_I net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_144_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_144_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4352__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3380_ _2775_ _2789_ _2791_ _2785_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5050_ dffram.data\[25\]\[1\] _1777_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4001_ dffram.data\[36\]\[2\] dffram.data\[37\]\[2\] _0797_ _0948_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_141_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5604__A1 _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5952_ net440 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_140_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _1679_ _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5883_ _2333_ _2328_ _2334_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ _1634_ _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4765_ dffram.data\[59\]\[2\] _1586_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3716_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6504_ _0461_ clknet_leaf_129_wb_clk_i net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ net404 _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3647_ _2926_ _2969_ _2972_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6435_ _0392_ clknet_leaf_63_wb_clk_i dffram.data\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input171_I sid_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3578_ _2926_ _2923_ _2927_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6366_ _0323_ clknet_leaf_94_wb_clk_i dffram.data\[43\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5317_ _1957_ _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _0254_ clknet_leaf_111_wb_clk_i dffram.data\[47\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold14 wbs_adr_i[22] net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_input32_I hellorld_do vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__A1 _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _1878_ _1909_ _1912_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold47 net510 net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold36 net504 net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 net490 net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3404__B _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold58 _0676_ net476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5179_ dffram.data\[23\]\[3\] _1862_ _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold69 wbs_dat_i[17] net487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_39_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3082__A1 net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5834__A1 _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4573__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4573__B2 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ net104 _1258_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_123_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4481_ net186 _1333_ _1375_ net37 _1376_ _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_3501_ _1473_ _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _0177_ clknet_leaf_123_wb_clk_i dffram.data\[51\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3432_ _2473_ _2350_ _2353_ _2477_ _2832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3363_ net233 _2773_ _2778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6151_ _0108_ clknet_leaf_173_wb_clk_i dffram.data\[28\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5490__I _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5102_ _1458_ _1813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4100__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6082_ _0039_ clknet_leaf_22_wb_clk_i dffram.data\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3294_ _2704_ _2721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_29_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5033_ dffram.data\[49\]\[3\] _1764_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3300__A2 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__I _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5935_ net423 _2360_ _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3064__A1 net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _2321_ _2318_ _2322_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4817_ _1611_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6002__A1 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _2277_ _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4748_ dffram.data\[37\]\[4\] _1577_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _1444_ _1526_ _1528_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6418_ _0375_ clknet_leaf_87_wb_clk_i dffram.data\[40\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _0306_ clknet_leaf_78_wb_clk_i dffram.data\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5816__A1 _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput126 qcpu_oeb[21] net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput115 qcpu_oeb[11] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput104 qcpu_do[31] net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput159 qcpu_sram_in[6] net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput137 qcpu_oeb[31] net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput148 qcpu_sram_addr[2] net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_99_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3823__I _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3913__S0 _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _0681_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__I0 _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5720_ _2212_ _2223_ _2227_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_102_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5651_ _2133_ _2167_ _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_26_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A1 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__B2 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _2134_ _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4602_ _1462_ _1470_ _1471_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4533_ net50 _1414_ _1408_ net17 _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_135_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ net179 _1344_ _1331_ net110 net62 _1354_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6203_ _0160_ clknet_leaf_19_wb_clk_i dffram.data\[39\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4395_ net133 _1304_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_99_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3733__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3415_ wb_counter\[29\] _2819_ _2820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _2700_ _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6134_ _0091_ clknet_leaf_170_wb_clk_i dffram.data\[55\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6065_ _0022_ clknet_leaf_26_wb_clk_i dffram.data\[58\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input134_I qcpu_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ dffram.data\[53\]\[5\] _1754_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3277_ _2692_ _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3285__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4785__A1 _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ _2359_ _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5849_ _2303_ _2311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4537__A1 _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output353_I net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3643__I _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__C2 _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3028__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__A1 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold88_I wbs_dat_i[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4528__B2 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4180_ dffram.data\[34\]\[5\] dffram.data\[35\]\[5\] _0946_ _1124_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3200_ _2642_ _2643_ _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3131_ net374 _2562_ _2579_ _2585_ _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3267__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3062_ _2455_ _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4464__C2 _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__S _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3964_ dffram.data\[20\]\[2\] dffram.data\[21\]\[2\] _0843_ _0911_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5703_ _2216_ _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3895_ _0708_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5634_ _2132_ _2169_ _2171_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__B2 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5565_ _2071_ _2120_ _2124_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ _2063_ _2078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4516_ net195 _1402_ _1403_ net92 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4447_ _1323_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_1_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_70_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _0074_ clknet_leaf_9_wb_clk_i dffram.data\[57\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3329_ _2704_ _2750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6048_ _0005_ clknet_leaf_19_wb_clk_i dffram.data\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4302__S0 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_169_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_169_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_9_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3497__A1 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3322__B _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__I _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__A1 _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5410__A2 _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3421__A1 _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3680_ _0634_ _0626_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__3709__C1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5174__A1 _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _1945_ _1977_ _1979_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ dffram.data\[46\]\[7\] dffram.data\[47\]\[7\] _0827_ _1243_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5281_ _1890_ _1928_ _1932_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5477__A2 _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4232_ dffram.data\[34\]\[6\] dffram.data\[35\]\[6\] _0757_ _1175_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ dffram.data\[14\]\[5\] dffram.data\[15\]\[5\] _0926_ _1107_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_52_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4437__B1 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4094_ _1035_ _1036_ _1037_ _1038_ _0976_ _0977_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3114_ _2547_ _2570_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ net393 _2470_ _2508_ _2509_ _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4988__A1 _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5938__I _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4996_ _1664_ _1439_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3947_ dffram.data\[44\]\[1\] dffram.data\[45\]\[1\] _0811_ _0895_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3412__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3458__I _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3878_ _0658_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5617_ dffram.data\[42\]\[3\] _2156_ _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6597_ _0554_ clknet_leaf_32_wb_clk_i dffram.data\[34\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ dffram.data\[18\]\[4\] _2113_ _2114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input62_I mc14500_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _2063_ _2065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3479__A1 _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output316_I net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3651__A1 _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5156__A1 _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_131_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _1627_ _1641_ _1645_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3801_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4781_ _1597_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3278__I _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _0477_ clknet_leaf_134_wb_clk_i net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3732_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _0408_ clknet_leaf_57_wb_clk_i dffram.data\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3663_ _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6382_ _0339_ clknet_leaf_88_wb_clk_i dffram.data\[17\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4103__S _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ _2013_ _2010_ _2014_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_170_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3594_ dffram.data\[60\]\[6\] _2934_ _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5333_ _1951_ _1964_ _1968_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3942__S _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _1921_ _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_10_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4215_ dffram.data\[14\]\[6\] dffram.data\[15\]\[6\] _0740_ _1158_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5195_ dffram.data\[50\]\[0\] _1876_ _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3741__I _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ _1084_ _1085_ _1086_ _1087_ _0968_ _1089_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4077_ dffram.data\[44\]\[3\] dffram.data\[45\]\[3\] _1022_ _1023_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3028_ _0863_ _0899_ _2477_ _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4979_ dffram.data\[26\]\[1\] _1730_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _0606_ clknet_leaf_48_wb_clk_i dffram.data\[61\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output266_I net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__I _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3872__A1 _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3624__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5578__I _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__I _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A1 _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold70_I wbs_dat_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3826__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_113_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3561__I _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ dffram.data\[34\]\[2\] dffram.data\[35\]\[2\] _0946_ _0947_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_144_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3615__A1 _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5951_ _2384_ _2357_ _2385_ _2371_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4902_ _1679_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5882_ dffram.data\[14\]\[6\] _2329_ _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _1634_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _1545_ _1585_ _1588_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3715_ _0659_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_60_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6503_ _0460_ clknet_leaf_132_wb_clk_i net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_114_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6434_ _0391_ clknet_leaf_63_wb_clk_i dffram.data\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4695_ _1478_ _1532_ _1537_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3646_ dffram.data\[9\]\[1\] _2970_ _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3577_ dffram.data\[60\]\[1\] _2924_ _2927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6365_ _0322_ clknet_leaf_94_wb_clk_i dffram.data\[43\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ _1957_ _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6296_ _0253_ clknet_leaf_111_wb_clk_i dffram.data\[47\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input164_I sid_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ dffram.data\[7\]\[1\] _1910_ _1912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold37 net497 net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold15 wbs_dat_i[6] net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold26 net489 net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I ay8913_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ _1811_ _1861_ _1865_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold59 wbs_adr_i[21] net477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold48 net512 net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4129_ _0886_ _1073_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4008__S _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3082__A2 _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__A1 _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3847__S _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5531__A1 _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3381__I _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5598__A1 _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_122_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A1 _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3500_ _2876_ _2873_ _2877_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4480_ _1337_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5771__I _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3431_ net436 _2554_ wb_sram_we _2831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3362_ wb_counter\[19\] _2776_ _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6150_ _0107_ clknet_leaf_176_wb_clk_i dffram.data\[28\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5101_ _1811_ _1804_ _1812_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6081_ _0038_ clknet_leaf_64_wb_clk_i dffram.data\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3293_ wb_counter\[7\] _2719_ _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_81_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5032_ _1748_ _1763_ _1767_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3300__A3 _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_10_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5934_ net282 _2372_ _2373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3064__A2 _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5865_ dffram.data\[14\]\[1\] _2319_ _2322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _1611_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ _2277_ _2278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4747_ _1569_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4678_ dffram.data\[30\]\[0\] _1527_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3629_ dffram.data\[61\]\[3\] _2957_ _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6417_ _0374_ clknet_leaf_87_wb_clk_i dffram.data\[40\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6348_ _0305_ clknet_leaf_79_wb_clk_i dffram.data\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _0236_ clknet_leaf_74_wb_clk_i dffram.data\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput127 qcpu_oeb[22] net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput116 qcpu_oeb[12] net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_73_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput105 qcpu_do[32] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput138 qcpu_oeb[32] net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5816__A2 _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput149 qcpu_sram_addr[3] net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__I _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5752__A1 _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4555__A2 _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3913__S1 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3980_ dffram.data\[14\]\[2\] dffram.data\[15\]\[2\] _0926_ _0927_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__I1 _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5991__A1 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _2152_ _2175_ _2180_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_102_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ dffram.data\[5\]\[5\] _1466_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5743__A1 _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5581_ _2134_ _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ net199 _1402_ _1403_ net96 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_26_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _1347_ _1363_ _1364_ net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_29_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6202_ _0159_ clknet_leaf_20_wb_clk_i dffram.data\[39\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3414_ _2670_ _2816_ _2819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4394_ _1303_ _1307_ net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3345_ net230 _2750_ _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6133_ _0090_ clknet_leaf_170_wb_clk_i dffram.data\[55\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6064_ _0021_ clknet_leaf_26_wb_clk_i dffram.data\[58\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3276_ _2691_ _2703_ _2706_ _2701_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5015_ _1558_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input127_I qcpu_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5917_ net213 net256 _2354_ _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5982__A1 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5848_ _2303_ _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input92_I qcpu_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5779_ _2264_ _2257_ _2265_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Left_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4021__S _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__B2 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3130_ _2580_ _2584_ _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__B2 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__A1 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__S0 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3267__A2 _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3061_ _2502_ _2519_ _2521_ _2523_ _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_89_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3019__A2 _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__I _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ dffram.data\[18\]\[2\] dffram.data\[19\]\[2\] _0705_ _0910_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3894_ dffram.data\[18\]\[1\] dffram.data\[19\]\[1\] _0705_ _0842_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5702_ _2104_ _2019_ _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__A1 _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ dffram.data\[17\]\[0\] _2170_ _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5564_ dffram.data\[44\]\[2\] _2121_ _2124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4515_ _1341_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5495_ _2076_ _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ net175 _1348_ _1350_ net22 _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_106_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4377_ _1253_ _1289_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_95_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _0073_ clknet_leaf_4_wb_clk_i dffram.data\[57\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3328_ wb_counter\[13\] _2748_ _2749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4575__I _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A1 _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6047_ _0004_ clknet_leaf_19_wb_clk_i dffram.data\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3259_ _2692_ _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4302__S1 _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A2 _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output296_I net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__A1 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4446__B2 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3829__I _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__A1 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3709__B1 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4300_ dffram.data\[44\]\[7\] dffram.data\[45\]\[7\] _1216_ _1242_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ dffram.data\[22\]\[6\] _1929_ _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4231_ dffram.data\[32\]\[6\] dffram.data\[33\]\[6\] _0754_ _1174_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4685__A1 _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ dffram.data\[12\]\[5\] dffram.data\[13\]\[5\] _0991_ _1106_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_74_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_52_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4437__A1 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4093_ dffram.data\[22\]\[4\] dffram.data\[23\]\[4\] _0709_ _1038_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3113_ net372 _2562_ _2551_ _2569_ _2570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4437__B2 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3044_ _1278_ _2489_ _2499_ _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4296__S0 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5937__A1 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ _1538_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3946_ dffram.data\[42\]\[1\] dffram.data\[43\]\[1\] _0809_ _0894_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input194_I sn76489_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ dffram.data\[24\]\[1\] dffram.data\[25\]\[1\] _0824_ _0825_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _2140_ _2155_ _2159_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6596_ _0553_ clknet_leaf_38_wb_clk_i dffram.data\[35\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5547_ _2105_ _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _2063_ _2064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input55_I mc14500_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4429_ _1327_ _1335_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XPHY_EDGE_ROW_92_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3479__A2 _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4428__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output309_I net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__I _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5864__I _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3167__A1 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__I _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4780_ _1597_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3800_ _0718_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3731_ _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5774__I _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_35_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _0407_ clknet_leaf_58_wb_clk_i dffram.data\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ design_select\[1\] _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_71_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6381_ _0338_ clknet_leaf_88_wb_clk_i dffram.data\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3593_ _1473_ _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5401_ dffram.data\[20\]\[5\] _2011_ _2014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3294__I _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5332_ dffram.data\[8\]\[6\] _1965_ _1968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _1858_ _1524_ _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4214_ dffram.data\[12\]\[6\] dffram.data\[13\]\[6\] _0991_ _1157_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5194_ _1874_ _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4145_ _1088_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3330__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4076_ _0781_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4853__I _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5083__A1 dffram.data\[39\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3027_ _1482_ _2493_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3469__I _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input207_I sn76489_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _1678_ _1729_ _1731_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ dffram.data\[50\]\[1\] dffram.data\[51\]\[1\] _0775_ _0877_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6648_ _0605_ clknet_4_5_0_wb_clk_i dffram.data\[61\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4897__A1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6579_ _0536_ clknet_leaf_121_wb_clk_i wb_rst_override vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output259_I net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3321__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5074__A1 _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3388__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_153_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_153_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5065__A1 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ net252 net440 _2385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4901_ _1664_ _1524_ _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _1473_ _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _1504_ _1633_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_8_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3379__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ dffram.data\[59\]\[1\] _1586_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4114__S _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4694_ dffram.data\[30\]\[7\] _1533_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6502_ _0459_ clknet_leaf_133_wb_clk_i net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3714_ dffram.data\[24\]\[0\] dffram.data\[25\]\[0\] _0662_ _0663_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6433_ _0390_ clknet_4_6_0_wb_clk_i dffram.data\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3645_ _2921_ _2969_ _2971_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3576_ _1448_ _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6364_ _0321_ clknet_leaf_96_wb_clk_i dffram.data\[43\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _1956_ _1649_ _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6295_ _0252_ clknet_leaf_100_wb_clk_i dffram.data\[47\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3752__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input157_I qcpu_sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1873_ _1909_ _1911_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xhold27 net494 net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold16 net474 net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 net495 net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5177_ dffram.data\[23\]\[2\] _1862_ _1865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold49 net515 net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5679__I _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4128_ _1069_ _1070_ _1071_ _1072_ _0765_ _0766_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_39_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I ay8913_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4059_ _0769_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5359__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_35_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4567__B1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__C2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3927__I _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3863__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3662__I design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3542__A1 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5295__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3430_ _0628_ net429 _2830_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3361_ _2614_ _2768_ _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6080_ _0037_ clknet_leaf_22_wb_clk_i dffram.data\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5100_ dffram.data\[24\]\[2\] _1805_ _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4089__A2 _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5031_ dffram.data\[49\]\[2\] _1764_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3292_ wb_counter\[4\] wb_counter\[5\] wb_counter\[6\] _2709_ _2719_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_100_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5038__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3948__S _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ net440 _2372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5864_ _1448_ _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4815_ _1553_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5795_ _2276_ _1859_ _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4013__A2 _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5210__A1 _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _1569_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_17_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _1525_ _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3628_ _2928_ _2956_ _2960_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5513__A2 _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6416_ _0373_ clknet_leaf_87_wb_clk_i dffram.data\[40\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _0304_ clknet_leaf_79_wb_clk_i dffram.data\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4578__I _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3559_ _2870_ _2909_ _2914_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6278_ _0235_ clknet_leaf_69_wb_clk_i dffram.data\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput117 qcpu_oeb[13] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5277__A1 _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput106 qcpu_do[3] net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput128 qcpu_oeb[23] net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput139 qcpu_oeb[3] net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5229_ dffram.data\[4\]\[3\] _1896_ _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3431__B wb_sram_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3515__A1 _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4476__C1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5112__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5440__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4600_ _1469_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5580_ _2133_ _1583_ _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4531_ _1413_ _1415_ net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__I _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4462_ net207 _1345_ _1277_ net109 net61 _1352_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_68_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3506__A1 _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _0158_ clknet_leaf_19_wb_clk_i dffram.data\[39\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3413_ _2765_ _2817_ _2818_ _2806_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4393_ net132 _1304_ _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3344_ wb_counter\[16\] _2761_ _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6132_ _0089_ clknet_leaf_170_wb_clk_i dffram.data\[55\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6063_ _0020_ clknet_leaf_26_wb_clk_i dffram.data\[58\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ net248 _2705_ _2706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5014_ _1752_ _1753_ _1755_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__I _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5916_ net257 _2357_ _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _2264_ _2304_ _2309_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5778_ dffram.data\[3\]\[3\] _2258_ _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input85_I qcpu_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4729_ _1476_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_75_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__I _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_150_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_134_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4212__S _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__A1 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3850__I _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3060_ _2506_ _2522_ _2488_ _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5661__A1 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__S1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5777__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _2214_ _2207_ _2215_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3962_ dffram.data\[16\]\[2\] dffram.data\[17\]\[2\] _0840_ _0909_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3893_ dffram.data\[16\]\[1\] dffram.data\[17\]\[1\] _0840_ _0841_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__I wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5632_ _2168_ _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5563_ _2068_ _2120_ _2123_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3727__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_130_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4514_ _1321_ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5494_ _1463_ _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4445_ _1349_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4376_ net126 _1268_ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_10_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6115_ _0072_ clknet_leaf_17_wb_clk_i dffram.data\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3327_ _2573_ wb_counter\[12\] _2738_ _2748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3760__I _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6046_ _0003_ clknet_leaf_7_wb_clk_i dffram.data\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3258_ _2689_ _2692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3189_ _2633_ _2634_ _2635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4591__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__C _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__I _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output289_I net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5891__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4207__S _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_178_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_178_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_107_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold93_I wbs_dat_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3709__B2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3709__A1 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__S _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _1005_ _1172_ _1067_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4161_ dffram.data\[10\]\[5\] dffram.data\[11\]\[5\] _0923_ _1105_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4676__I _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5634__A1 _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A2 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4092_ dffram.data\[20\]\[4\] dffram.data\[21\]\[4\] _0843_ _1037_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3112_ _2567_ _2568_ _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _2502_ _2504_ _2505_ _2507_ _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_78_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5300__I _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4117__S _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ _1697_ _1735_ _1740_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3945_ dffram.data\[40\]\[1\] dffram.data\[41\]\[1\] _0807_ _0893_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4296__S1 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3956__S _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5615_ dffram.data\[42\]\[2\] _2156_ _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3876_ _0661_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_27_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6595_ _0552_ clknet_leaf_39_wb_clk_i dffram.data\[35\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5546_ _2105_ _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input187_I sn76489_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5477_ _1984_ _2062_ _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_112_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__I _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4428_ net30 _1279_ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input48_I mc14500_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4359_ net119 _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3490__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6029_ net242 _2437_ _2444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3665__I design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6041__I net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3798__S0 _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5616__A1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__A2 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__I _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _0674_ _0676_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_56_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _2940_ _2975_ _2980_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3592_ _2936_ _2933_ _2937_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_75_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6380_ _0337_ clknet_leaf_97_wb_clk_i dffram.data\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5400_ _1821_ _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _1949_ _1964_ _1967_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5855__A1 _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _1892_ _1915_ _1920_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4213_ dffram.data\[10\]\[6\] dffram.data\[11\]\[6\] _0705_ _1156_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5193_ _1874_ _1875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4144_ _0688_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5607__A1 _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ dffram.data\[42\]\[3\] dffram.data\[43\]\[3\] _0954_ _1021_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3026_ net371 _2470_ _2486_ _2492_ _2493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_65_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input102_I qcpu_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4977_ dffram.data\[26\]\[0\] _1730_ _1731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3928_ dffram.data\[48\]\[1\] dffram.data\[49\]\[1\] _0875_ _0876_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _0604_ clknet_leaf_44_wb_clk_i dffram.data\[61\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3859_ dffram.data\[40\]\[0\] dffram.data\[41\]\[0\] _0807_ _0808_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4346__A1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6578_ _0535_ clknet_leaf_120_wb_clk_i wb_override_act vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5529_ _2082_ _2098_ _2101_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4649__A2 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output321_I net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3085__A1 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A1 net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold56_I wbs_dat_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5837__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__I _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_122_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5880_ _2331_ _2328_ _2332_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4900_ _1538_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _1632_ _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5785__I _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4762_ _1539_ _1585_ _1587_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__A1 dffram.data\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4693_ _1474_ _1532_ _1536_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_28_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _0458_ clknet_leaf_132_wb_clk_i net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3644_ dffram.data\[9\]\[0\] _2970_ _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6432_ _0389_ clknet_leaf_58_wb_clk_i dffram.data\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4879__A2 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _0320_ clknet_leaf_83_wb_clk_i dffram.data\[44\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3575_ _2921_ _2923_ _2925_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3000__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__S _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5314_ _1955_ _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6294_ _0251_ clknet_leaf_100_wb_clk_i dffram.data\[47\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5245_ dffram.data\[7\]\[0\] _1910_ _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4500__A1 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold17 net482 net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 net491 net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4500__B2 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5176_ _1808_ _1861_ _1864_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold39 net505 net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4127_ dffram.data\[38\]\[4\] dffram.data\[39\]\[4\] _0949_ _1072_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4058_ _0864_ _1003_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3067__A1 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _2475_ net212 _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4567__B2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output271_I net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output369_I net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput390 net390 wbs_dat_o[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_109_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3058__A1 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4215__S _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3853__I _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3360_ _2707_ _2775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3074__B _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3291_ _2708_ _2716_ _2717_ _2718_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5030_ _1746_ _1763_ _1766_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_49_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3049__A1 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A1 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _2367_ _2357_ net431 _2371_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_48_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5863_ _2316_ _2318_ _2320_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_62_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5794_ _1955_ _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4125__S _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4814_ _1619_ _1612_ _1620_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4745_ _1551_ _1570_ _1575_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4352__C _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3772__A2 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _1525_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6415_ _0372_ clknet_leaf_93_wb_clk_i dffram.data\[40\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3627_ dffram.data\[61\]\[2\] _2957_ _2960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _0303_ clknet_leaf_78_wb_clk_i dffram.data\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3558_ dffram.data\[29\]\[3\] _2910_ _2914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _0234_ clknet_leaf_74_wb_clk_i dffram.data\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput118 qcpu_oeb[14] net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_90_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3489_ _2868_ _2863_ _2869_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput107 qcpu_do[4] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input30_I blinker_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput129 qcpu_oeb[24] net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5228_ _1880_ _1895_ _1899_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4594__I _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5159_ dffram.data\[51\]\[4\] _1852_ _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4960__A1 _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__I _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3451__A1 _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3848__I _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ net49 _1414_ _1408_ net16 _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_124_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4951__A1 _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4461_ net178 _1348_ _1350_ net25 _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_40_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6200_ _0157_ clknet_leaf_20_wb_clk_i dffram.data\[39\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3412_ net243 _2814_ _2818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4392_ _1303_ _1306_ net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6131_ _0088_ clknet_leaf_6_wb_clk_i dffram.data\[56\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3343_ _2757_ _2756_ _2753_ _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6062_ _0019_ clknet_leaf_26_wb_clk_i dffram.data\[58\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ _2704_ _2705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ dffram.data\[53\]\[4\] _1754_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3758__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5915_ net440 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5846_ dffram.data\[38\]\[3\] _2305_ _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5777_ _2073_ _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _1278_ _2458_ _2460_ _2454_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3745__A2 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _1562_ _1555_ _1563_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I mc14500_sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ dffram.data\[58\]\[2\] _1512_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3493__I _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _0286_ clknet_leaf_105_wb_clk_i dffram.data\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3681__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3433__A1 net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3984__A2 _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__A1 _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _0769_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5700_ dffram.data\[11\]\[7\] _2208_ _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3892_ _0739_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ _2168_ _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_42_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5562_ dffram.data\[44\]\[1\] _2121_ _2123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3727__A2 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4513_ _1400_ _1401_ net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5493_ _2074_ _2064_ _2075_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _0649_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4375_ _1291_ _1295_ net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_1_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _0071_ clknet_leaf_18_wb_clk_i dffram.data\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3326_ _2732_ _2745_ _2746_ _2747_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6045_ _0002_ clknet_leaf_10_wb_clk_i dffram.data\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5101__A1 _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input132_I qcpu_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A3 _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3257_ _2690_ _2691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3188_ net270 _2627_ _2628_ _2634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5829_ dffram.data\[13\]\[4\] _2298_ _2299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__I _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output351_I net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6039__I _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5878__I _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4603__C2 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold86_I wbs_dat_i[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_147_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_147_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4022__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5331__A1 _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ dffram.data\[8\]\[5\] dffram.data\[9\]\[5\] _0703_ _1104_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3111_ net258 _2553_ _2557_ _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4091_ dffram.data\[18\]\[4\] dffram.data\[19\]\[4\] _0972_ _1036_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3645__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3042_ _2506_ wb_counter\[2\] _2484_ _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4993_ dffram.data\[26\]\[7\] _1736_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3944_ _0886_ _0891_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3875_ _0695_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _2138_ _2155_ _2158_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4133__S _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6594_ _0551_ clknet_leaf_36_wb_clk_i dffram.data\[35\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _2074_ _2106_ _2111_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5476_ _1438_ _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ net194 _1333_ _1325_ net45 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4867__I _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4358_ _1257_ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4289_ dffram.data\[54\]\[7\] dffram.data\[55\]\[7\] _1200_ _1231_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3309_ net254 _2721_ _2734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3636__A1 _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6028_ net276 _2433_ _2443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output399_I net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5561__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3798__S1 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4364__A2 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3882__S _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4116__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_142_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ dffram.data\[9\]\[7\] _2976_ _2980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3591_ dffram.data\[60\]\[5\] _2934_ _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3792__S _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__A2 _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5330_ dffram.data\[8\]\[5\] _1965_ _1967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5261_ dffram.data\[7\]\[7\] _1916_ _1920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4687__I _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4212_ dffram.data\[8\]\[6\] dffram.data\[9\]\[6\] _0703_ _1155_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_44_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4512__C1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5192_ _1830_ _1509_ _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4143_ dffram.data\[30\]\[5\] dffram.data\[31\]\[5\] _0904_ _1087_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4074_ dffram.data\[40\]\[3\] dffram.data\[41\]\[3\] _0807_ _1020_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _2487_ _2489_ _2491_ _2492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_65_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4976_ _1728_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3766__I _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3927_ _0771_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_132_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _0603_ clknet_leaf_44_wb_clk_i dffram.data\[61\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3858_ _0771_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__A1 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3789_ dffram.data\[10\]\[0\] dffram.data\[11\]\[0\] _0737_ _0738_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _0534_ clknet_leaf_149_wb_clk_i wb_counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5528_ dffram.data\[10\]\[5\] _2099_ _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input60_I mc14500_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _2003_ _2048_ _2051_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A3 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3609__A1 _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output314_I net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4038__S _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__S _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5837__A2 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _1631_ _1437_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_162_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_162_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5773__A1 _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ dffram.data\[59\]\[0\] _1586_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4692_ dffram.data\[30\]\[6\] _1533_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6500_ _0457_ clknet_leaf_136_wb_clk_i net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3643_ _2968_ _2970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6431_ _0388_ clknet_leaf_66_wb_clk_i dffram.data\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6362_ _0319_ clknet_leaf_89_wb_clk_i dffram.data\[44\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3574_ dffram.data\[60\]\[0\] _2924_ _2925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5313_ _1484_ _1053_ _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6293_ _0250_ clknet_leaf_102_wb_clk_i dffram.data\[47\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ _1908_ _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5175_ dffram.data\[23\]\[1\] _1862_ _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold29 net488 net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold18 _2354_ net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4126_ dffram.data\[36\]\[4\] dffram.data\[37\]\[4\] _0759_ _1071_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0997_ _0999_ _1000_ _1002_ _0871_ _0872_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_79_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3067__A2 _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3008_ _2474_ _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4880__I _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_130_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__A1 _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4959_ dffram.data\[27\]\[2\] _1716_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _0586_ clknet_leaf_45_wb_clk_i dffram.data\[60\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output264_I net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput380 net380 wbs_dat_o[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput391 net391 wbs_dat_o[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_126_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__A2 _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__I _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__A2 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5507__A1 _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5126__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4030__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3290_ _2700_ _2718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _2370_ _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5994__A1 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5862_ dffram.data\[14\]\[0\] _2319_ _2320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5793_ _2274_ _2267_ _2275_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4813_ dffram.data\[6\]\[3\] _1613_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4744_ dffram.data\[37\]\[3\] _1571_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4675_ _1486_ _1524_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _0371_ clknet_leaf_93_wb_clk_i dffram.data\[40\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3626_ _2926_ _2956_ _2959_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6345_ _0302_ clknet_leaf_78_wb_clk_i dffram.data\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3557_ _2868_ _2909_ _2913_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6276_ _0233_ clknet_leaf_69_wb_clk_i dffram.data\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input162_I sid_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3488_ dffram.data\[34\]\[2\] _2864_ _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5227_ dffram.data\[4\]\[2\] _1896_ _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput108 qcpu_do[5] net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput119 qcpu_oeb[15] net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input23_I ay8913_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _1844_ _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4109_ _0921_ _1052_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5089_ _1727_ _1649_ _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__A1 _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4476__B2 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A1 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4779__A2 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5976__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4226__S _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4251__I1 dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__I _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _1360_ _1362_ net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4003__I1 dffram.data\[39\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4391_ net131 _1304_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3411_ _2670_ _2816_ _2817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6130_ _0087_ clknet_leaf_6_wb_clk_i dffram.data\[56\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3342_ _2752_ _2759_ _2760_ _2747_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4467__A1 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6061_ _0018_ clknet_leaf_28_wb_clk_i dffram.data\[58\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3273_ _2689_ _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4467__B2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5012_ _1742_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3690__A2 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5967__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5914_ _2355_ _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5845_ _2262_ _2304_ _2308_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5776_ _2262_ _2257_ _2263_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ net245 _2459_ _2460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4727_ dffram.data\[2\]\[6\] _1556_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ _1449_ _1511_ _1514_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_75_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3609_ _2930_ _2943_ _2948_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput90 qcpu_do[19] net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4589_ dffram.data\[5\]\[3\] _1445_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6328_ _0285_ clknet_leaf_105_wb_clk_i dffram.data\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6259_ _0216_ clknet_leaf_114_wb_clk_i dffram.data\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3014__I net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4046__S _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3433__A2 _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A1 _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3885__S _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _0823_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_69_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4621__A1 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ _0823_ _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _2104_ _2167_ _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3188__A1 net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5561_ _2061_ _2120_ _2122_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_42_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5492_ dffram.data\[45\]\[3\] _2065_ _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4512_ net171 _1396_ _1359_ net44 net11 _1393_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_81_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _1330_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_44_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4374_ net125 _1294_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_95_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6113_ _0070_ clknet_leaf_17_wb_clk_i dffram.data\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3325_ _2700_ _2747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6044_ _0001_ clknet_leaf_12_wb_clk_i dffram.data\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3256_ _2689_ _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3112__A1 _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4860__A1 _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3187_ _2619_ wb_counter\[21\] _2633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input125_I qcpu_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_53_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_85_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ _2290_ _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input90_I qcpu_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ dffram.data\[12\]\[5\] _2250_ _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4223__S0 _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__A1 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__B2 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold79_I wbs_dat_i[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_116_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3110_ _2534_ wb_counter\[10\] _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4090_ dffram.data\[16\]\[4\] dffram.data\[17\]\[4\] _0840_ _1035_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4973__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4842__A1 _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ _2481_ _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4992_ _1695_ _1735_ _1739_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _0887_ _0888_ _0889_ _0890_ _0801_ _0802_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3874_ _0822_ net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5613_ dffram.data\[42\]\[1\] _2156_ _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _0550_ clknet_leaf_36_wb_clk_i dffram.data\[35\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ dffram.data\[18\]\[3\] _2107_ _2111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _2060_ _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3581__A1 _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ _1320_ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4357_ _1282_ _1283_ net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__5086__A1 _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4288_ dffram.data\[52\]\[7\] dffram.data\[53\]\[7\] _0660_ _1230_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3308_ wb_counter\[9\] _2727_ _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_87_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3239_ _2663_ wb_counter\[29\] _2677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6027_ _2439_ _2440_ _2442_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output294_I net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3324__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__I _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_109_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3590_ _1469_ _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3563__A1 _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5260_ _1890_ _1915_ _1919_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4211_ _0792_ _1153_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_118_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _1801_ _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4142_ dffram.data\[28\]\[5\] dffram.data\[29\]\[5\] _0795_ _1086_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4073_ _0805_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4115__I0 _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_84_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3024_ _2490_ _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4291__A2 _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_82_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _1728_ _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_127_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3926_ _0864_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5240__A1 _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6645_ _0602_ clknet_leaf_40_wb_clk_i dffram.data\[61\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input192_I sn76489_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3788_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6576_ _0533_ clknet_leaf_135_wb_clk_i wb_counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5527_ _2077_ _2098_ _2100_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3554__A1 dffram.data\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input53_I mc14500_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5458_ dffram.data\[1\]\[1\] _2049_ _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4409_ _1276_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4649__A4 _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5389_ _1810_ _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5059__A1 _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4121__I3 _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output307_I net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3957__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__S _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__I _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5298__A1 _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5412__I _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3867__I _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _1584_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3711_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4691_ _1470_ _1532_ _1535_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3642_ _2968_ _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6430_ _0387_ clknet_leaf_66_wb_clk_i dffram.data\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_131_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_131_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_141_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _0318_ clknet_leaf_82_wb_clk_i dffram.data\[44\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__A1 _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3573_ _2922_ _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _1953_ _1946_ _1954_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _0249_ clknet_leaf_99_wb_clk_i dffram.data\[47\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5289__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5243_ _1908_ _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5174_ _1802_ _1861_ _1863_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4125_ dffram.data\[34\]\[4\] dffram.data\[35\]\[4\] _0946_ _1070_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3978__S _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4056_ dffram.data\[62\]\[3\] dffram.data\[63\]\[3\] _1001_ _1002_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5461__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3007_ net213 _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_78_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input205_I sn76489_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__A1 _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4958_ _1683_ _1715_ _1718_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3909_ dffram.data\[8\]\[1\] dffram.data\[9\]\[1\] _0734_ _0857_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4889_ _1619_ _1666_ _1671_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6628_ _0585_ clknet_leaf_5_wb_clk_i dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3527__A1 _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4401__I _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6559_ _0516_ clknet_leaf_153_wb_clk_i wb_counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_113_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output257_I net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput370 net370 wbs_ack_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput381 net381 wbs_dat_o[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput392 net392 wbs_dat_o[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A1 _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5930_ _1480_ _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _2317_ _2319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5792_ dffram.data\[3\]\[7\] _2268_ _2275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4812_ _1550_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4743_ _1548_ _1570_ _1574_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6413_ _0370_ clknet_leaf_93_wb_clk_i dffram.data\[40\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4674_ _1523_ _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3625_ dffram.data\[61\]\[1\] _2957_ _2959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6344_ _0301_ clknet_leaf_78_wb_clk_i dffram.data\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3556_ dffram.data\[29\]\[2\] _2910_ _2913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6275_ _0232_ clknet_leaf_113_wb_clk_i dffram.data\[48\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3780__I1 dffram.data\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input155_I qcpu_sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3487_ _1454_ _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5226_ _1878_ _1895_ _1898_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput109 qcpu_do[6] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5157_ _1844_ _1851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_108_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4108_ _0749_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5088_ _1801_ _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input16_I ay8913_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4891__I _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4039_ dffram.data\[6\]\[3\] dffram.data\[7\]\[3\] _0852_ _0985_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3748__A1 _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4079__I2 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4400__A2 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4390_ _1303_ _1305_ net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_0_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ _2802_ _2812_ _2794_ _2809_ _2816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_110_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3341_ net229 _2750_ _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__I _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3880__I _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I ay8913_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _0017_ clknet_leaf_28_wb_clk_i dffram.data\[58\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_72_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ wb_counter\[3\] _2702_ _2703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5011_ _1742_ _1753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5416__A1 _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ net213 _2350_ _2354_ _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5844_ dffram.data\[38\]\[2\] _2305_ _2308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ dffram.data\[3\]\[2\] _2258_ _2263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2987_ _2457_ _2459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ _1561_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4657_ dffram.data\[58\]\[1\] _1512_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3608_ dffram.data\[19\]\[3\] _2944_ _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput91 qcpu_do[1] net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput80 qcpu_do[0] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4588_ _1459_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6327_ _0284_ clknet_leaf_127_wb_clk_i dffram.data\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__I _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3539_ _2895_ _2902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5655__A1 _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ _0215_ clknet_leaf_114_wb_clk_i dffram.data\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5209_ dffram.data\[50\]\[4\] _1886_ _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6189_ _0146_ clknet_leaf_156_wb_clk_i dffram.data\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3681__A3 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__S _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4241__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5646__A1 _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4237__S _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4621__A2 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3890_ _0825_ _0830_ _0832_ _0833_ _0836_ _0837_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_128_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5560_ dffram.data\[44\]\[0\] _2121_ _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5491_ _2073_ _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_38_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ net193 _1385_ _1386_ net90 _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_123_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4442_ _1337_ _1328_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4373_ _1249_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6112_ _0069_ clknet_leaf_17_wb_clk_i dffram.data\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_70_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3324_ net226 _2721_ _2746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6043_ _0000_ clknet_leaf_10_wb_clk_i dffram.data\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3255_ _2471_ net256 _2548_ _2689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_1_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3186_ _2561_ _2632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input118_I qcpu_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4612__A2 _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3785__I _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5827_ _2290_ _2297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _2206_ _2249_ _2251_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3179__A2 wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ dffram.data\[2\]\[2\] _1542_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input83_I qcpu_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _2196_ _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_116_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4223__S1 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output337_I net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A1 _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6483__D _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3695__I design_select\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_156_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_156_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3040_ net405 _2479_ _2505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4991_ dffram.data\[26\]\[6\] _1736_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3942_ dffram.data\[38\]\[1\] dffram.data\[39\]\[1\] _0799_ _0890_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_67_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3873_ _0752_ _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5612_ _2132_ _2155_ _2157_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6592_ _0549_ clknet_leaf_34_wb_clk_i dffram.data\[35\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_80_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5543_ _2071_ _2106_ _2110_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5474_ _1442_ _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4425_ net172 _1330_ _1331_ net91 net12 _1318_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_2_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__A1 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__B2 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4356_ net118 _1272_ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_6_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3307_ _2707_ _2732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4287_ dffram.data\[50\]\[7\] dffram.data\[51\]\[7\] _1216_ _1229_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_87_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3238_ _2668_ _2676_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6026_ _2441_ _2442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3169_ net380 _2609_ _2602_ _2617_ _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output287_I net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold91_I wbs_dat_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3260__A1 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4512__A1 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ _1149_ _1150_ _1151_ _1152_ _0836_ _0986_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4512__B2 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1828_ _1867_ _1872_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4141_ dffram.data\[26\]\[5\] dffram.data\[27\]\[5\] _0964_ _1085_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4072_ _0886_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3079__A1 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3023_ _2352_ _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6017__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4974_ _1727_ _1509_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3925_ _0866_ _0867_ _0869_ _0870_ _0871_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__3251__A1 _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6644_ _0601_ clknet_leaf_73_wb_clk_i dffram.data\[19\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3856_ _0694_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3787_ _0701_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_15_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6575_ _0532_ clknet_leaf_136_wb_clk_i wb_counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5526_ dffram.data\[10\]\[4\] _2099_ _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4160__S _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4751__A1 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input185_I sn76489_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5457_ _1998_ _2048_ _2050_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4408_ _1315_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input46_I mc14500_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5388_ _2003_ _2000_ _2004_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4339_ _1269_ _1271_ net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6009_ net237 _2426_ _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__A1 net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4990__A1 _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3769__C1 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _0658_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_16_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ dffram.data\[30\]\[5\] _1533_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3641_ _2276_ _2167_ _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _0317_ clknet_leaf_82_wb_clk_i dffram.data\[44\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3572_ _2922_ _2923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ dffram.data\[48\]\[7\] _1947_ _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_171_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_171_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _0248_ clknet_leaf_112_wb_clk_i dffram.data\[21\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _1907_ _1859_ _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5173_ dffram.data\[23\]\[0\] _1862_ _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4124_ dffram.data\[32\]\[4\] dffram.data\[33\]\[4\] _0754_ _1069_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput1 ay8913_do[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4055_ _0761_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3006_ _2472_ _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4155__S _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input100_I qcpu_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4421__B1 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ dffram.data\[27\]\[1\] _1716_ _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3994__S _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3775__A2 _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3908_ _0725_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4972__A1 _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ dffram.data\[55\]\[3\] _1667_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3793__I _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _0584_ clknet_leaf_6_wb_clk_i dffram.data\[29\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3839_ _0773_ _0776_ _0780_ _0783_ _0785_ _0787_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_104_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _0515_ clknet_leaf_154_wb_clk_i wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_95_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _2087_ _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_112_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6489_ _0446_ clknet_leaf_145_wb_clk_i net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput360 net360 qcpu_sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput371 net371 wbs_dat_o[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput393 net393 wbs_dat_o[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput382 net382 wbs_dat_o[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3033__I _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3463__A1 _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4263__I0 _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3454__A1 dffram.data\[36\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _2317_ _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4811_ _1617_ _1612_ _1618_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _2087_ _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4742_ dffram.data\[37\]\[2\] _1571_ _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4673_ _1487_ _1507_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6412_ _0369_ clknet_leaf_92_wb_clk_i dffram.data\[40\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3624_ _2921_ _2956_ _2958_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__A1 _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6343_ _0300_ clknet_leaf_77_wb_clk_i dffram.data\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3555_ _2866_ _2909_ _2912_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3486_ _2866_ _2863_ _2867_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6274_ _0231_ clknet_leaf_113_wb_clk_i dffram.data\[48\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5225_ dffram.data\[4\]\[1\] _1896_ _1898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5131__A1 _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input148_I qcpu_sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1814_ _1845_ _1850_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4107_ _1048_ _1049_ _1050_ _1051_ _0928_ _0929_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_108_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5087_ _1442_ _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3445__A1 _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ dffram.data\[4\]\[3\] dffram.data\[5\]\[3\] _0983_ _0984_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3788__I _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5989_ net265 _2411_ _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4945__A1 _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5508__I _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output367_I net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5243__I _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3340_ _2756_ _2758_ _2759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1553_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_72_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3271_ wb_counter\[0\] _2496_ wb_counter\[2\] _2702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_108_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5912_ net214 _2353_ _2354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5843_ _2260_ _2304_ _2307_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__A1 dffram.data\[54\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5774_ _2070_ _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2986_ _2457_ _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4725_ _1472_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _1444_ _1511_ _1513_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput70 mc14500_sram_addr[5] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3607_ _2928_ _2943_ _2947_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5352__A1 _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1458_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput81 qcpu_do[10] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6651__CLK clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3538_ _2870_ _2896_ _2901_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6326_ _0283_ clknet_leaf_129_wb_clk_i dffram.data\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput92 qcpu_do[20] net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3469_ _2848_ _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6257_ _0214_ clknet_leaf_115_wb_clk_i dffram.data\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5208_ _1874_ _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6188_ _0145_ clknet_leaf_163_wb_clk_i dffram.data\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5139_ _1817_ _1838_ _1840_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_4_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_101_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A2 _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3981__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3657__A1 _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__B _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4082__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4253__S _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__A2 _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__I _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5490_ _1458_ _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4510_ _1398_ _1399_ net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_0_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4441_ _1340_ _1343_ _1346_ net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_79_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4372_ _1291_ _1293_ net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_0_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6111_ _0068_ clknet_leaf_170_wb_clk_i dffram.data\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3323_ wb_counter\[12\] _2742_ _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3254_ _2371_ _2351_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6042_ net281 _2376_ _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3185_ _2624_ _2631_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5826_ _2264_ _2291_ _2296_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A1 _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5757_ dffram.data\[12\]\[4\] _2250_ _2251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _1547_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input76_I mc14500_sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _2076_ _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5325__A1 _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4639_ dffram.data\[31\]\[5\] _1498_ _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6309_ _0266_ clknet_leaf_128_wb_clk_i dffram.data\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3041__I _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3976__I _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4600__I _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4248__S _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_125_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _1693_ _1735_ _1738_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3941_ dffram.data\[36\]\[1\] dffram.data\[37\]\[1\] _0797_ _0889_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6660_ _0617_ clknet_leaf_74_wb_clk_i dffram.data\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3872_ _0768_ _0791_ _0804_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_144_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A1 _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ dffram.data\[42\]\[0\] _2156_ _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6591_ _0548_ clknet_leaf_35_wb_clk_i dffram.data\[35\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5542_ dffram.data\[18\]\[2\] _2107_ _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5473_ _2017_ _2054_ _2059_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4424_ _1276_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _1281_ _1282_ net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_10_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3126__I _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout405 net279 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_111_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3306_ _2729_ _2731_ _2451_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4286_ dffram.data\[48\]\[7\] dffram.data\[49\]\[7\] _1200_ _1228_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input130_I qcpu_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6025_ _2362_ _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3237_ net391 _2654_ _2669_ _2675_ _2676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_87_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3168_ _2615_ _2616_ _2617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3099_ net287 _2553_ _2557_ _2558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_25_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3796__I _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4597__A2 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5809_ _2266_ _2284_ _2286_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__C1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4068__S _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3260__A2 _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4140_ dffram.data\[24\]\[5\] dffram.data\[25\]\[5\] _0671_ _1084_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4115__I2 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _1013_ _1014_ _1015_ _1016_ _0801_ _0802_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__3079__A2 _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3022_ _2488_ _2489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5776__A1 _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4973_ _1485_ _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3924_ _0745_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6643_ _0600_ clknet_leaf_84_wb_clk_i dffram.data\[19\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3855_ _0792_ _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3786_ dffram.data\[8\]\[0\] dffram.data\[9\]\[0\] _0734_ _0735_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _0531_ clknet_leaf_134_wb_clk_i wb_counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5525_ _2091_ _2099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_22_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input178_I sid_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5456_ dffram.data\[1\]\[0\] _2049_ _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4407_ _0620_ _0635_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ dffram.data\[20\]\[1\] _2001_ _2004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4338_ _1253_ _1270_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input39_I mc14500_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ dffram.data\[6\]\[7\] dffram.data\[7\]\[7\] _1209_ _1211_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6008_ net271 _2422_ _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5519__A1 _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3242__A2 _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output397_I net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5758__A1 _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4325__I _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3769__C2 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _2940_ _2962_ _2967_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4261__S _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3571_ _1647_ _2118_ _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4733__A2 _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _0247_ clknet_leaf_112_wb_clk_i dffram.data\[21\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5310_ _1827_ _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__I _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ _1430_ _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4497__B2 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5172_ _1860_ _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ _1005_ _1066_ _1067_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput2 ay8913_do[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4054_ dffram.data\[60\]\[3\] dffram.data\[61\]\[3\] _0868_ _1000_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__A1 net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3005_ _2471_ _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4421__A1 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4421__B2 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4956_ _1678_ _1715_ _1717_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_35_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3907_ _0848_ _0850_ _0851_ _0853_ _0854_ _0690_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4887_ _1617_ _1666_ _1670_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3838_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6626_ _0583_ clknet_4_0_0_wb_clk_i dffram.data\[29\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6557_ _0514_ clknet_leaf_152_wb_clk_i wb_counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5508_ _1476_ _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3769_ net221 _0717_ _0640_ net151 _0643_ net70 _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_70_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ _0445_ clknet_leaf_144_wb_clk_i net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput350 net350 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput361 net361 qcpu_sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ dffram.data\[46\]\[2\] _2036_ _2039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_58_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput372 net372 wbs_dat_o[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput383 net383 wbs_dat_o[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput394 net394 wbs_dat_o[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4660__A1 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output312_I net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_97_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4145__I _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4263__I1 _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5704__I _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__S0 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5979__A1 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4055__I _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4810_ dffram.data\[6\]\[2\] _1613_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5790_ _2272_ _2267_ _2273_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _1545_ _1570_ _1573_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4672_ _1478_ _1517_ _1522_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _0368_ clknet_leaf_83_wb_clk_i dffram.data\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3623_ dffram.data\[61\]\[0\] _2957_ _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5903__A1 _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6342_ _0299_ clknet_leaf_54_wb_clk_i dffram.data\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3554_ dffram.data\[29\]\[1\] _2910_ _2912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ dffram.data\[34\]\[1\] _2864_ _2867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6273_ _0230_ clknet_leaf_113_wb_clk_i dffram.data\[48\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_90_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5224_ _1873_ _1895_ _1897_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5155_ dffram.data\[51\]\[3\] _1846_ _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4106_ dffram.data\[14\]\[4\] dffram.data\[15\]\[4\] _0926_ _1051_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5086_ _1760_ _1795_ _1800_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4037_ _0665_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4642__A1 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input210_I sn76489_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5988_ _2412_ _2413_ _2408_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4939_ _1685_ _1702_ _1706_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6609_ _0566_ clknet_leaf_3_wb_clk_i dffram.data\[33\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__I _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output262_I net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3979__I _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5434__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3270_ _2691_ _2698_ _2699_ _2701_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_72_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__A1 _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3889__I _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ net215 _2352_ _2353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5842_ dffram.data\[38\]\[1\] _2305_ _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5773_ _2260_ _2257_ _2261_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5609__I _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _1559_ _1555_ _1560_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2985_ _2455_ _2350_ _2456_ _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4655_ dffram.data\[58\]\[0\] _1512_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput71 mc14500_sram_gwe net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3606_ dffram.data\[19\]\[2\] _2944_ _2947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4586_ net248 _1451_ _1457_ net156 _1452_ net75 _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_115_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput60 mc14500_do[5] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput82 qcpu_do[11] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3537_ dffram.data\[32\]\[3\] _2897_ _2901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6325_ _0282_ clknet_leaf_127_wb_clk_i dffram.data\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3363__A1 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput93 qcpu_do[21] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input160_I qcpu_sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3468_ _2848_ _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6256_ _0213_ clknet_leaf_115_wb_clk_i dffram.data\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _0144_ clknet_leaf_115_wb_clk_i dffram.data\[49\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5207_ _1874_ _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3399_ net241 _2730_ _2807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input21_I ay8913_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ dffram.data\[52\]\[4\] _1839_ _1840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_4_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5069_ dffram.data\[39\]\[0\] _1790_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3354__A1 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__I _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3106__A1 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ net174 _1344_ _1345_ net203 net21 _1318_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_80_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__B1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3345__A1 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ net123 _1284_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6110_ _0067_ clknet_leaf_169_wb_clk_i dffram.data\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3322_ _2743_ _2744_ _2451_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6041_ net247 _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3253_ _2668_ _2688_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_13_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3184_ net383 _2609_ _2625_ _2630_ _2631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_105_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5825_ dffram.data\[13\]\[3\] _2292_ _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _2242_ _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5687_ _2204_ _2197_ _2205_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3584__A1 _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4707_ _1453_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_20_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _1465_ _1497_ _1499_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input69_I mc14500_sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4569_ _1443_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5089__A1 _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _0265_ clknet_leaf_128_wb_clk_i dffram.data\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6239_ _0196_ clknet_leaf_129_wb_clk_i dffram.data\[50\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4836__A1 _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_40_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3575__A1 _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput250 net434 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3940_ dffram.data\[34\]\[1\] dffram.data\[35\]\[1\] _0795_ _0888_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5252__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3802__A2 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _0806_ _0817_ _0819_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_165_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_165_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5610_ _2154_ _2156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6590_ _0547_ clknet_leaf_35_wb_clk_i dffram.data\[35\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5541_ _2068_ _2106_ _2109_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ dffram.data\[1\]\[7\] _2055_ _2059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4423_ _1315_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _0626_ _0652_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_6_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3305_ net253 _2730_ _2731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4285_ _0805_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6024_ net241 _2437_ _2440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3236_ _2671_ _2674_ _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3167_ net266 _2604_ _2605_ _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input123_I qcpu_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3098_ _2556_ _2557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4174__S _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2981__I _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__C1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5808_ dffram.data\[15\]\[4\] _2285_ _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5739_ _2210_ _2236_ _2239_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3557__A1 _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3309__A1 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6514__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4285__A2 _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A1 _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__S _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3548__A1 _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold77_I wbs_dat_i[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__S _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4070_ dffram.data\[38\]\[3\] dffram.data\[39\]\[3\] _0949_ _1016_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5473__A1 _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3021_ _2455_ _2488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4972_ _1697_ _1721_ _1726_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3923_ _0764_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6642_ _0599_ clknet_leaf_73_wb_clk_i dffram.data\[19\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3854_ _0794_ _0796_ _0798_ _0800_ _0801_ _0802_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4521__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3785_ _0702_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6573_ _0530_ clknet_leaf_136_wb_clk_i wb_counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5524_ _2091_ _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_113_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _2047_ _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_62_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ _1290_ _1314_ net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_93_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5386_ _1807_ _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4169__S _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _0638_ _0651_ net405 _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_105_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4268_ dffram.data\[4\]\[7\] dffram.data\[5\]\[7\] _1209_ _1210_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6007_ _2425_ _2427_ _2419_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3219_ net275 _2649_ _2650_ _2660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4199_ _0696_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__A1 _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output292_I net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3769__A1 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3769__B2 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _1443_ _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1892_ _1901_ _1906_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__I _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5171_ _1860_ _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4122_ _0789_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5446__A1 _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4053_ dffram.data\[58\]\[3\] dffram.data\[59\]\[3\] _0998_ _0999_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 ay8913_do[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3004_ net214 _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4955_ dffram.data\[27\]\[0\] _1716_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3906_ _0835_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ dffram.data\[55\]\[2\] _1667_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3837_ _0687_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5347__I _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _0582_ clknet_leaf_7_wb_clk_i dffram.data\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3768_ _0657_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input190_I sn76489_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0513_ clknet_leaf_151_wb_clk_i wb_counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _2085_ _2078_ _2086_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3699_ _0649_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6487_ _0444_ clknet_leaf_147_wb_clk_i net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput340 net340 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput351 net351 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput362 net362 qcpu_sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input51_I mc14500_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ _2003_ _2035_ _2038_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5369_ _1943_ _1986_ _1991_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput373 net373 wbs_dat_o[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput384 net384 wbs_dat_o[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput395 net395 wbs_dat_o[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_126_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4426__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output305_I net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4023__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3782__S0 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_169_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4272__S _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4740_ dffram.data\[37\]\[1\] _1571_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4671_ dffram.data\[58\]\[7\] _1518_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6410_ _0367_ clknet_leaf_85_wb_clk_i dffram.data\[16\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3622_ _2955_ _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _0298_ clknet_leaf_77_wb_clk_i dffram.data\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _2861_ _2909_ _2911_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3484_ _1448_ _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6272_ _0229_ clknet_leaf_118_wb_clk_i dffram.data\[48\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5667__A1 _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ dffram.data\[4\]\[0\] _1896_ _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5154_ _1811_ _1845_ _1849_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4105_ dffram.data\[12\]\[4\] dffram.data\[13\]\[4\] _0991_ _1050_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_108_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5085_ dffram.data\[39\]\[7\] _1796_ _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4036_ dffram.data\[2\]\[3\] dffram.data\[3\]\[3\] _0849_ _0982_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input203_I sn76489_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5987_ net230 _2404_ _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4938_ dffram.data\[28\]\[2\] _1703_ _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5077__I _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ dffram.data\[56\]\[4\] _1658_ _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input99_I qcpu_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _0565_ clknet_leaf_30_wb_clk_i dffram.data\[33\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6539_ _0496_ clknet_leaf_137_wb_clk_i net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5830__A1 _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5897__A1 _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4624__A2 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ net255 net222 _2351_ _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_115_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5841_ _2255_ _2304_ _2306_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ dffram.data\[3\]\[1\] _2258_ _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2984_ wb_feedback_delay _1483_ _2456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4723_ dffram.data\[2\]\[5\] _1556_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4654_ _1510_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput72 mc14500_sram_in[0] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput50 mc14500_do[24] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3605_ _2926_ _2943_ _2946_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4585_ _0641_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput61 mc14500_do[6] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4560__B2 _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4560__A1 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3536_ _2868_ _2896_ _2900_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6324_ _0281_ clknet_leaf_129_wb_clk_i dffram.data\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput83 qcpu_do[12] net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput94 qcpu_do[22] net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_110_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6255_ _0212_ clknet_leaf_164_wb_clk_i dffram.data\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input153_I qcpu_sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3467_ _2325_ _2849_ _2854_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5206_ _1816_ _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6186_ _0143_ clknet_leaf_114_wb_clk_i dffram.data\[49\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3398_ _2792_ _2804_ _2805_ _2806_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5360__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ _1831_ _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5068_ _1788_ _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input14_I ay8913_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ dffram.data\[26\]\[3\] dffram.data\[27\]\[3\] _0964_ _0965_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4171__S0 _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4379__A1 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4704__I _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_134_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3354__A2 _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4087__S _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A1 _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4614__I _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__B2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4370_ _1291_ _1292_ net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_74_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3321_ net225 _2730_ _2744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3252_ net395 _2491_ _2669_ _2687_ _2688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6040_ _2449_ _2450_ _2451_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input6_I ay8913_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _2626_ _2629_ _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_87_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3281__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5824_ _2262_ _2291_ _2295_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _2242_ _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5686_ dffram.data\[11\]\[3\] _2198_ _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ _1545_ _1541_ _1546_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ dffram.data\[31\]\[4\] _1498_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4533__A1 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__B2 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ net404 _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_102_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1390_ _1391_ net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _0264_ clknet_leaf_109_wb_clk_i dffram.data\[20\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3519_ _2882_ _2890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5089__A2 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _0195_ clknet_leaf_129_wb_clk_i dffram.data\[50\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6169_ _0126_ clknet_leaf_171_wb_clk_i dffram.data\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6038__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__A1 _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A1 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__I _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__B2 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_56_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3714__S _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4127__I1 dffram.data\[39\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4609__I _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput251 net433 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput240 net456 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6029__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3263__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3870_ _0818_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5540_ dffram.data\[18\]\[1\] _2107_ _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4280__S _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _2015_ _2054_ _2058_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4422_ _1319_ _1329_ net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_134_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4353_ net117 _1268_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4284_ _1222_ _1223_ _1224_ _1225_ _1196_ _0714_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_6_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3304_ _2726_ _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_111_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6023_ net275 _2433_ _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3235_ net277 _2672_ _2673_ _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3166_ _2596_ _2614_ _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3097_ _2555_ _2556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input116_I qcpu_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__C2 _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3254__A1 _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5807_ _2277_ _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3999_ _0756_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ dffram.data\[40\]\[5\] _2237_ _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I qcpu_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_131_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__A1 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _2150_ _2188_ _2192_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4506__B2 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output335_I net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_142_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3245__A1 net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3508__I _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3020_ wb_override_act _2487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4275__S _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4971_ dffram.data\[27\]\[7\] _1722_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ dffram.data\[62\]\[1\] dffram.data\[63\]\[1\] _0762_ _0870_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_82_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4984__A1 _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6641_ _0598_ clknet_leaf_84_wb_clk_i dffram.data\[19\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ _0689_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4802__I _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _0695_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6572_ _0529_ clknet_leaf_148_wb_clk_i wb_counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5523_ _2074_ _2092_ _2097_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5454_ _2047_ _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _0637_ net138 _1312_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_100_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5385_ _1998_ _2000_ _2002_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4336_ net144 _1268_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4267_ _0826_ _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_leaf_31_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4198_ _1137_ _1138_ _1139_ _1140_ _0968_ _1089_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6006_ net236 _2426_ _2427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3218_ _2641_ wb_counter\[26\] _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__S _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3149_ _2578_ _2600_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4712__I _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output285_I net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3950__A2 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A1 _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3769__A2 _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A1 _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4430__A3 _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5143__A1 _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5170_ _1858_ _1859_ _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _1062_ _1063_ _1064_ _1065_ _0881_ _0883_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__3457__A1 _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _0756_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput4 ay8913_do[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3003_ _2469_ _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4954_ _1714_ _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ dffram.data\[6\]\[1\] dffram.data\[7\]\[1\] _0852_ _0853_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4885_ _1615_ _1666_ _1669_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3836_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_6_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _0581_ clknet_leaf_178_wb_clk_i dffram.data\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3767_ _0704_ _0706_ _0710_ _0712_ _0713_ _0715_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_7_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6555_ _0512_ clknet_leaf_154_wb_clk_i wb_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5506_ dffram.data\[45\]\[6\] _2079_ _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input183_I sn76489_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ _0634_ _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6486_ _0443_ clknet_leaf_144_wb_clk_i net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput341 net341 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput330 net330 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput352 net352 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ dffram.data\[46\]\[1\] _2036_ _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput363 net363 rst_ay8913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input44_I mc14500_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ dffram.data\[47\]\[3\] _1987_ _1991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput396 net396 wbs_dat_o[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput374 net374 wbs_dat_o[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput385 net385 wbs_dat_o[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4319_ net124 _1258_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5299_ _1816_ _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_410 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_126_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4707__I _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A3 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3620__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3439__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4939__A1 _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _1474_ _1517_ _1521_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3621_ _2955_ _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _0297_ clknet_leaf_54_wb_clk_i dffram.data\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3914__A2 _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3552_ dffram.data\[29\]\[0\] _2910_ _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_133_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ _2861_ _2863_ _2865_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6271_ _0228_ clknet_leaf_119_wb_clk_i dffram.data\[48\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ _1894_ _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5153_ dffram.data\[51\]\[2\] _1846_ _1849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4104_ dffram.data\[10\]\[4\] dffram.data\[11\]\[4\] _0923_ _1049_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5084_ _1758_ _1795_ _1799_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_142_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4035_ dffram.data\[0\]\[3\] dffram.data\[1\]\[3\] _0980_ _0981_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5986_ net264 _2411_ _2412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4937_ _1683_ _1702_ _1705_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4868_ _1650_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3819_ _0696_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6607_ _0564_ clknet_leaf_31_wb_clk_i dffram.data\[33\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _1565_ _1604_ _1609_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6538_ _0495_ clknet_leaf_137_wb_clk_i net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _0426_ clknet_leaf_42_wb_clk_i dffram.data\[62\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4397__A2 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4900__I _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4283__S _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ dffram.data\[38\]\[0\] _2305_ _2306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5771_ _2067_ _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ net215 _2455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4722_ _1558_ _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput40 mc14500_do[15] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4653_ _1510_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput73 mc14500_sram_in[1] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput51 mc14500_do[25] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3604_ dffram.data\[19\]\[1\] _2944_ _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput62 mc14500_do[7] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4584_ _1441_ _1455_ _1456_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6323_ _0280_ clknet_leaf_99_wb_clk_i dffram.data\[46\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4560__A2 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3535_ dffram.data\[32\]\[2\] _2897_ _2900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput84 qcpu_do[13] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput95 qcpu_do[23] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3466_ dffram.data\[35\]\[3\] _2850_ _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6254_ _0211_ clknet_leaf_164_wb_clk_i dffram.data\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1882_ _1875_ _1883_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__I _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _0142_ clknet_leaf_114_wb_clk_i dffram.data\[49\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3397_ _2370_ _2806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5136_ _1831_ _1838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input146_I qcpu_sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _1788_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4018_ _0661_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4171__S1 _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5088__I _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2355_ _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3051__A2 _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output365_I net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4303__A2 _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5319__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3320_ _2693_ _2741_ _2742_ _2743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3251_ _2685_ _2686_ _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3182_ net269 _2627_ _2628_ _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3910__S _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5823_ dffram.data\[13\]\[2\] _2292_ _2295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5754_ _2204_ _2243_ _2248_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5685_ _2073_ _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4705_ dffram.data\[2\]\[1\] _1542_ _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _1490_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4567_ net223 _1312_ _0642_ net153 _0645_ net72 _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_6306_ _0263_ clknet_leaf_110_wb_clk_i dffram.data\[20\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4498_ net167 _1383_ _1388_ net40 net7 _1379_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_3518_ _2882_ _2889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3449_ _2327_ _2841_ _2843_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4188__S _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _0194_ clknet_leaf_129_wb_clk_i dffram.data\[50\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6168_ _0125_ clknet_leaf_171_wb_clk_i dffram.data\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5119_ _1825_ _1818_ _1826_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6099_ _0056_ clknet_4_1_0_wb_clk_i dffram.data\[59\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__I _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5549__A1 _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4509__C1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__I _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput241 net454 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput230 net447 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput252 net464 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_hold15_I wbs_dat_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4625__I _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3263__A2 _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5470_ dffram.data\[1\]\[6\] _2055_ _2058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ net183 _1322_ _1325_ net34 _1328_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5712__A1 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3905__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4352_ net405 _0638_ _1280_ _0635_ net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xclkbuf_leaf_174_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_174_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_111_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4283_ dffram.data\[62\]\[7\] dffram.data\[63\]\[7\] _1194_ _1225_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5191__I _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3303_ _2725_ _2728_ _2729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6022_ _2436_ _2438_ _2430_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3234_ _2555_ _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3165_ wb_counter\[18\] _2614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5779__A1 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3096_ _2471_ _2554_ _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_25_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4451__B2 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__A1 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input109_I qcpu_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5806_ _2277_ _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ dffram.data\[32\]\[2\] dffram.data\[33\]\[2\] _0793_ _0945_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5737_ _2206_ _2236_ _2238_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5951__A1 _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input74_I mc14500_sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5668_ dffram.data\[41\]\[6\] _2189_ _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5599_ _2081_ _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ _1484_ _1040_ _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_40_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output328_I net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_149_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4445__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5942__A1 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_51_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4681__A1 _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1695_ _1721_ _1725_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ dffram.data\[60\]\[1\] dffram.data\[61\]\[1\] _0868_ _0869_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _0597_ clknet_leaf_76_wb_clk_i dffram.data\[19\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ _0764_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6571_ _0528_ clknet_leaf_136_wb_clk_i wb_counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5522_ dffram.data\[10\]\[3\] _2093_ _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3783_ _0725_ _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5453_ _1907_ _1633_ _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4404_ _1302_ _1313_ net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5384_ dffram.data\[20\]\[0\] _2001_ _2002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4335_ _1249_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6433__CLK clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4266_ dffram.data\[2\]\[7\] dffram.data\[3\]\[7\] _1189_ _1208_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4672__A1 _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4197_ dffram.data\[30\]\[6\] dffram.data\[31\]\[6\] _0728_ _1140_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6005_ _2390_ _2426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3217_ _2646_ _2658_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3148_ net377 _2587_ _2579_ _2599_ _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_124_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4275__I1 dffram.data\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3079_ net399 _2518_ _2538_ _2539_ _2540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_49_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__A1 net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3786__I0 dffram.data\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_28_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output278_I net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_144_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_37_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4266__I1 dffram.data\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4903__I _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold82_I wbs_dat_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3519__I _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_46_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5734__I _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ dffram.data\[54\]\[4\] dffram.data\[55\]\[4\] _0779_ _1065_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4286__S _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4051_ dffram.data\[56\]\[3\] dffram.data\[57\]\[3\] _0865_ _0997_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 ay8913_do[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3457__A2 _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3002_ _2352_ _2469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4406__A1 _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _1714_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _0668_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6623_ _0580_ clknet_leaf_177_wb_clk_i dffram.data\[29\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4884_ dffram.data\[55\]\[1\] _1667_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ _0680_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3766_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6554_ _0511_ clknet_leaf_150_wb_clk_i wb_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _2084_ _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6485_ _0442_ clknet_leaf_132_wb_clk_i net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3697_ _0647_ _0619_ _0625_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5436_ _1998_ _2035_ _2037_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input176_I sid_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput331 net331 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput342 net342 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput353 net353 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput320 net320 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput364 net364 rst_blinker vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5367_ _1941_ _1986_ _1990_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4893__A1 _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput375 net375 wbs_dat_o[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput386 net386 wbs_dat_o[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4318_ _1257_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5298_ _1943_ _1936_ _1944_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput397 net397 wbs_dat_o[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input37_I mc14500_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__S _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ dffram.data\[26\]\[7\] dffram.data\[27\]\[7\] _0778_ _1191_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmultiplexer_411 irq[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_126_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5070__A1 _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3620__A2 _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5125__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ _1647_ _2062_ _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3551_ _2908_ _2910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5464__I _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3482_ dffram.data\[34\]\[0\] _2864_ _2865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6270_ _0227_ clknet_leaf_119_wb_clk_i dffram.data\[48\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5221_ _1894_ _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5152_ _1808_ _1845_ _1848_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4103_ dffram.data\[8\]\[4\] dffram.data\[9\]\[4\] _0703_ _1048_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5083_ dffram.data\[39\]\[6\] _1796_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3712__I _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4034_ _0661_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _2399_ _2411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4936_ dffram.data\[28\]\[1\] _1703_ _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4867_ _1650_ _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _0755_ _0758_ _0760_ _0763_ _0765_ _0766_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_6606_ _0563_ clknet_leaf_31_wb_clk_i dffram.data\[33\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4798_ dffram.data\[63\]\[7\] _1605_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3366__A1 wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6537_ _0494_ clknet_leaf_137_wb_clk_i net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3749_ _0692_ _0693_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _0425_ clknet_leaf_42_wb_clk_i dffram.data\[62\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6399_ _0356_ clknet_leaf_54_wb_clk_i dffram.data\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ dffram.data\[0\]\[3\] _2022_ _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4866__A1 _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3622__I _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output310_I net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4229__S0 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5284__I _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_128_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5770_ _2255_ _2257_ _2259_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2982_ _2452_ _2360_ _2453_ _2454_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_84_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4721_ _1468_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _1504_ _1509_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput30 blinker_do[1] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ _2921_ _2943_ _2945_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput52 mc14500_do[26] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_126_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput41 mc14500_do[16] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput63 mc14500_do[8] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3899__A2 _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5194__I _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4583_ dffram.data\[5\]\[2\] _1445_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput74 mc14500_sram_in[2] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6322_ _0279_ clknet_leaf_99_wb_clk_i dffram.data\[46\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3534_ _2866_ _2896_ _2899_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput85 qcpu_do[14] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput96 qcpu_do[24] net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3465_ _2323_ _2849_ _2853_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6253_ _0210_ clknet_leaf_164_wb_clk_i dffram.data\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4848__A1 _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ dffram.data\[50\]\[3\] _1876_ _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5922__I _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6184_ _0141_ clknet_leaf_117_wb_clk_i dffram.data\[49\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3396_ net240 _2790_ _2805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5135_ _1814_ _1832_ _1837_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input139_I qcpu_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _1568_ _1489_ _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5273__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ dffram.data\[24\]\[3\] dffram.data\[25\]\[3\] _0824_ _0963_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5968_ _2397_ _2398_ _2396_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4919_ _1689_ _1690_ _1692_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_43_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5899_ _2337_ _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__B1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output260_I net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3511__A1 _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_max_cap404_I _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3578__A1 _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3250_ net281 _2672_ _2673_ _2686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3181_ _2556_ _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4058__A2 _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5822_ _2260_ _2291_ _2294_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5753_ dffram.data\[12\]\[3\] _2244_ _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3569__A1 _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4230__A2 _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _1544_ _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5684_ _2202_ _2197_ _2203_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_96_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3437__I _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4635_ _1490_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4566_ _1440_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6305_ _0262_ clknet_leaf_106_wb_clk_i dffram.data\[20\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3517_ _2870_ _2883_ _2888_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5652__I _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4497_ net189 _1385_ _1386_ net86 _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_input256_I wbs_we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3448_ dffram.data\[36\]\[4\] _2842_ _2843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4297__A2 _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6236_ _0193_ clknet_leaf_129_wb_clk_i dffram.data\[50\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3379_ net237 _2790_ _2791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6167_ _0124_ clknet_leaf_174_wb_clk_i dffram.data\[26\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5118_ dffram.data\[24\]\[6\] _1819_ _1826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6098_ _0055_ clknet_leaf_23_wb_clk_i dffram.data\[59\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5246__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _1741_ _1776_ _1778_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_178_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A1 _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput220 net473 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput253 net442 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput231 net463 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput242 net455 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3810__I _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4906__I _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5960__A2 _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3257__I _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _1326_ _1327_ _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_41_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4351_ net116 _1277_ _0652_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4289__S _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4282_ dffram.data\[60\]\[7\] dffram.data\[61\]\[7\] _1194_ _1224_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3302_ _2726_ _2727_ _2728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6021_ net240 _2437_ _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3233_ _2475_ _2672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5228__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3164_ _2601_ _2613_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4816__I _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3720__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3095_ _2474_ net212 _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _2264_ _2278_ _2283_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3997_ _0770_ _0943_ _0790_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__I _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5736_ dffram.data\[40\]\[4\] _2237_ _2238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5667_ _2148_ _2188_ _2191_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4618_ _1199_ _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input67_I mc14500_sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _2144_ _2145_ _2147_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4549_ _1426_ net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5382__I _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5467__A1 _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6219_ _0176_ clknet_leaf_118_wb_clk_i dffram.data\[52\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3831__S _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3805__I _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__I _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4636__I _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3920_ _0736_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5630__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__I2 _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ dffram.data\[38\]\[0\] dffram.data\[39\]\[0\] _0799_ _0800_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3782_ _0726_ _0727_ _0729_ _0730_ _0682_ _0690_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_6_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6570_ _0527_ clknet_leaf_148_wb_clk_i wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _2071_ _2092_ _2096_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _2017_ _2041_ _2046_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4403_ _0637_ net137 _1312_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__3715__I _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5383_ _1999_ _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4334_ _1262_ _1267_ net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3172__A2 wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4265_ dffram.data\[0\]\[7\] dffram.data\[1\]\[7\] _1192_ _1207_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6004_ net270 _2422_ _2425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5930__I _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4196_ dffram.data\[28\]\[6\] dffram.data\[29\]\[6\] _0795_ _1139_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3216_ net388 _2654_ _2647_ _2657_ _2658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3147_ _2597_ _2598_ _2599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input121_I qcpu_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input219_I wbs_adr_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ _2467_ _2525_ _2469_ _2539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5719_ dffram.data\[16\]\[6\] _2224_ _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4360__A1 _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4456__I _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3360__I _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__A1 _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__I _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold75_I wbs_dat_i[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4351__A1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4050_ _0970_ _0979_ _0988_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xinput6 ay8913_do[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5851__A1 _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3001_ _2467_ _2459_ _2468_ _2466_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4952_ _1486_ _1583_ _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ dffram.data\[4\]\[1\] dffram.data\[5\]\[1\] _0728_ _0851_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4883_ _1610_ _1666_ _1668_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3834_ dffram.data\[54\]\[0\] dffram.data\[55\]\[0\] _0782_ _0783_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6622_ _0579_ clknet_leaf_178_wb_clk_i dffram.data\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3765_ _0687_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6553_ _0510_ clknet_leaf_151_wb_clk_i wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5504_ _1472_ _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_95_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3696_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6484_ _0441_ clknet_leaf_130_wb_clk_i net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5435_ dffram.data\[46\]\[0\] _2036_ _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput310 net310 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput343 net343 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput332 net332 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4342__A1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput321 net321 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput354 net354 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput365 net365 rst_hellorld vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5366_ dffram.data\[47\]\[2\] _1987_ _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input169_I sid_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput376 net376 wbs_dat_o[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput387 net387 wbs_dat_o[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4317_ _1248_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5297_ dffram.data\[48\]\[3\] _1937_ _1944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput398 net398 wbs_dat_o[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ dffram.data\[24\]\[7\] dffram.data\[25\]\[7\] _1189_ _1190_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmultiplexer_412 irq[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_126_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5842__A1 dffram.data\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4179_ dffram.data\[32\]\[5\] dffram.data\[33\]\[5\] _0754_ _1123_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_104_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output290_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3767__S0 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5833__A1 dffram.data\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Left_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3550_ _2908_ _2909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3481_ _2862_ _2864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5220_ _1431_ _1700_ _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_90_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5151_ dffram.data\[51\]\[1\] _1846_ _1848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4102_ _0792_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5082_ _1756_ _1795_ _1798_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5824__A1 _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _0908_ _0978_ _0723_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_108_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _2409_ _2410_ _2408_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _1678_ _1702_ _1704_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3063__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6001__A1 net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4866_ _1619_ _1651_ _1656_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4797_ _1562_ _1604_ _1608_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3817_ _0745_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6605_ _0562_ clknet_leaf_30_wb_clk_i dffram.data\[33\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3748_ _0691_ _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _0493_ clknet_leaf_136_wb_clk_i net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _0424_ clknet_leaf_61_wb_clk_i dffram.data\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3679_ _0633_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6398_ _0355_ clknet_leaf_53_wb_clk_i dffram.data\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ _2005_ _2021_ _2025_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5349_ dffram.data\[21\]\[4\] _1978_ _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4000__S _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5815__A1 _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4734__I _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output303_I net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4229__S1 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__I _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__I _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3293__A1 wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3045__A1 net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2981_ _2441_ _2454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4793__A1 _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ _1554_ _1555_ _1557_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _1508_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_168_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_168_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput20 ay8913_do[27] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput31 blinker_do[2] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5475__I _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3602_ dffram.data\[19\]\[0\] _2944_ _2945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput53 mc14500_do[27] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput42 mc14500_do[17] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput64 mc14500_do[9] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4582_ _1454_ _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput75 mc14500_sram_in[3] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ _0278_ clknet_leaf_99_wb_clk_i dffram.data\[46\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3533_ dffram.data\[32\]\[1\] _2897_ _2899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput86 qcpu_do[15] net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput97 qcpu_do[25] net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3464_ dffram.data\[35\]\[2\] _2850_ _2853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6252_ _0209_ clknet_leaf_164_wb_clk_i dffram.data\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5203_ _1813_ _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6183_ _0140_ clknet_leaf_161_wb_clk_i dffram.data\[49\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3395_ wb_counter\[25\] _2803_ _2804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5134_ dffram.data\[52\]\[3\] _1833_ _1837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5065_ _1760_ _1782_ _1787_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4016_ _0962_ net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3284__A1 wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input201_I sn76489_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ net225 _2391_ _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4918_ dffram.data\[54\]\[4\] _1691_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _2337_ _2344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input97_I qcpu_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4536__A1 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ dffram.data\[57\]\[6\] _1642_ _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4536__B2 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_73_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_168_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _0476_ clknet_leaf_150_wb_clk_i net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_31_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4729__I _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__I0 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold8_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_82_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3275__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4527__A1 _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3180_ _2581_ _2627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5821_ dffram.data\[13\]\[1\] _2292_ _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5752_ _2202_ _2243_ _2247_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4766__A1 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ net403 _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5683_ dffram.data\[11\]\[2\] _2198_ _2203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4518__A1 _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _1460_ _1491_ _1496_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_116_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4565_ _1431_ _1439_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ _0261_ clknet_leaf_106_wb_clk_i dffram.data\[20\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3516_ dffram.data\[33\]\[3\] _2884_ _2888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4496_ _1387_ _1389_ net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_139_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3447_ _2834_ _2842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6235_ _0192_ clknet_leaf_113_wb_clk_i dffram.data\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input151_I qcpu_sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3378_ _2692_ _2790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6166_ _0123_ clknet_leaf_175_wb_clk_i dffram.data\[26\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ _0054_ clknet_leaf_23_wb_clk_i dffram.data\[59\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5117_ _1824_ _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ dffram.data\[25\]\[0\] _1777_ _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input12_I ay8913_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__B1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4057__I0 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3009__A1 _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4509__B2 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__A1 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output370_I net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput210 sn76489_do[9] net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput243 net462 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput254 net466 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput232 net458 net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput221 net471 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_98_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4296__I0 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__A2 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3420__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4350_ _0623_ _0636_ _1278_ _1252_ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_50_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3301_ _2723_ _2724_ _2719_ _2727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_39_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4281_ dffram.data\[58\]\[7\] dffram.data\[59\]\[7\] _0778_ _1223_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_111_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6020_ _2359_ _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3232_ _2663_ _2670_ _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input4_I ay8913_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ net379 _2609_ _2602_ _2612_ _2613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_87_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3094_ _2520_ _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5804_ dffram.data\[15\]\[3\] _2279_ _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4739__A1 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_112_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _0939_ _0940_ _0941_ _0942_ _0881_ _0883_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_45_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _2229_ _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_118_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ dffram.data\[41\]\[5\] _2189_ _2191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input199_I sn76489_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5164__A1 _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4617_ _1482_ net469 _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_131_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5663__I _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ dffram.data\[43\]\[4\] _2146_ _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4548_ net103 _1411_ _1407_ net57 _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__A1 _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4479_ _1324_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_111_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _0175_ clknet_leaf_119_wb_clk_i dffram.data\[52\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3868__I3 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _0106_ clknet_leaf_174_wb_clk_i dffram.data\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4427__B1 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4978__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__I _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_69_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A1 _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3850_ _0753_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5394__A1 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3268__I _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3781_ dffram.data\[6\]\[0\] dffram.data\[7\]\[0\] _0671_ _0730_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5520_ dffram.data\[10\]\[2\] _2093_ _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3944__A2 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5483__I _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5451_ dffram.data\[46\]\[7\] _2042_ _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _1311_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5382_ _1999_ _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_10_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ net143 _1263_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4264_ _1199_ _1205_ _0722_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6003_ _2423_ _2424_ _2419_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3215_ _2655_ _2656_ _2657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4195_ dffram.data\[26\]\[6\] dffram.data\[27\]\[6\] _0964_ _1138_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3146_ net263 _2582_ _2583_ _2598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3077_ _2534_ _2535_ _2536_ _2537_ _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_input114_I qcpu_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__A1 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ _2210_ _2223_ _2226_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3979_ _0739_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ dffram.data\[17\]\[7\] _2176_ _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3906__I _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output333_I net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4737__I _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5568__I _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3926__A2 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold68_I wbs_dat_i[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3816__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4351__A2 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__I _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3551__I _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 ay8913_do[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3000_ net251 _2462_ _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_99_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5478__I _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4951_ _1697_ _1708_ _1713_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3902_ dffram.data\[2\]\[1\] dffram.data\[3\]\[1\] _0849_ _0850_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ dffram.data\[55\]\[0\] _1667_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3833_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6621_ _0578_ clknet_leaf_10_wb_clk_i dffram.data\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3764_ _0681_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6552_ _0509_ clknet_leaf_151_wb_clk_i wb_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_27_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5503_ _2082_ _2078_ _2083_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3695_ design_select\[2\] _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_70_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5119__A1 _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A2 _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _0440_ clknet_leaf_130_wb_clk_i net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5434_ _2034_ _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_95_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput300 net300 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput344 net344 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput333 net333 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput322 net322 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput311 net311 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput355 net355 qcpu_sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _1939_ _1986_ _1989_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput366 net366 rst_mc14500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput377 net377 wbs_dat_o[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4316_ _1251_ _1256_ net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5296_ _1813_ _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput399 net399 wbs_dat_o[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput388 net388 wbs_dat_o[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4247_ _0777_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xmultiplexer_413 irq[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_126_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4178_ _1005_ _1121_ _1067_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3129_ net260 _2582_ _2583_ _2584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3605__A1 _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3908__A2 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output283_I net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3767__S1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3687__A4 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A2 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3480_ _2862_ _2863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_77_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A1 _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_102_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_90_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5150_ _1802_ _1845_ _1847_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ _1042_ _1043_ _1044_ _1045_ _0854_ _0986_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5081_ dffram.data\[39\]\[5\] _1796_ _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4032_ _0971_ _0973_ _0974_ _0975_ _0976_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_108_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5983_ net229 _2404_ _2410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ dffram.data\[28\]\[0\] _1703_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_111_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5001__I _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ dffram.data\[56\]\[3\] _1652_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4796_ dffram.data\[63\]\[6\] _1605_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3816_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6604_ _0561_ clknet_leaf_28_wb_clk_i dffram.data\[34\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5760__A1 _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3747_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3456__I _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6535_ _0492_ clknet_leaf_137_wb_clk_i net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input181_I sid_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__B1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_158_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ _0423_ clknet_leaf_47_wb_clk_i dffram.data\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3678_ design_select\[0\] _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_3_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6397_ _0354_ clknet_leaf_53_wb_clk_i dffram.data\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_120_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ dffram.data\[0\]\[2\] _2022_ _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input42_I mc14500_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _1970_ _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5279_ _1888_ _1928_ _1931_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__A1 _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5581__I _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _1506_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_72_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 ay8913_do[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput21 ay8913_do[2] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3601_ _2942_ _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput32 hellorld_do net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput54 mc14500_do[28] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput43 mc14500_do[18] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6320_ _0277_ clknet_leaf_99_wb_clk_i dffram.data\[46\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4581_ _1453_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput76 mc14500_sram_in[4] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput65 mc14500_sram_addr[0] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3532_ _2861_ _2896_ _2898_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 qcpu_do[16] net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput98 qcpu_do[26] net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_137_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3463_ _2321_ _2849_ _2852_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6251_ _0208_ clknet_leaf_68_wb_clk_i dffram.data\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5202_ _1880_ _1875_ _1881_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6182_ _0139_ clknet_leaf_161_wb_clk_i dffram.data\[49\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3394_ _2802_ _2795_ _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5133_ _1811_ _1832_ _1836_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3940__S _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5064_ dffram.data\[25\]\[7\] _1783_ _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4015_ _0932_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4481__A1 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__B2 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ net259 _2386_ _2397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5897_ _2325_ _2338_ _2343_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4917_ _1679_ _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_43_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ _1625_ _1641_ _1644_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5733__A1 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4779_ _1504_ _1489_ _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3744__B1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6518_ _0475_ clknet_leaf_158_wb_clk_i net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _0406_ clknet_leaf_56_wb_clk_i dffram.data\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__S _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3898__I1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__I _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold50_I wbs_cyc_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ _2255_ _2291_ _2293_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_85_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5751_ dffram.data\[12\]\[2\] _2244_ _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5486__I _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _1539_ _1541_ _1543_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5682_ _2070_ _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4633_ dffram.data\[31\]\[3\] _1492_ _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4564_ _1438_ _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_124_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6303_ _0260_ clknet_leaf_103_wb_clk_i dffram.data\[20\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3515_ _2868_ _2883_ _2887_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4495_ net166 _1383_ _1388_ net39 net6 _1379_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_6234_ _0191_ clknet_leaf_108_wb_clk_i dffram.data\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3446_ _2834_ _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3377_ _2786_ _2788_ _2789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6165_ _0122_ clknet_leaf_174_wb_clk_i dffram.data\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input144_I qcpu_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6096_ _0053_ clknet_leaf_26_wb_clk_i dffram.data\[59\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5116_ _1472_ _1824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _1775_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4454__A1 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__B2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3009__A2 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5949_ net286 _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5954__A1 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__I _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output363_I net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3193__A1 net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6020__I _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4693__A1 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput200 sn76489_do[25] net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput211 wb_rst_i net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput233 net449 net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput244 net460 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput222 net468 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput255 wbs_stb_i net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4996__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3755__S _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3300_ _2481_ net256 _2549_ _2726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4280_ dffram.data\[56\]\[7\] dffram.data\[57\]\[7\] _1189_ _1222_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_111_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3231_ wb_counter\[28\] _2670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3162_ _2610_ _2611_ _2612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3093_ _2534_ wb_counter\[8\] _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _2262_ _2278_ _2282_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3995_ dffram.data\[54\]\[2\] dffram.data\[55\]\[2\] _0782_ _0942_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _2229_ _2236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_118_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5665_ _2144_ _2188_ _2190_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_152_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_152_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5944__I _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4616_ net255 net222 _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5596_ _2134_ _2146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4547_ _1425_ net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _1373_ _1374_ net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6217_ _0174_ clknet_leaf_118_wb_clk_i dffram.data\[52\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3429_ net426 _2829_ _1481_ _2830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _0105_ clknet_leaf_173_wb_clk_i dffram.data\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4427__A1 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4427__B2 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6079_ _0036_ clknet_leaf_18_wb_clk_i dffram.data\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2989__A1 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__I _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4210__S0 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__A1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__I _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__A2 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4277__S0 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ dffram.data\[4\]\[0\] dffram.data\[5\]\[0\] _0728_ _0729_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _2015_ _2041_ _2045_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_113_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4401_ _0717_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_97_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5146__A2 _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5381_ _1858_ _1700_ _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4332_ _1262_ _1266_ net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4263_ _1201_ _1202_ _1203_ _1204_ _0680_ _0688_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6002_ net235 _2415_ _2424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3214_ net274 _2649_ _2650_ _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4194_ dffram.data\[24\]\[6\] dffram.data\[25\]\[6\] _0671_ _1137_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3145_ _2596_ wb_counter\[15\] _2597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5004__I _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3076_ _2472_ wb_counter\[6\] _2488_ _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5082__A1 _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__I _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input107_I qcpu_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3459__I _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ dffram.data\[12\]\[2\] dffram.data\[13\]\[2\] _0740_ _0925_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ dffram.data\[16\]\[5\] _2224_ _2226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3396__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input72_I mc14500_sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _2150_ _2175_ _2179_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _1983_ _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A1 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output326_I net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3320__A1 _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3871__A2 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5073__A1 dffram.data\[39\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput8 ay8913_do[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ dffram.data\[28\]\[7\] _1709_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4811__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3901_ _0828_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4881_ _1665_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3832_ _0707_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6620_ _0577_ clknet_leaf_2_wb_clk_i dffram.data\[32\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6551_ _0508_ clknet_leaf_155_wb_clk_i wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5502_ dffram.data\[45\]\[5\] _2079_ _2083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5494__I _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3763_ dffram.data\[22\]\[0\] dffram.data\[23\]\[0\] _0711_ _0712_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_148_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4104__S _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3694_ _0631_ _0645_ net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_95_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6482_ _0439_ clknet_leaf_129_wb_clk_i net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5433_ _2034_ _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput301 net301 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput334 net334 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput323 net323 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5364_ dffram.data\[47\]\[1\] _1987_ _1989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3925__I0 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput312 net312 io_oeb[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput345 net345 io_out[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput356 net356 qcpu_sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput367 net367 rst_qcpu vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4315_ _1255_ _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput378 net378 wbs_dat_o[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5295_ _1941_ _1936_ _1942_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput389 net389 wbs_dat_o[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4246_ _0694_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4177_ _1117_ _1118_ _1119_ _1120_ _0835_ _1088_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xmultiplexer_414 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_3128_ _2556_ _2583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3059_ wb_counter\[4\] _2522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3917__I _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output276_I net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__I _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4483__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold80_I wbs_dat_i[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3907__I0 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3532__A1 _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5080_ _1752_ _1795_ _1797_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4100_ dffram.data\[6\]\[4\] dffram.data\[7\]\[4\] _0852_ _1045_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4031_ _0714_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ net263 _2400_ _2409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3599__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4933_ _1701_ _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _1617_ _1651_ _1655_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_59_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4795_ _1559_ _1604_ _1607_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3815_ _0680_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6603_ _0560_ clknet_leaf_28_wb_clk_i dffram.data\[34\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3746_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6534_ _0491_ clknet_leaf_137_wb_clk_i net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6465_ _0422_ clknet_leaf_47_wb_clk_i dffram.data\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3771__B2 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3771__A1 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3677_ _0620_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5416_ _2003_ _2021_ _2024_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input174_I sid_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ _0353_ clknet_leaf_52_wb_clk_i dffram.data\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__I net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5347_ _1970_ _1977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3523__A1 _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ dffram.data\[22\]\[5\] _1929_ _1931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input35_I mc14500_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4229_ _1168_ _1169_ _1170_ _1171_ _0835_ _1088_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4484__C1 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__A1 _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4009__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__B1 _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output393_I net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5102__I _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4242__A2 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput11 ay8913_do[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput22 ay8913_do[3] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3600_ _2942_ _2943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4580_ net245 _1451_ _0642_ net155 _1452_ net74 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
Xinput33 io_in[0] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput55 mc14500_do[29] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput44 mc14500_do[19] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3531_ dffram.data\[32\]\[0\] _2897_ _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput77 mc14500_sram_in[5] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput66 mc14500_sram_addr[1] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput88 qcpu_do[17] net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3462_ dffram.data\[35\]\[1\] _2850_ _2852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6250_ _0207_ clknet_leaf_68_wb_clk_i dffram.data\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput99 qcpu_do[27] net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ dffram.data\[50\]\[2\] _1876_ _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6181_ _0138_ clknet_leaf_164_wb_clk_i dffram.data\[49\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3393_ wb_counter\[24\] _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5132_ dffram.data\[52\]\[2\] _1833_ _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_177_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_177_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_106_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5258__A1 _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _1758_ _1782_ _1786_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4337__B net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ _0938_ _0944_ _0952_ _0960_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_90_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5430__A1 _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5965_ _2393_ _2394_ _2396_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5896_ dffram.data\[62\]\[3\] _2339_ _2343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_101_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ _1679_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4847_ dffram.data\[57\]\[5\] _1642_ _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _1565_ _1591_ _1596_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__A1 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5682__I _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3729_ net147 _0677_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3744__B2 net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6517_ _0474_ clknet_leaf_150_wb_clk_i net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_140_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _0405_ clknet_leaf_57_wb_clk_i dffram.data\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _0336_ clknet_leaf_100_wb_clk_i dffram.data\[42\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_54_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4457__C1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3930__I _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A2 _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3735__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4202__S _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__C1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5767__I _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5750_ _2200_ _2243_ _2246_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5681_ _2200_ _2197_ _2201_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ dffram.data\[2\]\[0\] _1542_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _1455_ _1491_ _1495_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4563_ _1433_ _1437_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4494_ _1324_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6302_ _0259_ clknet_leaf_103_wb_clk_i dffram.data\[20\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3514_ dffram.data\[33\]\[2\] _2884_ _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3445_ _2325_ _2835_ _2840_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6233_ _0190_ clknet_leaf_108_wb_clk_i dffram.data\[23\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5007__I _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3376_ _2787_ _2782_ _2788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6164_ _0121_ clknet_leaf_175_wb_clk_i dffram.data\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6095_ _0052_ clknet_leaf_33_wb_clk_i dffram.data\[59\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5115_ _1822_ _1818_ _1823_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input137_I qcpu_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1775_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5651__A1 _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_74_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4057__I2 _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__I _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5948_ _2382_ _2383_ _2381_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5879_ dffram.data\[14\]\[5\] _2329_ _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3197__I _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3861__S _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput201 sn76489_do[26] net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6530__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput245 net430 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput234 net425 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput212 net467 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput223 net419 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput256 wbs_we_i net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_98_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4491__I _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3835__I _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3230_ _2549_ _2669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3570__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ net265 _2604_ _2605_ _2611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_87_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3092_ _2550_ _2551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5497__I _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5802_ dffram.data\[15\]\[2\] _2279_ _2282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3994_ dffram.data\[52\]\[2\] dffram.data\[53\]\[2\] _0878_ _0941_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5733_ _2204_ _2230_ _2235_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3946__S _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ dffram.data\[41\]\[4\] _2189_ _2190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5595_ _2134_ _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4615_ _1481_ _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4546_ net101 _1411_ _1407_ net55 _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_131_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_121_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4477_ net185 _1333_ _1350_ net3 _1339_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__3970__I1 dffram.data\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6216_ _0173_ clknet_leaf_119_wb_clk_i dffram.data\[52\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _2525_ _2350_ _2456_ _2829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5872__A1 _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3480__I _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _0104_ clknet_leaf_16_wb_clk_i dffram.data\[54\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4675__A2 _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3359_ _2752_ _2772_ _2774_ _2764_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5624__A1 _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _0035_ clknet_leaf_67_wb_clk_i dffram.data\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5029_ dffram.data\[49\]\[1\] _1764_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4017__S _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5870__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5863__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4486__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_82_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4277__S1 _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4400_ _1302_ _1310_ net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5380_ _1801_ _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_10_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ net142 _1263_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4262_ dffram.data\[22\]\[7\] dffram.data\[23\]\[7\] _0660_ _1204_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 dffram.data\[38\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ net269 _2422_ _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3213_ _2641_ wb_counter\[25\] _2655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4193_ _1136_ net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3144_ _2571_ _2596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3075_ net285 _2520_ _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_177_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__A1 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3977_ dffram.data\[10\]\[2\] dffram.data\[11\]\[2\] _0923_ _0924_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5716_ _2206_ _2223_ _2225_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ dffram.data\[17\]\[6\] _2176_ _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input65_I mc14500_sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5578_ _2060_ _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4529_ _1324_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4300__S _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5845__A1 _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output319_I net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6026__I _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A1 _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 ay8913_do[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3075__A1 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ dffram.data\[0\]\[1\] dffram.data\[1\]\[1\] _0662_ _0848_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6013__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4880_ _1665_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3831_ dffram.data\[52\]\[0\] dffram.data\[53\]\[0\] _0779_ _0780_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3762_ _0708_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6550_ _0507_ clknet_leaf_155_wb_clk_i wb_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ _2081_ _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3693_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_70_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _0438_ clknet_leaf_132_wb_clk_i net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_27_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5432_ _1984_ _2033_ _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput335 net335 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput324 net324 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5363_ _1934_ _1986_ _1988_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput313 net313 io_oeb[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput302 net302 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput346 net346 io_out[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput357 net357 qcpu_sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4314_ _0638_ _0645_ _0651_ _1254_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4120__S _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput368 net368 rst_sid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5294_ dffram.data\[48\]\[2\] _1937_ _1942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput379 net379 wbs_dat_o[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4245_ _1187_ net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_143_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4176_ dffram.data\[54\]\[5\] dffram.data\[55\]\[5\] _0779_ _1120_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmultiplexer_415 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_3127_ _2581_ _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input217_I wbs_adr_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3066__A1 _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ net283 _2520_ _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6004__A1 net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5685__I _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3369__A2 wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output269_I net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3933__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4177__S0 _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__I _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4557__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold73_I wbs_dat_i[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_77_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3907__I1 _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A1 _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4030_ _0784_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5285__A2 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_108_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3048__A1 _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _2406_ _2407_ _2408_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3599__A2 _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4932_ _1701_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__A1 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6602_ _0559_ clknet_leaf_29_wb_clk_i dffram.data\[34\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4863_ dffram.data\[56\]\[2\] _1652_ _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4548__B2 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4794_ dffram.data\[63\]\[5\] _1605_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3814_ dffram.data\[62\]\[0\] dffram.data\[63\]\[0\] _0762_ _0763_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3745_ _0692_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _0490_ clknet_leaf_139_wb_clk_i net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3954__S _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _0421_ clknet_leaf_47_wb_clk_i dffram.data\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3771__A2 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3676_ _0627_ _0631_ net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5415_ dffram.data\[0\]\[1\] _2022_ _2024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3753__I _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _0352_ clknet_leaf_98_wb_clk_i dffram.data\[41\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4720__A1 _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _1943_ _1971_ _1976_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input167_I sid_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5277_ _1884_ _1928_ _1930_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4228_ dffram.data\[54\]\[6\] dffram.data\[55\]\[6\] _0779_ _1171_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_34_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input28_I ay8913_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4159_ _0792_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3039__A1 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3421__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__A1 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_43_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4539__B2 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__A1 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__S _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__I _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__I _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4778__A1 _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3838__I _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput12 ay8913_do[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput23 ay8913_do[4] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput45 mc14500_do[1] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput34 mc14500_do[0] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3530_ _2895_ _2897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput78 mc14500_sram_in[6] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput67 mc14500_sram_addr[2] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 mc14500_do[2] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput89 qcpu_do[18] net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3461_ _2316_ _2849_ _2851_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4702__A1 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ _1810_ _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6180_ _0137_ clknet_leaf_165_wb_clk_i dffram.data\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3392_ _2792_ _2800_ _2801_ _2785_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5131_ _1808_ _1832_ _1835_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5062_ dffram.data\[25\]\[6\] _1783_ _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4013_ _0806_ _0959_ _0819_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_146_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_146_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5964_ _2395_ _2396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5895_ _2323_ _2338_ _2342_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3441__A1 _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4915_ _1553_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _1621_ _1641_ _1643_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ dffram.data\[59\]\[7\] _1592_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3744__A2 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__I _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _0473_ clknet_leaf_149_wb_clk_i net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4941__A1 _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3728_ _0646_ design_select\[1\] design_select\[0\] _0624_ _0677_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_71_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _0404_ clknet_leaf_59_wb_clk_i dffram.data\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _2938_ _2975_ _2979_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _0335_ clknet_leaf_100_wb_clk_i dffram.data\[42\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5329_ _1945_ _1964_ _1966_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3898__I3 _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output301_I net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5873__I _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4448__B1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__I _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5680_ dffram.data\[11\]\[1\] _2198_ _2201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4700_ _1540_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5176__A1 _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ dffram.data\[31\]\[2\] _1492_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4223__I0 _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4562_ _0666_ _1436_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6301_ _0258_ clknet_leaf_103_wb_clk_i dffram.data\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3513_ _2866_ _2883_ _2886_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4493_ net188 _1385_ _1386_ net85 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3444_ dffram.data\[36\]\[3\] _2836_ _2840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6232_ _0189_ clknet_leaf_113_wb_clk_i dffram.data\[23\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6163_ _0120_ clknet_leaf_172_wb_clk_i dffram.data\[27\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3375_ wb_counter\[21\] _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6094_ _0051_ clknet_leaf_29_wb_clk_i dffram.data\[59\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5114_ dffram.data\[24\]\[5\] _1819_ _1823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5045_ _1727_ _1633_ _1775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5651__A2 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3478__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5947_ net251 _2377_ _2383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5878_ _1469_ _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input95_I qcpu_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__I _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_117_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_43_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4829_ _1432_ _1505_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4914__A1 _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4390__A2 _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output349_I net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput202 sn76489_do[27] net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_126_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput224 net453 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput235 net461 net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput213 net438 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput246 net448 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_135_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_128_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3708__A2 design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4381__A2 _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _2596_ wb_counter\[17\] _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xhold1 net514 net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3091_ _2549_ _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_167_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5801_ _2260_ _2278_ _2281_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5732_ dffram.data\[40\]\[3\] _2231_ _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3993_ dffram.data\[50\]\[2\] dffram.data\[51\]\[2\] _0775_ _0940_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5663_ _2181_ _2189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5594_ _2076_ _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _1480_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4545_ _1424_ net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_131_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4372__A2 _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3962__S _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4476_ net163 _1316_ _1317_ net82 net36 _1352_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_41_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__A1 _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4857__I _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6215_ _0172_ clknet_leaf_161_wb_clk_i dffram.data\[52\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3427_ _2487_ _2459_ _2828_ _2541_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6146_ _0103_ clknet_leaf_169_wb_clk_i dffram.data\[54\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3358_ net232 _2773_ _2774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_161_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_161_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6077_ _0034_ clknet_leaf_18_wb_clk_i dffram.data\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3289_ net251 _2705_ _2717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input10_I ay8913_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _1741_ _1763_ _1765_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output299_I net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5312__A1 _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3626__A1 _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4208__S _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A1 _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4007__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__A1 _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _1262_ _1265_ net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_50_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4261_ dffram.data\[20\]\[7\] dffram.data\[21\]\[7\] _0660_ _1203_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5303__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__I _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6000_ _2399_ _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3212_ _2490_ _2654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input2_I ay8913_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _1110_ _1135_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_59_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3143_ _2578_ _2595_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3617__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3074_ _1161_ _1186_ _2476_ _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5301__I _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__S _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3976_ _0736_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5715_ dffram.data\[16\]\[4\] _2224_ _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3756__I _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5790__A1 _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5646_ _2148_ _2175_ _2178_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input197_I sn76489_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _2088_ _2126_ _2131_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4528_ net198 _1402_ _1403_ net95 _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4459_ net206 _1322_ _1361_ net24 _1339_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_input58_I mc14500_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4587__I _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__C1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6129_ _0086_ clknet_leaf_5_wb_clk_i dffram.data\[56\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5211__I _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3084__A2 wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3666__I design_select\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__A1 _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__I _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3075__A2 _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3777__S _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3830_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3761_ dffram.data\[20\]\[0\] dffram.data\[21\]\[0\] _0709_ _0710_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5500_ _1468_ _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3576__I _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3692_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6480_ _0437_ clknet_leaf_133_wb_clk_i net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5791__I _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _1523_ _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput325 net325 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5362_ dffram.data\[47\]\[0\] _1987_ _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3925__I2 _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput314 net314 io_oeb[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput303 net303 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput369 net369 rst_sn76489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput347 net347 io_out[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput336 net336 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput358 net358 qcpu_sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4313_ _0632_ net182 _1253_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _1810_ _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_61_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _1161_ _1186_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_143_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4175_ dffram.data\[52\]\[5\] dffram.data\[53\]\[5\] _0828_ _1119_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmultiplexer_416 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_3126_ _2475_ _2581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I qcpu_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3057_ _2474_ _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A1 _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3369__A3 wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0901_ _0902_ _0903_ _0905_ _0836_ _0837_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_73_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _1632_ _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__S1 _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output331_I net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4780__I _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A1 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_hold66_I wbs_dat_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4221__S _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5116__I _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_108_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4493__B2 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _2395_ _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_121_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4931_ _1486_ _1700_ _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5993__A1 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _1615_ _1651_ _1654_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_103_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3813_ _0761_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _0558_ clknet_leaf_30_wb_clk_i dffram.data\[34\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4793_ _1554_ _1604_ _1606_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3744_ net219 _0675_ _0685_ net149 _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6532_ _0489_ clknet_leaf_137_wb_clk_i net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _0420_ clknet_leaf_39_wb_clk_i dffram.data\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3675_ _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4131__S _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5414_ _1998_ _2021_ _2023_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6394_ _0351_ clknet_leaf_98_wb_clk_i dffram.data\[41\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__I1 dffram.data\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5345_ dffram.data\[21\]\[3\] _1972_ _1976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3970__S _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5276_ dffram.data\[22\]\[4\] _1929_ _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_68_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4227_ dffram.data\[52\]\[6\] dffram.data\[53\]\[6\] _0828_ _1170_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4484__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4484__A1 net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3287__A2 wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4158_ _1098_ _1099_ _1100_ _1101_ _0836_ _0986_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4089_ _0823_ _1033_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3109_ _2547_ _2566_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output281_I net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__A1 _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5727__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput13 ay8913_do[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 ay8913_do[5] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 mc14500_do[20] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput35 mc14500_do[10] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_107_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput68 mc14500_sram_addr[3] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput79 mc14500_sram_in[7] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput57 mc14500_do[30] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ dffram.data\[35\]\[0\] _2850_ _2851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ net239 _2790_ _2801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ dffram.data\[52\]\[1\] _1833_ _1835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _1756_ _1782_ _1785_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4012_ _0953_ _0955_ _0956_ _0958_ _0815_ _0816_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__4466__A1 _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5963_ _2362_ _2395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5966__A1 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4914_ _1687_ _1680_ _1688_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5894_ dffram.data\[62\]\[2\] _2339_ _2342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5718__A1 _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4845_ dffram.data\[57\]\[4\] _1642_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_115_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4776_ _1562_ _1591_ _1595_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3727_ net217 _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6515_ _0472_ clknet_leaf_149_wb_clk_i net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_125_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3764__I _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6446_ _0403_ clknet_leaf_52_wb_clk_i dffram.data\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3658_ dffram.data\[9\]\[6\] _2976_ _2979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3589_ _2932_ _2933_ _2935_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6377_ _0334_ clknet_leaf_101_wb_clk_i dffram.data\[42\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ dffram.data\[8\]\[4\] _1965_ _1966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input40_I mc14500_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4595__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4457__B2 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A1 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ dffram.data\[7\]\[6\] _1916_ _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3004__I net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4232__I1 dffram.data\[35\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4448__A1 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4448__B2 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_157_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _1449_ _1491_ _1494_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _0257_ clknet_leaf_103_wb_clk_i dffram.data\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3726__A3 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ net211 _1434_ _1435_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_13_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3512_ dffram.data\[33\]\[1\] _2884_ _2886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4492_ _1341_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3443_ _2323_ _2835_ _2839_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6231_ _0188_ clknet_leaf_107_wb_clk_i dffram.data\[23\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _0119_ clknet_leaf_172_wb_clk_i dffram.data\[27\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5113_ _1821_ _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3374_ wb_counter\[22\] _2786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6093_ _0050_ clknet_leaf_33_wb_clk_i dffram.data\[59\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5304__I _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5044_ _1760_ _1769_ _1774_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3111__A1 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4611__A1 dffram.data\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ net285 _2372_ _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5877_ _2327_ _2328_ _2330_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _1629_ _1622_ _1630_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4214__I1 dffram.data\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input88_I qcpu_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4759_ _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3494__I _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3427__C _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_83_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6429_ _0386_ clknet_leaf_66_wb_clk_i dffram.data\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_12_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_8_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput236 net451 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput225 net452 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput203 sn76489_do[2] net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput214 net441 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput247 net450 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4850__A1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3669__I _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5884__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3708__A3 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3341__A1 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3353__B _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold2 net223 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3090_ _2548_ _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__I _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3579__I _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5800_ dffram.data\[15\]\[1\] _2279_ _2281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3992_ dffram.data\[48\]\[2\] dffram.data\[49\]\[2\] _0875_ _0939_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5731_ _2202_ _2230_ _2234_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5662_ _2181_ _2188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5593_ _2142_ _2135_ _2143_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4613_ net211 _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4544_ net100 _1411_ _1407_ net54 _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_64_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4475_ _1336_ _1371_ _1372_ net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _0171_ clknet_leaf_157_wb_clk_i dffram.data\[52\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3426_ net420 _2462_ _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6145_ _0102_ clknet_leaf_16_wb_clk_i dffram.data\[54\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _2704_ _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input142_I qcpu_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _0033_ clknet_leaf_18_wb_clk_i dffram.data\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5027_ dffram.data\[49\]\[0\] _1764_ _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3288_ wb_counter\[6\] _2715_ _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_130_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3399__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5929_ net245 _2368_ _2369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__A1 _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5076__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold96_I wbs_dat_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A1 _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3562__A1 dffram.data\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3862__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ dffram.data\[18\]\[7\] dffram.data\[19\]\[7\] _1200_ _1202_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _1116_ _1122_ _1128_ _1134_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3211_ _2646_ _2653_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3142_ net376 _2587_ _2579_ _2594_ _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_128_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3073_ _2472_ _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4814__A1 _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3975_ dffram.data\[8\]\[2\] dffram.data\[9\]\[2\] _0734_ _0922_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5714_ _2216_ _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5645_ dffram.data\[17\]\[5\] _2176_ _2178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5576_ dffram.data\[44\]\[7\] _2127_ _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3553__A1 _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _1410_ _1412_ net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3943__I3 _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4868__I _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4458_ _1349_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3305__A1 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3409_ _2792_ _2813_ _2815_ _2806_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4389_ net130 _1304_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_102_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6128_ _0085_ clknet_leaf_5_wb_clk_i dffram.data\[56\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5699__I _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _0016_ clknet_leaf_15_wb_clk_i dffram.data\[31\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4805__A1 _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4108__I _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3012__I _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__A2 _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__A1 _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4044__S _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3544__A1 _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3682__I design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5049__A1 _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4219__S _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4018__I _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4024__A2 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3760_ _0708_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3691_ _0622_ _0618_ design_select\[0\] _0639_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5430_ _2017_ _2027_ _2032_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout405_I net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput326 net326 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5361_ _1985_ _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput315 net315 io_oeb[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput304 net304 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput337 net337 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput348 net348 io_out[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput359 net359 qcpu_sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _0623_ _0621_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_61_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _1939_ _1936_ _1940_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4243_ _1167_ _1173_ _1179_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_143_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_406 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_93_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4174_ dffram.data\[50\]\[5\] dffram.data\[51\]\[5\] _1007_ _1118_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xmultiplexer_417 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_3125_ _2572_ wb_counter\[12\] _2580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3056_ _1055_ _1082_ _2503_ _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_89_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3968__S _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input105_I qcpu_do[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3958_ dffram.data\[30\]\[2\] dffram.data\[31\]\[2\] _0904_ _0905_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3889_ _0689_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input70_I mc14500_sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5628_ _2152_ _2161_ _2166_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _2119_ _2121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__A1 _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__I net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output324_I net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4039__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__C1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__A1 _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold59_I wbs_adr_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5442__A1 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _1699_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ dffram.data\[56\]\[1\] _1652_ _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3812_ _0701_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6600_ _0557_ clknet_leaf_32_wb_clk_i dffram.data\[34\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4792_ dffram.data\[63\]\[4\] _1605_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3743_ net68 _0683_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6531_ _0488_ clknet_leaf_137_wb_clk_i net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6462_ _0419_ clknet_leaf_46_wb_clk_i dffram.data\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3674_ wb_override_act net33 _0629_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_136_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6393_ _0350_ clknet_leaf_98_wb_clk_i dffram.data\[41\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5413_ dffram.data\[0\]\[0\] _2022_ _2023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5344_ _1941_ _1971_ _1975_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _1921_ _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4226_ dffram.data\[50\]\[6\] dffram.data\[51\]\[6\] _1007_ _1169_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5681__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ dffram.data\[6\]\[5\] dffram.data\[7\]\[5\] _0669_ _1101_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3108_ net402 _2562_ _2551_ _2565_ _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4236__A2 _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _1029_ _1030_ _1031_ _1032_ _0968_ _0837_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_3039_ _0932_ _0961_ _2503_ _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4881__I _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output274_I net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_147_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A1 _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__I _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 ay8913_do[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput25 ay8913_do[6] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput36 mc14500_do[11] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput69 mc14500_sram_addr[4] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 mc14500_do[21] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput58 mc14500_do[3] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__I _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ wb_counter\[24\] _2795_ _2800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3870__I _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5060_ dffram.data\[25\]\[5\] _1783_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4011_ dffram.data\[46\]\[2\] dffram.data\[47\]\[2\] _0957_ _0958_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5962_ net224 _2391_ _2394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5966__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4913_ dffram.data\[54\]\[3\] _1681_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5893_ _2321_ _2338_ _2341_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ _1634_ _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ dffram.data\[59\]\[6\] _1592_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3729__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4241__I2 _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3726_ _0622_ _0619_ _0639_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__4142__S _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_155_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_155_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6514_ _0471_ clknet_4_8_0_wb_clk_i net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_114_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _0402_ clknet_leaf_52_wb_clk_i dffram.data\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3657_ _2936_ _2975_ _2978_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input172_I sid_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3588_ dffram.data\[60\]\[4\] _2934_ _2935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6376_ _0333_ clknet_leaf_95_wb_clk_i dffram.data\[42\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5327_ _1957_ _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input33_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ _1888_ _1915_ _1918_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5189_ dffram.data\[23\]\[7\] _1868_ _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4209_ dffram.data\[6\]\[6\] dffram.data\[7\]\[6\] _0669_ _1152_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5500__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__A1 _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__S _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4081__B1 _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__I _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4223__I2 _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ net152 _0641_ _1288_ _0717_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_TAPCELL_ROW_41_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_133_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3511_ _2861_ _2883_ _2885_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4491_ _1321_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_123_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3442_ dffram.data\[36\]\[2\] _2836_ _2839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _0187_ clknet_leaf_126_wb_clk_i dffram.data\[23\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__I net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3373_ _2775_ _2783_ _2784_ _2785_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_21_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6161_ _0118_ clknet_leaf_172_wb_clk_i dffram.data\[27\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5112_ _1468_ _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5636__A1 _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6092_ _0049_ clknet_leaf_29_wb_clk_i dffram.data\[59\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5043_ dffram.data\[49\]\[7\] _1770_ _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3742__S0 _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5945_ _2379_ _2380_ _2381_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ dffram.data\[14\]\[4\] _2329_ _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4827_ dffram.data\[6\]\[7\] _1623_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _1504_ _1583_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3709_ _0654_ _0640_ _0643_ _0655_ _0656_ _0657_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_4689_ _1465_ _1532_ _1534_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _0385_ clknet_leaf_64_wb_clk_i dffram.data\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6359_ _0316_ clknet_leaf_90_wb_clk_i dffram.data\[44\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput226 net445 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput215 net502 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput204 sn76489_do[3] net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput237 net459 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput248 net422 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3015__I _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A2 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A1 _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A1 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold3 _2361_ net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _0864_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5730_ dffram.data\[40\]\[2\] _2231_ _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _2142_ _2182_ _2187_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__A1 _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ dffram.data\[43\]\[3\] _2136_ _2143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4612_ _1462_ _1478_ _1479_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4543_ _1422_ _1423_ net344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A1 _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ net184 _1322_ _1361_ net2 _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_96_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ _0170_ clknet_4_8_0_wb_clk_i dffram.data\[52\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3425_ _2452_ _2730_ _2826_ _2827_ _1481_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_40_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6144_ _0101_ clknet_leaf_169_wb_clk_i dffram.data\[54\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3356_ _2614_ _2768_ _2772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6075_ _0032_ clknet_leaf_15_wb_clk_i dffram.data\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3287_ _2522_ wb_counter\[5\] _2709_ _2715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input135_I qcpu_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5026_ _1762_ _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4832__A2 _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6034__A1 net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__I _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_170_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_170_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5928_ _2355_ _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _2276_ _2033_ _2317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3571__A2 _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output354_I net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold89_I wbs_dat_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3011__A1 _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4240__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4198__S0 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4190_ _1019_ _1133_ _1080_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4511__B2 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3210_ net387 _2632_ _2647_ _2652_ _2653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_66_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3141_ _2592_ _2593_ _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_128_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3072_ _2511_ _2533_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A1 net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3974_ _0805_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_75_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5713_ _2216_ _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3250__A1 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5644_ _2144_ _2175_ _2177_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5575_ _2085_ _2126_ _2130_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__S _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4526_ net94 _1411_ _1408_ net15 _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ net177 _1316_ _1317_ net108 net60 _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__4189__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__B2 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__A1 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3408_ net242 _2814_ _2815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4388_ _1249_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6127_ _0084_ clknet_leaf_10_wb_clk_i dffram.data\[56\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3339_ _2757_ _2753_ _2758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6058_ _0015_ clknet_leaf_6_wb_clk_i dffram.data\[31\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _1750_ _1743_ _1751_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4041__I0 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__S _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A1 _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3203__I _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3783__A2 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4034__I _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A1 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _0631_ _0642_ net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4032__I0 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ _1985_ _1986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4732__A1 _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput316 net316 io_oeb[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput305 net305 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput338 net338 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput327 net327 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput349 net349 io_out[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _0625_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5291_ dffram.data\[48\]\[1\] _1937_ _1940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4242_ _1019_ _1184_ _1080_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ dffram.data\[48\]\[5\] dffram.data\[49\]\[5\] _0813_ _1117_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_143_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_407 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_109_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xmultiplexer_418 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_3124_ _2550_ _2579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4799__A1 _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3055_ _2469_ _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3471__A1 _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3957_ _0668_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_34_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3888_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5627_ dffram.data\[42\]\[7\] _2162_ _2166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5558_ _2119_ _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input63_I mc14500_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4509_ net170 _1396_ _1378_ net89 net10 _1393_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_5489_ _2071_ _2064_ _2072_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_137_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output317_I net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3023__I _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3214__A1 net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__C2 _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__A1 _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__A1 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4190__A2 _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_176_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_7_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _1610_ _1651_ _1653_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3811_ dffram.data\[60\]\[0\] dffram.data\[61\]\[0\] _0759_ _0760_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4791_ _1597_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _0487_ clknet_4_10_0_wb_clk_i net379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _0663_ _0667_ _0670_ _0672_ _0682_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_126_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _0418_ clknet_leaf_46_wb_clk_i dffram.data\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3673_ _0628_ wb_override_act _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6392_ _0349_ clknet_leaf_86_wb_clk_i dffram.data\[41\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5412_ _2020_ _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ dffram.data\[21\]\[2\] _1972_ _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _1921_ _1928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4225_ dffram.data\[48\]\[6\] dffram.data\[49\]\[6\] _0813_ _1168_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ dffram.data\[4\]\[5\] dffram.data\[5\]\[5\] _0983_ _1100_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3107_ _2563_ _2564_ _2565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ dffram.data\[30\]\[4\] dffram.data\[31\]\[4\] _0904_ _1032_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3038_ _2476_ _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ dffram.data\[26\]\[5\] _1736_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _0616_ clknet_leaf_72_wb_clk_i dffram.data\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_12_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4402__I _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4172__A2 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output267_I net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__A3 _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3435__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5188__A1 _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4235__I0 _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3738__A2 _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold71_I wbs_dat_i[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4935__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput15 ay8913_do[22] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 ay8913_do[7] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput37 mc14500_do[12] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 mc14500_do[22] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_123_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 mc14500_do[4] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _0781_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5961_ net258 _2386_ _2393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3426__A1 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _1550_ _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5892_ dffram.data\[62\]\[1\] _2339_ _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4843_ _1634_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4774_ _1559_ _1591_ _1594_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3725_ net66 _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _0470_ clknet_leaf_135_wb_clk_i net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6444_ _0401_ clknet_leaf_56_wb_clk_i dffram.data\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3656_ dffram.data\[9\]\[5\] _2976_ _2978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3587_ _2922_ _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6375_ _0332_ clknet_leaf_95_wb_clk_i dffram.data\[42\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _1957_ _1964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input165_I sid_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_124_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5257_ dffram.data\[7\]\[5\] _1916_ _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_54_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4208_ dffram.data\[4\]\[6\] dffram.data\[5\]\[6\] _0983_ _1151_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input26_I ay8913_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1825_ _1867_ _1871_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4139_ _1083_ net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3417__A1 _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3432__A4 _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A1 _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A1 _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__I _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3408__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4307__I _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4908__A1 _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ dffram.data\[33\]\[0\] _2884_ _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _1382_ _1384_ net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_69_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3441_ _2321_ _2835_ _2838_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5333__A1 _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4136__A2 _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3881__I _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3372_ _2370_ _2785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6160_ _0117_ clknet_leaf_172_wb_clk_i dffram.data\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5111_ _1817_ _1818_ _1820_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6091_ _0048_ clknet_4_4_0_wb_clk_i dffram.data\[37\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3647__A1 _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _1758_ _1769_ _1773_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5944_ _2363_ _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5875_ _2317_ _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _1564_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4375__A2 _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _1582_ _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__3992__S _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3708_ _0646_ design_select\[1\] _0624_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_70_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ dffram.data\[30\]\[4\] _1533_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6427_ _0384_ clknet_leaf_75_wb_clk_i dffram.data\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3639_ dffram.data\[61\]\[7\] _2963_ _2967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3791__I _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _0315_ clknet_leaf_91_wb_clk_i dffram.data\[44\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5309_ _1951_ _1946_ _1952_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _0246_ clknet_leaf_110_wb_clk_i dffram.data\[21\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput227 net444 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput216 wbs_adr_i[2] net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput205 sn76489_do[4] net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3638__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput238 net457 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput249 net435 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_92_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4063__S _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold4 net480 net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4238__S _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__I _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3990_ _0933_ _0934_ _0935_ _0936_ _0871_ _0872_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_57_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3876__I _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ dffram.data\[41\]\[3\] _2183_ _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ dffram.data\[5\]\[7\] _1466_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5591_ _2073_ _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4542_ net53 _1325_ _1357_ net20 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4473_ net162 _1344_ _1331_ net81 net35 _1354_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__5306__A1 _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3424_ wb_counter\[31\] _2825_ _2726_ _2827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6212_ _0169_ clknet_leaf_162_wb_clk_i dffram.data\[52\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3116__I _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3355_ _2371_ _2771_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6143_ _0100_ clknet_leaf_175_wb_clk_i dffram.data\[54\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6074_ _0031_ clknet_leaf_15_wb_clk_i dffram.data\[30\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3286_ _2708_ _2713_ _2714_ _2701_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4148__S _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _1762_ _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input128_I qcpu_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5793__A1 _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5927_ net405 _2367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5858_ _1443_ _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input93_I qcpu_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5545__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ dffram.data\[3\]\[6\] _2268_ _2273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4809_ _1547_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4410__I _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5784__A1 _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3890__S0 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__A2 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6099__CLK clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4198__S1 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3140_ net262 _2582_ _2583_ _2593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_128_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3071_ net398 _2518_ _2531_ _2532_ _2533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_82_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5712_ _2204_ _2217_ _2222_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3973_ _0725_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A1 _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ dffram.data\[17\]\[4\] _2176_ _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5574_ dffram.data\[44\]\[6\] _2127_ _2130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4525_ _1341_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4456_ _1323_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4189__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4387_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ _2692_ _2814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3338_ wb_counter\[14\] _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6126_ _0083_ clknet_leaf_178_wb_clk_i dffram.data\[56\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6057_ _0014_ clknet_leaf_6_wb_clk_i dffram.data\[31\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3269_ _2700_ _2701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3069__A2 _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5008_ dffram.data\[53\]\[3\] _1744_ _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5766__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output297_I net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_166_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_79_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__I _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4251__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2991__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__I1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput317 net317 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput306 net306 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput339 net339 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput328 net328 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4310_ net113 _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5290_ _1807_ _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4241_ _1180_ _1181_ _1182_ _1183_ _0785_ _0787_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4985__I _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A1 _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4172_ _0733_ _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_408 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3123_ _2546_ _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3054_ _2511_ _2517_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_149_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_149_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5748__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3956_ dffram.data\[28\]\[2\] dffram.data\[29\]\[2\] _0831_ _0903_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__S _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5626_ _2150_ _2161_ _2165_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3887_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input195_I sn76489_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2982__A1 _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5557_ _1984_ _2118_ _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ dffram.data\[45\]\[2\] _2065_ _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4508_ net192 _1381_ _1375_ net43 _1376_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__3782__I0 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4439_ _1320_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input56_I mc14500_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__A1 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__B2 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _0066_ clknet_leaf_169_wb_clk_i dffram.data\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5987__A1 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5739__A1 _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4411__A1 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4135__I _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__B2 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5911__A1 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__S0 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5978__A1 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3810_ _0736_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4045__I _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4790_ _1597_ _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3741_ _0689_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6460_ _0417_ clknet_leaf_46_wb_clk_i dffram.data\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3672_ wb_rst_override _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_136_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6391_ _0348_ clknet_leaf_94_wb_clk_i dffram.data\[41\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5411_ _2020_ _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _1939_ _1971_ _1974_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5273_ _1882_ _1922_ _1927_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4224_ _0733_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4155_ dffram.data\[2\]\[5\] dffram.data\[3\]\[5\] _0829_ _1099_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3106_ net288 _2553_ _2557_ _2564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4086_ dffram.data\[28\]\[4\] dffram.data\[29\]\[4\] _0831_ _1031_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4156__S _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input110_I qcpu_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3037_ _2472_ _2502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input208_I sn76489_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4988_ _1689_ _1735_ _1737_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3939_ dffram.data\[32\]\[1\] dffram.data\[33\]\[1\] _0793_ _0887_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6658_ _0615_ clknet_leaf_73_wb_clk_i dffram.data\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_46_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _2154_ _2155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6589_ _0546_ clknet_leaf_36_wb_clk_i dffram.data\[35\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5514__I _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3435__A2 _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4632__A1 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3199__A1 net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 ay8913_do[23] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 ay8913_do[8] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput49 mc14500_do[23] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput38 mc14500_do[13] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold64_I wbs_dat_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3371__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4171__I0 _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__A2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ _2389_ _2392_ _2381_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5891_ _2316_ _2338_ _2340_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4911_ _1685_ _1680_ _1686_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _1619_ _1635_ _1640_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ dffram.data\[59\]\[5\] _1592_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3724_ _0647_ _0636_ _0634_ _0625_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6512_ _0469_ clknet_leaf_161_wb_clk_i design_select\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3655_ _2932_ _2975_ _2977_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6443_ _0400_ clknet_leaf_59_wb_clk_i dffram.data\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3586_ _2922_ _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6374_ _0331_ clknet_leaf_95_wb_clk_i dffram.data\[42\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3362__A1 wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _1943_ _1958_ _1963_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input158_I qcpu_sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _1884_ _1915_ _1917_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4207_ dffram.data\[2\]\[6\] dffram.data\[3\]\[6\] _0829_ _1150_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5187_ dffram.data\[23\]\[6\] _1868_ _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4862__A1 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_164_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_164_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ _1055_ _1082_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_3_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input19_I ay8913_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4069_ dffram.data\[36\]\[3\] dffram.data\[37\]\[3\] _0797_ _1015_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__I _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4413__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5244__I _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_100_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A1 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3592__A1 _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4216__S0 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3440_ dffram.data\[36\]\[1\] _2836_ _2838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3371_ net236 _2773_ _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4541__B1 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6090_ _0047_ clknet_leaf_38_wb_clk_i dffram.data\[37\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5110_ dffram.data\[24\]\[4\] _1819_ _1820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5041_ dffram.data\[49\]\[6\] _1770_ _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5097__A1 _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4072__A2 _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5943_ net250 _2377_ _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5874_ _2317_ _2328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ _1627_ _1622_ _1628_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4756_ _1506_ _1437_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _1525_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3707_ net216 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_31_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3638_ _2938_ _2962_ _2966_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6426_ _0383_ clknet_leaf_73_wb_clk_i dffram.data\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _0314_ clknet_leaf_91_wb_clk_i dffram.data\[44\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3569_ _2880_ _2915_ _2920_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3335__A1 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5308_ dffram.data\[48\]\[6\] _1947_ _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6288_ _0245_ clknet_leaf_109_wb_clk_i dffram.data\[21\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput217 wbs_adr_i[3] net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput206 sn76489_do[5] net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5239_ dffram.data\[4\]\[7\] _1902_ _1906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput228 net443 net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput239 net465 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4408__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5260__A1 _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5315__A2 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__A1 dffram.data\[39\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold5 net248 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _1477_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5003__A1 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5590_ _2140_ _2135_ _2141_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3565__A1 _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3892__I _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4541_ net202 _1356_ _1342_ net99 _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4472_ _1369_ _1370_ net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_110_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _0168_ clknet_leaf_115_wb_clk_i dffram.data\[24\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3423_ wb_counter\[31\] _2825_ _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_111_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6142_ _0099_ clknet_leaf_156_wb_clk_i dffram.data\[54\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3354_ net231 _2765_ _2770_ _2771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6073_ _0030_ clknet_leaf_15_wb_clk_i dffram.data\[30\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ net250 _2705_ _2714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5024_ _1664_ _1633_ _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5242__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5926_ _2365_ net427 _2364_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ _2274_ _2310_ _2315_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ _2084_ _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4808_ _1615_ _1612_ _1616_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input86_I qcpu_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4739_ _1539_ _1570_ _1572_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_156_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _0366_ clknet_leaf_83_wb_clk_i dffram.data\[16\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3307__I _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4808__A1 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__S1 _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__S _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3070_ _2464_ _2525_ _2469_ _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_128_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3887__I _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ dffram.data\[16\]\[3\] _2218_ _2222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3972_ _0915_ _0916_ _0917_ _0918_ _0854_ _0690_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_57_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_114_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ _2168_ _2176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _2082_ _2126_ _2129_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3538__A1 _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4524_ net197 _1381_ _1388_ net48 _1337_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _1336_ _1355_ _1358_ net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_123_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4386_ _1297_ _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3406_ _2812_ _2810_ _2813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6125_ _0082_ clknet_leaf_9_wb_clk_i dffram.data\[56\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3337_ wb_counter\[15\] _2756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input140_I qcpu_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__A1 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6056_ _0013_ clknet_leaf_7_wb_clk_i dffram.data\[31\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3268_ _1480_ _2700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3069__A3 _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3199_ net272 _2627_ _2628_ _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5007_ _1550_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3797__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_132_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5766__A2 _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ wb_feedback_delay _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold94_I wbs_dat_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__I2 _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput307 net307 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput329 net329 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput318 net318 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4240_ dffram.data\[46\]\[6\] dffram.data\[47\]\[6\] _0811_ _1183_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4171_ _1111_ _1112_ _1113_ _1114_ _0744_ _0746_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3122_ _2547_ _2577_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_143_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_409 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_93_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3053_ net396 _2470_ _2515_ _2516_ _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3955_ dffram.data\[26\]\[2\] dffram.data\[27\]\[2\] _0829_ _0902_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_34_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5625_ dffram.data\[42\]\[6\] _2162_ _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3886_ _0679_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5337__I _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5556_ _1699_ _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input188_I sn76489_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5487_ _2070_ _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4507_ _1395_ _1397_ net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3782__I1 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _1315_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5684__A1 _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I mc14500_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4369_ net122 _1284_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5436__A1 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6108_ _0065_ clknet_leaf_171_wb_clk_i dffram.data\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6039_ _2441_ _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4416__I _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5911__A2 _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4270__S1 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3230__I _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3740_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4262__S _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3671_ _0620_ _0621_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_82_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5157__I _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6390_ _0347_ clknet_leaf_97_wb_clk_i dffram.data\[41\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5410_ _1907_ _2019_ _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_24_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5341_ dffram.data\[21\]\[1\] _1972_ _1974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ dffram.data\[22\]\[3\] _1923_ _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4223_ _1162_ _1163_ _1164_ _1165_ _0744_ _0746_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_4154_ dffram.data\[0\]\[5\] dffram.data\[1\]\[5\] _0980_ _1098_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5418__A1 _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4085_ dffram.data\[26\]\[4\] dffram.data\[27\]\[4\] _0964_ _1030_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3105_ _2534_ wb_counter\[9\] _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5620__I _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3036_ _1482_ _2501_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input103_I qcpu_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ dffram.data\[26\]\[4\] _1736_ _1737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3938_ _0699_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6657_ _0614_ clknet_leaf_72_wb_clk_i dffram.data\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3869_ _0718_ _0721_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5067__I _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5608_ _2133_ _2090_ _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6588_ _0545_ clknet_leaf_39_wb_clk_i dffram.data\[36\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5539_ _2061_ _2106_ _2108_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_76_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5657__A1 _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_86_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_15_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output322_I net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 ay8913_do[24] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput28 ay8913_do[9] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 mc14500_do[14] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A1 _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5890_ dffram.data\[62\]\[0\] _2339_ _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4910_ dffram.data\[54\]\[2\] _1681_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ dffram.data\[57\]\[3\] _1636_ _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3895__I _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4772_ _1554_ _1591_ _1593_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6511_ _0468_ clknet_leaf_161_wb_clk_i design_select\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3723_ dffram.data\[30\]\[0\] dffram.data\[31\]\[0\] _0671_ _0672_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3654_ dffram.data\[9\]\[4\] _2976_ _2977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6442_ _0399_ clknet_leaf_59_wb_clk_i dffram.data\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5887__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ _0330_ clknet_leaf_94_wb_clk_i dffram.data\[42\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3585_ _1464_ _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5324_ dffram.data\[8\]\[3\] _1959_ _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5255_ dffram.data\[7\]\[4\] _1916_ _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4206_ dffram.data\[0\]\[6\] dffram.data\[1\]\[6\] _0980_ _1149_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4167__S _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5186_ _1822_ _1867_ _1870_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ _1061_ _1068_ _1074_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_3_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4068_ dffram.data\[34\]\[3\] dffram.data\[35\]\[3\] _0946_ _1014_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5811__A1 _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3019_ _2473_ _2478_ _2480_ _2485_ _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_133_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output272_I net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5525__I _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__A1 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__I _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5869__A1 _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4216__S1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6040__B _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__B2 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3370_ wb_counter\[21\] _2782_ _2783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _1756_ _1769_ _1772_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_53_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ net284 _2372_ _2379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5873_ _1464_ _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4824_ dffram.data\[6\]\[6\] _1623_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4514__I _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _1565_ _1576_ _1581_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3706_ net65 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA_clkbuf_leaf_146_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _1525_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3637_ dffram.data\[61\]\[6\] _2963_ _2966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6425_ _0382_ clknet_leaf_75_wb_clk_i dffram.data\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input170_I sid_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _0313_ clknet_leaf_92_wb_clk_i dffram.data\[44\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__S0 _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3568_ dffram.data\[29\]\[7\] _2916_ _2920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4532__B2 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5307_ _1824_ _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_8_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ _0244_ clknet_leaf_106_wb_clk_i dffram.data\[21\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3499_ dffram.data\[34\]\[5\] _2874_ _2877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput218 wbs_adr_i[4] net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput207 sn76489_do[6] net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input31_I blinker_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5238_ _1890_ _1901_ _1905_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput229 net446 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3099__A1 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _1488_ _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6037__A1 net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4424__I _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4523__A1 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold6 _2374_ net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_96_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6028__A1 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4134__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_27_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4540_ _1420_ _1421_ net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4762__A1 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ net210 _1333_ _1361_ net28 _1328_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_64_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6210_ _0167_ clknet_leaf_116_wb_clk_i dffram.data\[24\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3422_ _2670_ wb_counter\[29\] wb_counter\[30\] _2816_ _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XPHY_EDGE_ROW_36_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _0098_ clknet_leaf_175_wb_clk_i dffram.data\[54\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3353_ _2768_ _2769_ _2690_ _2770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6072_ _0029_ clknet_leaf_14_wb_clk_i dffram.data\[30\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3284_ wb_counter\[5\] _2712_ _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_139_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5023_ _1760_ _1753_ _1761_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A1 net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5242__A2 _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5925_ net426 _2360_ _2366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_24_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ dffram.data\[38\]\[7\] _2311_ _2315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4807_ dffram.data\[6\]\[1\] _1613_ _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ _2270_ _2267_ _2271_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4180__S _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2999_ design_select\[4\] _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4753__A1 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ dffram.data\[37\]\[0\] _1571_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input79_I mc14500_sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4669_ dffram.data\[58\]\[6\] _1518_ _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6408_ _0365_ clknet_leaf_89_wb_clk_i dffram.data\[16\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6339_ _0296_ clknet_leaf_81_wb_clk_i dffram.data\[45\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3492__A1 _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4090__S _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__I _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3233__I _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3483__A1 _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4265__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_141_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ dffram.data\[6\]\[2\] dffram.data\[7\]\[2\] _0852_ _0918_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3235__A1 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _2202_ _2217_ _2221_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_18_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5641_ _2168_ _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ dffram.data\[44\]\[5\] _2127_ _2129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4735__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _1406_ _1409_ net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4454_ net205 _1356_ _1357_ net23 _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4385_ _1298_ _1301_ net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5160__A1 _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3405_ wb_counter\[27\] _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6124_ _0081_ clknet_leaf_7_wb_clk_i dffram.data\[56\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3336_ _2752_ _2754_ _2755_ _2747_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6055_ _0012_ clknet_leaf_177_wb_clk_i dffram.data\[31\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input133_I qcpu_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3267_ net245 _2693_ _2699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5006_ _1748_ _1743_ _1749_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3474__A1 dffram.data\[35\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3198_ _2641_ wb_counter\[23\] _2642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4175__S _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4974__A1 _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ net256 _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _2303_ _2305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4041__I3 _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output352_I net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3465__A1 _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_99_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold87_I wbs_dat_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__I3 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput308 net308 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput319 net319 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5443__I _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ dffram.data\[62\]\[5\] dffram.data\[63\]\[5\] _1001_ _1114_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3121_ net373 _2562_ _2551_ _2576_ _2577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_143_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3052_ _0632_ _2489_ _2499_ _2516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3208__A1 net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4956__A1 _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ dffram.data\[24\]\[2\] dffram.data\[25\]\[2\] _0824_ _0901_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3885_ dffram.data\[30\]\[1\] dffram.data\[31\]\[1\] _0669_ _0833_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5624_ _2148_ _2161_ _2164_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5555_ _2088_ _2112_ _2117_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4184__A2 _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_158_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_158_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5486_ _1453_ _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4506_ net169 _1396_ _1388_ net42 net9 _1393_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4437_ net102 _1342_ _1325_ net56 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5133__A1 _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _0064_ clknet_leaf_23_wb_clk_i dffram.data\[63\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4368_ _1287_ _1291_ net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_74_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ dffram.data\[42\]\[7\] dffram.data\[43\]\[7\] _1209_ _1241_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3319_ _2573_ _2738_ _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ net246 _2376_ _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4947__A1 _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_86_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3670_ _0623_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5363__A1 _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ _1934_ _1971_ _1973_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5115__A1 _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5271_ _1880_ _1922_ _1926_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4222_ dffram.data\[62\]\[6\] dffram.data\[63\]\[6\] _1001_ _1165_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4153_ _0908_ _1096_ _1040_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4084_ dffram.data\[24\]\[4\] dffram.data\[25\]\[4\] _0824_ _1029_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3104_ _2561_ _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3429__A1 net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3035_ net382 _2470_ _2498_ _2500_ _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_39_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _1728_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3937_ _0770_ _0884_ _0790_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__I _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__I _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6656_ _0613_ clknet_leaf_75_wb_clk_i dffram.data\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3868_ _0808_ _0810_ _0812_ _0814_ _0815_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_61_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _0544_ clknet_leaf_40_wb_clk_i dffram.data\[36\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5607_ _2152_ _2145_ _2153_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5354__A1 _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3799_ _0719_ _0720_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5538_ dffram.data\[18\]\[0\] _2107_ _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input61_I mc14500_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _2013_ _2054_ _2057_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_55_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_107_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output315_I net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5593__A1 _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__A2 _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 ay8913_do[25] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput29 blinker_do[0] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__I2 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__C2 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__B1 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4273__S _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ _1617_ _1635_ _1639_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_138_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5584__A1 _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4771_ dffram.data\[59\]\[4\] _1592_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5168__I _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _0467_ clknet_leaf_120_wb_clk_i design_select\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_136_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3722_ _0668_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3653_ _2968_ _2976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6441_ _0398_ clknet_leaf_60_wb_clk_i dffram.data\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6372_ _0329_ clknet_leaf_95_wb_clk_i dffram.data\[42\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5887__A2 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4800__I _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3584_ _2930_ _2923_ _2931_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5323_ _1941_ _1958_ _1962_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5254_ _1908_ _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5631__I _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4205_ _0770_ _1147_ _1040_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5185_ dffram.data\[23\]\[5\] _1868_ _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4136_ _1019_ _1079_ _1080_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4247__I _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4067_ dffram.data\[32\]\[3\] dffram.data\[33\]\[3\] _0793_ _1013_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_175_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3018_ _2482_ _2483_ _2484_ _2485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A1 _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__I _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_173_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_173_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4969_ dffram.data\[27\]\[6\] _1722_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_22_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _0596_ clknet_leaf_78_wb_clk_i dffram.data\[19\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_102_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output265_I net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_89_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5318__A1 dffram.data\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4268__S _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3900__S _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5941_ _2375_ _2378_ _2364_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5872_ _2325_ _2318_ _2326_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5557__A1 _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4823_ _1561_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4754_ dffram.data\[37\]\[7\] _1577_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3032__A2 _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5309__A1 _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3705_ net146 _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__4517__C1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _1460_ _1526_ _1531_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3636_ _2936_ _2962_ _2965_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6424_ _0381_ clknet_leaf_75_wb_clk_i dffram.data\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _0312_ clknet_leaf_79_wb_clk_i dffram.data\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3966__S1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3567_ _2878_ _2915_ _2919_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6286_ _0243_ clknet_leaf_106_wb_clk_i dffram.data\[21\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5306_ _1949_ _1946_ _1950_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input163_I sid_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5237_ dffram.data\[4\]\[6\] _1902_ _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3498_ _1469_ _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput208 sn76489_do[7] net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput219 wbs_adr_i[5] net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input24_I ay8913_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5168_ _1857_ _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5099_ _1810_ _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4119_ dffram.data\[52\]\[4\] dffram.data\[53\]\[4\] _0878_ _1064_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output382_I net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5720__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold7 net513 net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A1 _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4134__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ net181 _1316_ _1317_ net112 net64 _1359_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ _2765_ _2823_ _2824_ _2541_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3352_ wb_counter\[16\] _2761_ wb_counter\[17\] _2769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6140_ _0097_ clknet_leaf_175_wb_clk_i dffram.data\[54\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5181__I _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3283_ _2522_ _2709_ _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6071_ _0028_ clknet_leaf_11_wb_clk_i dffram.data\[30\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5022_ dffram.data\[53\]\[7\] _1754_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__I _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ net268 _2357_ _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _2272_ _2310_ _2314_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4806_ _1544_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_111_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5786_ dffram.data\[3\]\[5\] _2268_ _2271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2998_ _2464_ _2458_ _2465_ _2466_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4737_ _1569_ _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5950__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4668_ _1470_ _1517_ _1520_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6407_ _0364_ clknet_leaf_89_wb_clk_i dffram.data\[16\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3619_ _2940_ _2949_ _2954_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5702__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6338_ _0295_ clknet_leaf_82_wb_clk_i dffram.data\[45\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6269_ _0226_ clknet_leaf_120_wb_clk_i dffram.data\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__I _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_141_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4432__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ dffram.data\[4\]\[2\] dffram.data\[5\]\[2\] _0728_ _0917_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_48_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4281__S _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2994__A1 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _2142_ _2169_ _2174_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5571_ _2077_ _2126_ _2128_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4522_ net47 _1407_ _1408_ net14 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3794__I0 dffram.data\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4453_ _1349_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__A1 _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3404_ _2807_ _2811_ _2451_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4384_ net129 _1294_ _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6123_ _0080_ clknet_leaf_27_wb_clk_i dffram.data\[57\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3335_ net228 _2750_ _2755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ wb_counter\[2\] _2697_ _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6054_ _0011_ clknet_leaf_177_wb_clk_i dffram.data\[31\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_0_Left_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5005_ dffram.data\[53\]\[2\] _1744_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3197_ _2571_ _2641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input126_I qcpu_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5907_ _2335_ _2344_ _2349_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4974__A2 _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ _2303_ _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input91_I qcpu_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ dffram.data\[3\]\[0\] _2258_ _2259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3162__A1 _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold2_I net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4662__A1 _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3509__I _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__I _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput309 net309 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3120_ _2574_ _2575_ _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4276__S _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3051_ _2502_ _2512_ _2513_ _2514_ _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3839__S0 _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3953_ _0900_ net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_63_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4803__I _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3884_ dffram.data\[28\]\[1\] dffram.data\[29\]\[1\] _0831_ _0832_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ dffram.data\[42\]\[5\] _2162_ _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3767__I0 _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ dffram.data\[18\]\[7\] _2113_ _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5381__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5485_ _2068_ _2064_ _2069_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _1330_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4436_ _1341_ _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4367_ _1290_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6106_ _0063_ clknet_leaf_24_wb_clk_i dffram.data\[63\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_127_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3318_ _2573_ _2738_ _2741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4298_ dffram.data\[40\]\[7\] dffram.data\[41\]\[7\] _0827_ _1240_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4186__S _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4644__A1 _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3249_ _2482_ wb_counter\[31\] _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6037_ net280 _2368_ _2449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output295_I net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__S0 _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3329__I _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__B1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__C2 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__I0 _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3135__A1 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A1 _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_72_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_31_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__I _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_81_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5270_ dffram.data\[22\]\[2\] _1923_ _1926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4221_ dffram.data\[60\]\[6\] dffram.data\[61\]\[6\] _0737_ _1164_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4874__A1 _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3903__S _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4152_ _1092_ _1093_ _1094_ _1095_ _0976_ _0977_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_4083_ _1028_ net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3103_ _2490_ _2561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3034_ _0628_ _2489_ _2499_ _2500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_90_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_165_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5051__A1 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _1728_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3936_ _0876_ _0877_ _0879_ _0880_ _0881_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_74_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6655_ _0612_ clknet_leaf_55_wb_clk_i dffram.data\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3867_ _0786_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input193_I sn76489_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3798_ _0735_ _0738_ _0741_ _0743_ _0744_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6586_ _0543_ clknet_leaf_40_wb_clk_i dffram.data\[36\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5606_ dffram.data\[43\]\[7\] _2146_ _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5537_ _2105_ _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input54_I mc14500_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ dffram.data\[1\]\[5\] _2055_ _2057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4419_ _0637_ net32 _0652_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5399_ _2009_ _2010_ _2012_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4708__I _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_107_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output308_I net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5042__A1 _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 ay8913_do[26] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_138_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5274__I _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3723__S _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__B2 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A1 _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3595__A1 _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _1584_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3721_ dffram.data\[28\]\[0\] dffram.data\[29\]\[0\] _0669_ _0670_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3652_ _2968_ _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6440_ _0397_ clknet_leaf_49_wb_clk_i dffram.data\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5336__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3583_ dffram.data\[60\]\[3\] _2924_ _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _0328_ clknet_leaf_96_wb_clk_i dffram.data\[43\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5322_ dffram.data\[8\]\[2\] _1959_ _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5253_ _1908_ _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4204_ _1143_ _1144_ _1145_ _1146_ _0976_ _0977_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_5184_ _1817_ _1867_ _1869_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_71_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4135_ _0818_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _1005_ _1011_ _0790_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3017_ _2455_ _2484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input206_I sn76489_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ _1693_ _1721_ _1724_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3919_ dffram.data\[58\]\[1\] dffram.data\[59\]\[1\] _0757_ _0867_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4899_ _1629_ _1672_ _1677_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6638_ _0595_ clknet_leaf_79_wb_clk_i dffram.data\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4535__B1 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5094__I _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_142_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_142_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6569_ _0526_ clknet_leaf_147_wb_clk_i wb_counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output258_I net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__A1 _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4066__A2 _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3718__S _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold62_I wbs_dat_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4348__I _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5940_ net249 _2377_ _2378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4462__C1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4083__I _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5871_ dffram.data\[14\]\[3\] _2319_ _2326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A1 _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5557__A2 _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ _1625_ _1622_ _1626_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4753_ _1562_ _1576_ _1580_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3568__A1 dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3704_ _0630_ _0653_ net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_83_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6423_ _0380_ clknet_leaf_55_wb_clk_i dffram.data\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4684_ dffram.data\[30\]\[3\] _1527_ _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ dffram.data\[61\]\[5\] _2963_ _2965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4517__C2 _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6354_ _0311_ clknet_leaf_84_wb_clk_i dffram.data\[18\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3566_ dffram.data\[29\]\[6\] _2916_ _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5642__I _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6285_ _0242_ clknet_leaf_106_wb_clk_i dffram.data\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3497_ _2872_ _2873_ _2875_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5305_ dffram.data\[48\]\[5\] _1947_ _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input156_I qcpu_sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5236_ _1888_ _1901_ _1904_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput209 sn76489_do[8] net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5493__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5167_ _1429_ _0722_ _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _1453_ _1810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4118_ dffram.data\[50\]\[4\] dffram.data\[51\]\[4\] _1007_ _1063_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input17_I ay8913_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ _0921_ _0994_ _0750_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4194__S _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3559__A1 _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3949__I3 _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold8 net234 net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5236__A1 _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3420_ net246 _2814_ _2824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ _2767_ _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I ay8913_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3282_ _2708_ _2710_ _2711_ _2701_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_29_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6070_ _0027_ clknet_leaf_176_wb_clk_i dffram.data\[30\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3911__S _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5021_ _1564_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__I _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ _2358_ net421 _2364_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ dffram.data\[38\]\[6\] _2311_ _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_66_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4805_ _1610_ _1612_ _1614_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5785_ _2081_ _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2997_ _2441_ _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4736_ _1569_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4667_ dffram.data\[58\]\[5\] _1518_ _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6406_ _0363_ clknet_leaf_88_wb_clk_i dffram.data\[16\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3618_ dffram.data\[19\]\[7\] _2950_ _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5702__A2 _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6337_ _0294_ clknet_leaf_81_wb_clk_i dffram.data\[45\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4598_ net250 _1451_ _1457_ net158 _1452_ net77 _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_101_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3549_ _1727_ _2062_ _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_110_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6268_ _0225_ clknet_leaf_119_wb_clk_i dffram.data\[48\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5219_ _1892_ _1885_ _1893_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6199_ _0156_ clknet_leaf_12_wb_clk_i dffram.data\[39\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3952__A1 _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4099__S _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5457__A1 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__I _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3530__I _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ dffram.data\[44\]\[4\] _2127_ _2128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_61_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4521_ _1349_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _1321_ _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3403_ _2726_ _2808_ _2810_ _2811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_102_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4383_ _1298_ _1300_ net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3705__I net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5448__A1 _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6122_ _0079_ clknet_leaf_27_wb_clk_i dffram.data\[57\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3334_ wb_counter\[14\] _2753_ _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5920__I _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3265_ _2483_ _2496_ _2697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6053_ _0010_ clknet_leaf_10_wb_clk_i dffram.data\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5004_ _1547_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_68_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3196_ _2624_ _2640_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input119_I qcpu_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5906_ dffram.data\[62\]\[7\] _2345_ _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5837_ _1568_ _2033_ _2303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_101_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5768_ _2256_ _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ dffram.data\[2\]\[4\] _1556_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input84_I qcpu_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ _2087_ _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_112_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__A1 _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_112_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_110_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5678__A1 _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_143_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3050_ _2506_ wb_counter\[3\] _2484_ _2514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_155_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4405__A2 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4292__S _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3839__S1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3952_ _0863_ _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3883_ _0665_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5622_ _2144_ _2161_ _2163_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5553_ _2085_ _2112_ _2116_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__I1 _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ net191 _1385_ _1386_ net88 _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_42_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5484_ dffram.data\[45\]\[1\] _2065_ _2069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5669__A1 _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4435_ _1248_ _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_1_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4366_ _1288_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6105_ _0062_ clknet_leaf_24_wb_clk_i dffram.data\[63\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3317_ _2732_ _2739_ _2740_ _2718_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4297_ _0769_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3248_ _2668_ _2684_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6036_ _2447_ _2448_ _2442_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5841__A1 _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_167_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_167_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3179_ _2619_ wb_counter\[20\] _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4255__S1 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output288_I net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__B2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5832__A1 _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold92_I wbs_dat_i[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3071__A1 net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_136_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5735__I _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__A1 dffram.data\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ dffram.data\[58\]\[6\] dffram.data\[59\]\[6\] _0998_ _1163_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4151_ dffram.data\[22\]\[5\] dffram.data\[23\]\[5\] _0709_ _1095_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4287__S _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ _0996_ _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3102_ _2547_ _2560_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3033_ _2490_ _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _1687_ _1729_ _1734_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3935_ _0882_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6654_ _0611_ clknet_leaf_56_wb_clk_i dffram.data\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ _0784_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5605_ _2087_ _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3797_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6585_ _0542_ clknet_leaf_40_wb_clk_i dffram.data\[36\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5536_ _2105_ _2106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4562__A1 _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3365__A2 wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input186_I sn76489_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5467_ _2009_ _2054_ _2056_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4418_ net29 _1279_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input47_I mc14500_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5398_ dffram.data\[20\]\[4\] _2011_ _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4349_ _0634_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4197__S _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__I _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6019_ net274 _2433_ _2436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3053__A1 net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__A1 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4856__A2 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3903__I1 dffram.data\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__A1 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A2 _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3044__A1 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3720_ _0668_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_28_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _2930_ _2969_ _2974_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__I _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__A1 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__B2 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3582_ _1459_ _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6370_ _0327_ clknet_leaf_99_wb_clk_i dffram.data\[43\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _1939_ _1958_ _1961_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5252_ _1882_ _1909_ _1914_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4203_ dffram.data\[22\]\[6\] dffram.data\[23\]\[6\] _0709_ _1146_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5183_ dffram.data\[23\]\[4\] _1868_ _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3713__I _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4809__I _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _1075_ _1076_ _1077_ _1078_ _0785_ _0787_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_74_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4065_ _1006_ _1008_ _1009_ _1010_ _0881_ _0883_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3016_ wb_counter\[0\] _2483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5024__A2 _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input101_I qcpu_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3035__A1 net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4967_ dffram.data\[27\]\[5\] _1722_ _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4783__A1 _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ dffram.data\[55\]\[7\] _1673_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3918_ dffram.data\[56\]\[1\] dffram.data\[57\]\[1\] _0865_ _0866_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6637_ _0594_ clknet_leaf_78_wb_clk_i dffram.data\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3849_ dffram.data\[36\]\[0\] dffram.data\[37\]\[0\] _0797_ _0798_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__B2 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _0525_ clknet_leaf_147_wb_clk_i wb_counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5519_ _2068_ _2092_ _2095_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__S _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6499_ _0456_ clknet_leaf_144_wb_clk_i net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_89_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output320_I net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A2 _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__S0 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3026__A1 net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4774__A1 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4526__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__B2 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold55_I wbs_adr_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4462__B1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _1459_ _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ dffram.data\[6\]\[5\] _1623_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ dffram.data\[37\]\[6\] _1577_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3703_ _0621_ _0652_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4683_ _1455_ _1526_ _1530_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6422_ _0379_ clknet_leaf_55_wb_clk_i dffram.data\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3634_ _2932_ _2962_ _2964_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4517__A1 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__B2 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _0310_ clknet_leaf_81_wb_clk_i dffram.data\[18\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A1 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3565_ _2876_ _2915_ _2918_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5304_ _1821_ _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6284_ _0241_ clknet_leaf_107_wb_clk_i dffram.data\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3496_ dffram.data\[34\]\[4\] _2874_ _2875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5235_ dffram.data\[4\]\[5\] _1902_ _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input149_I qcpu_sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5166_ _1828_ _1851_ _1856_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4117_ dffram.data\[48\]\[4\] dffram.data\[49\]\[4\] _0875_ _1062_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5097_ _1808_ _1804_ _1809_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4048_ _0989_ _0990_ _0992_ _0993_ _0928_ _0929_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_78_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5999_ _2420_ _2421_ _2419_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__I3 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A1 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4508__B2 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output270_I net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output368_I net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput290 net290 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xhold9 _2366_ net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_96_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4047__I0 dffram.data\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4912__I _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3350_ _2757_ _2756_ _2753_ _2766_ _2767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_110_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5020_ _1758_ _1753_ _1759_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3281_ net249 _2705_ _2711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3486__A1 _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4295__S _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5922_ _2363_ _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ _2270_ _2310_ _2313_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5918__I _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5784_ _2266_ _2267_ _2269_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4804_ dffram.data\[6\]\[0\] _1613_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4735_ _1568_ _1439_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_72_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2996_ net250 _2462_ _2465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _1465_ _1517_ _1519_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _0362_ clknet_leaf_92_wb_clk_i dffram.data\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3617_ _2938_ _2949_ _2953_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5653__I _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4210__I0 _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _1462_ _1465_ _1467_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6336_ _0293_ clknet_leaf_90_wb_clk_i dffram.data\[45\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3548_ _2880_ _2902_ _2907_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3479_ _2847_ _2090_ _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6267_ _0224_ clknet_leaf_107_wb_clk_i dffram.data\[22\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5218_ dffram.data\[50\]\[7\] _1886_ _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6198_ _0155_ clknet_leaf_13_wb_clk_i dffram.data\[39\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3901__I _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ dffram.data\[51\]\[0\] _1846_ _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3348__I _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5154__A1 _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_145_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4968__A1 _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3640__A1 _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _1354_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4451_ net176 _1344_ _1331_ net107 net59 _1354_ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__5145__A1 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _2802_ _2795_ _2809_ _2810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_141_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4382_ net128 _1294_ _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6121_ _0078_ clknet_leaf_27_wb_clk_i dffram.data\[57\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3333_ wb_counter\[11\] wb_counter\[12\] wb_counter\[13\] _2737_ _2753_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3264_ _2691_ _2695_ _2696_ _2466_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6052_ _0009_ clknet_leaf_10_wb_clk_i dffram.data\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4817__I _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5003_ _1746_ _1743_ _1747_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3195_ net385 _2632_ _2625_ _2639_ _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5905_ _2333_ _2344_ _2348_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5836_ _2274_ _2297_ _2302_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5767_ _2256_ _2257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ _2212_ _2207_ _2213_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4718_ _1540_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input77_I mc14500_sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4649_ net211 _0666_ _1434_ _1435_ _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_79_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5383__I _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6319_ _0276_ clknet_leaf_101_wb_clk_i dffram.data\[46\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_92_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_89_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_18_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3631__I _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output400_I net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5558__I _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A1 _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _0874_ _0885_ _0892_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3613__A1 _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3882_ dffram.data\[26\]\[1\] dffram.data\[27\]\[1\] _0829_ _0830_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ dffram.data\[42\]\[4\] _2162_ _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5552_ dffram.data\[18\]\[6\] _2113_ _2116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4503_ _1392_ _1394_ net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _2067_ _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3716__I _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4434_ _1337_ _1339_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4365_ _0627_ _0653_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6104_ _0061_ clknet_leaf_38_wb_clk_i dffram.data\[63\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3316_ net224 _2721_ _2740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4296_ _1234_ _1235_ _1236_ _1237_ _1196_ _0786_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_6035_ net244 _2376_ _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input131_I qcpu_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3247_ net394 _2491_ _2669_ _2683_ _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3178_ _2550_ _2625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_136_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_136_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_135_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ dffram.data\[13\]\[0\] _2292_ _2293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3827__S _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output350_I net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__A2 _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3071__A2 _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold85_I wbs_dat_i[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ dffram.data\[20\]\[5\] dffram.data\[21\]\[5\] _0809_ _1094_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3101_ net401 _2518_ _2551_ _2559_ _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4081_ _1004_ _1012_ _1018_ _1026_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4367__I _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput190 sn76489_do[16] net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3032_ _2473_ _2494_ _2495_ _2497_ _2498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_76_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4229__I3 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5587__A1 _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4983_ dffram.data\[26\]\[3\] _1730_ _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3934_ _0687_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6653_ _0610_ clknet_leaf_55_wb_clk_i dffram.data\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3865_ dffram.data\[46\]\[0\] dffram.data\[47\]\[0\] _0813_ _0814_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5604_ _2150_ _2145_ _2151_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6584_ _0541_ clknet_leaf_43_wb_clk_i dffram.data\[36\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3796_ _0688_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5535_ _2104_ _2090_ _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3446__I _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ dffram.data\[1\]\[4\] _2055_ _2056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input179_I sid_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5511__A1 _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4417_ _1324_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ _1999_ _2011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4348_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4279_ _1198_ _1206_ _1213_ _1220_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_107_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6018_ _2434_ _2435_ _2430_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output398_I net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5750__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4553__A2 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3091__I _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3292__A2 wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3650_ dffram.data\[9\]\[3\] _2970_ _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _2928_ _2923_ _2929_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5741__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ dffram.data\[8\]\[1\] _1959_ _1961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4298__S _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ dffram.data\[7\]\[3\] _1910_ _1914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4202_ dffram.data\[20\]\[6\] dffram.data\[21\]\[6\] _0809_ _1145_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5182_ _1860_ _1868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4133_ dffram.data\[46\]\[4\] dffram.data\[47\]\[4\] _0957_ _1078_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4064_ dffram.data\[54\]\[3\] dffram.data\[55\]\[3\] _0782_ _1010_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3015_ _2481_ _2482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _1689_ _1721_ _1723_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3917_ _0753_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4897_ _1627_ _1672_ _1676_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6636_ _0593_ clknet_leaf_48_wb_clk_i dffram.data\[60\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3848_ _0761_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3779_ _0665_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4535__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6567_ _0524_ clknet_leaf_147_wb_clk_i wb_counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5518_ dffram.data\[10\]\[1\] _2093_ _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_131_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _0455_ clknet_leaf_144_wb_clk_i net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5449_ dffram.data\[46\]\[6\] _2042_ _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3904__I _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__A1 _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4146__S1 _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output313_I net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__A1 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_151_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_151_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4471__B2 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__A1 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A1 _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4462__A1 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4462__B2 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4820_ _1558_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_34_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4065__I1 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4751_ _1559_ _1576_ _1579_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_78_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_90_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ _0648_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_71_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4682_ dffram.data\[30\]\[2\] _1527_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6421_ _0378_ clknet_leaf_52_wb_clk_i dffram.data\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3633_ dffram.data\[61\]\[4\] _2963_ _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ _0309_ clknet_leaf_83_wb_clk_i dffram.data\[18\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3564_ dffram.data\[29\]\[5\] _2916_ _2918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6283_ _0240_ clknet_leaf_69_wb_clk_i dffram.data\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3495_ _2862_ _2874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5303_ _1945_ _1946_ _1948_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5234_ _1884_ _1901_ _1903_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5165_ dffram.data\[51\]\[7\] _1852_ _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4116_ _0864_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ dffram.data\[24\]\[1\] _1805_ _1809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4047_ dffram.data\[14\]\[3\] dffram.data\[15\]\[3\] _0926_ _0993_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input211_I wb_rst_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ net233 _2415_ _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _1695_ _1708_ _1712_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5953__A1 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _0576_ clknet_leaf_2_wb_clk_i dffram.data\[32\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output263_I net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput280 net280 custom_settings[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput291 net291 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_96_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_135_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3247__A2 _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_174_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3280_ _2522_ _2709_ _2710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4683__A1 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5921_ _2362_ _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5852_ dffram.data\[38\]\[5\] _2311_ _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4038__I1 dffram.data\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ dffram.data\[3\]\[4\] _2268_ _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3719__I _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__A1 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4803_ _1611_ _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4734_ _1567_ _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2995_ design_select\[3\] _2464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_127_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4665_ dffram.data\[58\]\[4\] _1518_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ _0361_ clknet_leaf_89_wb_clk_i dffram.data\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3616_ dffram.data\[19\]\[6\] _2950_ _2953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4596_ dffram.data\[5\]\[4\] _1466_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _0292_ clknet_leaf_90_wb_clk_i dffram.data\[45\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3547_ dffram.data\[32\]\[7\] _2903_ _2907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input161_I sid_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_110_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3478_ _1443_ _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6266_ _0223_ clknet_leaf_107_wb_clk_i dffram.data\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5217_ _1827_ _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6197_ _0154_ clknet_leaf_11_wb_clk_i dffram.data\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input22_I ay8913_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _1844_ _1846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5079_ dffram.data\[39\]\[4\] _1796_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2988__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A2 _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4268__I1 dffram.data\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4923__I _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5917__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3539__I _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4450_ _1323_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_80_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4381_ _1298_ _1299_ net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3156__A1 _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3401_ wb_counter\[25\] wb_counter\[26\] _2809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6120_ _0077_ clknet_leaf_5_wb_clk_i dffram.data\[57\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3332_ _2707_ _2752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3274__I _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4656__A1 _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3263_ net234 _2693_ _2696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6051_ _0008_ clknet_leaf_134_wb_clk_i wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3194_ _2637_ _2638_ _2639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5002_ dffram.data\[53\]\[1\] _1744_ _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 dffram.data\[39\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5904_ dffram.data\[62\]\[6\] _2345_ _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4833__I _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ dffram.data\[13\]\[7\] _2298_ _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ _1907_ _2195_ _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5697_ dffram.data\[11\]\[6\] _2208_ _2213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4717_ _1540_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4648_ _0682_ _1505_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _0644_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3942__I0 dffram.data\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__A1 _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ _0275_ clknet_leaf_101_wb_clk_i dffram.data\[46\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_92_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6249_ _0206_ clknet_leaf_68_wb_clk_i dffram.data\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_58_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5072__A1 _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_33_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_133_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3094__I _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4350__A3 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4638__A1 _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold90 wbs_dat_i[19] net508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5063__A1 _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ _0806_ _0897_ _0819_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3881_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_73_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5620_ _2154_ _2162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _2082_ _2112_ _2115_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_51_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4502_ net168 _1383_ _1378_ net87 net8 _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__3767__I3 _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5482_ _1447_ _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3129__A1 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4433_ _1327_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4364_ _0636_ _0635_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6103_ _0060_ clknet_leaf_36_wb_clk_i dffram.data\[63\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4295_ dffram.data\[38\]\[7\] dffram.data\[39\]\[7\] _1192_ _1237_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3732__I _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3315_ _2735_ _2738_ _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3246_ _2681_ _2682_ _2683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6034_ net278 _2368_ _2447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3177_ _2546_ _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input124_I qcpu_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4101__I0 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4801__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _2290_ _2292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ dffram.data\[12\]\[1\] _2244_ _2246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_176_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_176_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_143_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_105_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4183__I3 _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3642__I _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4096__A2 _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5569__I _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A1 _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold78_I wbs_dat_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3817__I _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3100_ _2552_ _2558_ _2559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4080_ _1019_ _1025_ _0819_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput180 sid_do[8] net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3031_ _2482_ _2496_ _2484_ _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput191 sn76489_do[17] net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5479__I _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3598__A1 _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _1685_ _1729_ _1733_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3933_ _0784_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3928__S _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6652_ _0609_ clknet_leaf_47_wb_clk_i dffram.data\[61\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3864_ _0771_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5603_ dffram.data\[43\]\[6\] _2146_ _2151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _0540_ clknet_leaf_43_wb_clk_i dffram.data\[36\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3795_ _0681_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _1857_ _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3770__A1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5465_ _2047_ _2055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_76_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _1999_ _2010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4347_ _1248_ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4278_ _1188_ _1219_ _0749_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_107_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3229_ _2363_ _2668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6017_ net239 _2426_ _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5027__A1 dffram.data\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3589__A1 _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__B1 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output293_I net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3513__A1 _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_73_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_116_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3580_ dffram.data\[60\]\[2\] _2924_ _2929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_125_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5250_ _1880_ _1909_ _1913_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4201_ dffram.data\[18\]\[6\] dffram.data\[19\]\[6\] _0972_ _1144_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4378__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5181_ _1860_ _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_71_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4132_ dffram.data\[44\]\[4\] dffram.data\[45\]\[4\] _1022_ _1077_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4063_ dffram.data\[52\]\[3\] dffram.data\[53\]\[3\] _0878_ _1009_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3014_ net214 _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5009__A1 _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4965_ dffram.data\[27\]\[4\] _1722_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _0695_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ dffram.data\[55\]\[6\] _1673_ _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _0592_ clknet_leaf_50_wb_clk_i dffram.data\[60\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3847_ dffram.data\[34\]\[0\] dffram.data\[35\]\[0\] _0795_ _0796_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3778_ dffram.data\[2\]\[0\] dffram.data\[3\]\[0\] _0666_ _0727_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6566_ _0523_ clknet_leaf_146_wb_clk_i wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_6_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input191_I sn76489_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _2061_ _2092_ _2094_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3743__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5672__I _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6497_ _0454_ clknet_leaf_142_wb_clk_i net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input52_I mc14500_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _2013_ _2041_ _2044_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5379_ _1953_ _1992_ _1997_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5248__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3920__I _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output306_I net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5420__A1 _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_120_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5723__A2 _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_164_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__I _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3830__I _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4750_ dffram.data\[37\]\[5\] _1577_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3701_ _0630_ _0651_ net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4681_ _1449_ _1526_ _1529_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6420_ _0377_ clknet_leaf_55_wb_clk_i dffram.data\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3632_ _2955_ _2963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6351_ _0308_ clknet_leaf_80_wb_clk_i dffram.data\[18\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3725__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5302_ dffram.data\[48\]\[4\] _1947_ _1948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3563_ _2872_ _2915_ _2917_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6282_ _0239_ clknet_leaf_72_wb_clk_i dffram.data\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3494_ _2862_ _2873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ dffram.data\[4\]\[4\] _1902_ _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5164_ _1825_ _1851_ _1855_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4115_ _1056_ _1057_ _1058_ _1059_ _0871_ _0872_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_120_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3740__I _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5095_ _1807_ _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4046_ dffram.data\[12\]\[3\] dffram.data\[13\]\[3\] _0991_ _0992_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5650__A1 _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input204_I sn76489_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4205__A2 _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__A1 _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ net267 _2411_ _2420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4948_ dffram.data\[28\]\[6\] _1709_ _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5953__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4879_ _1664_ _1489_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _0575_ clknet_leaf_3_wb_clk_i dffram.data\[32\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6549_ _0506_ clknet_leaf_158_wb_clk_i wb_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5469__A1 _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput270 net270 custom_settings[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3851__S _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput281 net281 custom_settings[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput292 net292 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4746__I _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3097__I _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A1 _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3560__I _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _1480_ _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_88_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5487__I _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5851_ _2266_ _2310_ _2312_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5782_ _2256_ _2268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4802_ _1611_ _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2994_ _0647_ _2458_ _2463_ _2454_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4733_ _1429_ _0818_ _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6403_ _0360_ clknet_leaf_75_wb_clk_i dffram.data\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4664_ _1510_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3615_ _2936_ _2949_ _2952_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4595_ _1440_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6334_ _0291_ clknet_leaf_91_wb_clk_i dffram.data\[45\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3546_ _2878_ _2902_ _2906_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6265_ _0222_ clknet_leaf_107_wb_clk_i dffram.data\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input154_I qcpu_sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3477_ _2335_ _2855_ _2860_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5216_ _1890_ _1885_ _1891_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__A1 dffram.data\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _0153_ clknet_leaf_12_wb_clk_i dffram.data\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5147_ _1844_ _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4566__I _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _1788_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input15_I ay8913_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ dffram.data\[22\]\[3\] dffram.data\[23\]\[3\] _0711_ _0975_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5397__I _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4362__A1 _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5862__A1 dffram.data\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5917__A2 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4380_ net127 _1294_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3400_ wb_counter\[25\] _2803_ wb_counter\[26\] _2808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3331_ _2732_ _2749_ _2751_ _2747_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6050_ _0007_ clknet_leaf_19_wb_clk_i dffram.data\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3262_ _2483_ _2496_ _2695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input7_I ay8913_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3193_ net271 _2627_ _2628_ _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5001_ _1544_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_68_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5903_ _2331_ _2344_ _2347_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5834_ _2272_ _2297_ _2301_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_17_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ _2060_ _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5696_ _2084_ _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4592__B2 net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _1553_ _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _1088_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_60_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4344__A1 _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4578_ _1311_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6317_ _0274_ clknet_leaf_102_wb_clk_i dffram.data\[46\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_92_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3942__I1 dffram.data\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3529_ _2895_ _2896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6248_ _0205_ clknet_leaf_114_wb_clk_i dffram.data\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6179_ _0136_ clknet_leaf_117_wb_clk_i dffram.data\[53\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3083__A1 _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_98_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_36_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_27_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6021__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4583__A1 dffram.data\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__S _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5835__A1 dffram.data\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold91 wbs_dat_i[20] net509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold80 wbs_dat_i[30] net498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_89_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3074__A1 _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__A1 net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5765__I _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5550_ dffram.data\[18\]\[5\] _2113_ _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _2061_ _2064_ _2066_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4501_ _0650_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ net31 _1279_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4363_ net121 _1268_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ _0059_ clknet_leaf_36_wb_clk_i dffram.data\[63\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4294_ dffram.data\[36\]\[7\] dffram.data\[37\]\[7\] _1192_ _1236_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3314_ _2737_ _2738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5826__A1 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _2445_ _2446_ _2442_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3245_ net280 _2672_ _2673_ _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3176_ _2601_ _2623_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4844__I _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input117_I qcpu_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__A2 _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5817_ _2290_ _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4014__B1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _2194_ _2243_ _2245_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4565__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input82_I qcpu_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5679_ _2067_ _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_103_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_145_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_145_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4020__S _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output336_I net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3056__A1 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__A2 _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__I _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3833__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput170 sid_do[18] net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput181 sid_do[9] net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3295__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ wb_counter\[1\] _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput192 sn76489_do[18] net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_19_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4981_ dffram.data\[26\]\[2\] _1730_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__A1 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ dffram.data\[54\]\[1\] dffram.data\[55\]\[1\] _0782_ _0880_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3863_ dffram.data\[44\]\[0\] dffram.data\[45\]\[0\] _0811_ _0812_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6651_ _0608_ clknet_4_5_0_wb_clk_i dffram.data\[61\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5602_ _2084_ _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4105__S _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _0539_ clknet_leaf_42_wb_clk_i dffram.data\[36\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5533_ _2088_ _2098_ _2103_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3794_ dffram.data\[14\]\[0\] dffram.data\[15\]\[0\] _0742_ _0743_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5464_ _2047_ _2054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4415_ _0683_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5395_ _1816_ _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4346_ _1271_ _1275_ net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4277_ _1214_ _1215_ _1217_ _1218_ _0834_ _0882_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4158__S0 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6016_ net273 _2433_ _2434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3228_ _2646_ _2667_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4574__I net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3159_ _2561_ _2609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4538__B2 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_154_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3653__I _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__A1 _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3029__A1 net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold90_I wbs_dat_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ dffram.data\[16\]\[6\] dffram.data\[17\]\[6\] _0742_ _1143_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _1814_ _1861_ _1866_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_71_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4131_ dffram.data\[42\]\[4\] dffram.data\[43\]\[4\] _0954_ _1076_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4062_ dffram.data\[50\]\[3\] dffram.data\[51\]\[3\] _1007_ _1008_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3013_ net257 _2479_ _2480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4768__A1 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4964_ _1714_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _0839_ _0847_ _0856_ _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_73_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4895_ _1625_ _1672_ _1675_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6634_ _0591_ clknet_leaf_50_wb_clk_i dffram.data\[60\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3991__A2 _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3846_ _0756_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ dffram.data\[0\]\[0\] dffram.data\[1\]\[0\] _0662_ _0726_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6565_ _0522_ clknet_leaf_146_wb_clk_i wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5516_ dffram.data\[10\]\[0\] _2093_ _2094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6496_ _0453_ clknet_leaf_142_wb_clk_i net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input184_I sn76489_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ dffram.data\[46\]\[5\] _2042_ _2044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4569__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5378_ dffram.data\[47\]\[7\] _1993_ _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input45_I mc14500_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4329_ net141 _1263_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A1 _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4479__I _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__I _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__I3 _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3700_ _0650_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_138_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3973__A2 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ dffram.data\[30\]\[1\] _1527_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3631_ _2955_ _2962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6350_ _0307_ clknet_leaf_80_wb_clk_i dffram.data\[18\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4922__A1 _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3562_ dffram.data\[29\]\[4\] _2916_ _2917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5301_ _1935_ _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ _0238_ clknet_leaf_70_wb_clk_i dffram.data\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3493_ _1464_ _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3489__A1 _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _1894_ _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5163_ dffram.data\[51\]\[6\] _1852_ _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4114_ dffram.data\[62\]\[4\] dffram.data\[63\]\[4\] _1001_ _1059_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5094_ _1447_ _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4289__I0 dffram.data\[54\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4045_ _0708_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3661__A1 _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5996_ _2417_ _2418_ _2419_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3468__I _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4947_ _1693_ _1708_ _1711_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3413__A1 _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4878_ _1663_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3829_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5166__A1 _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ _0574_ clknet_leaf_4_wb_clk_i dffram.data\[32\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6548_ _0505_ clknet_leaf_157_wb_clk_i wb_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6479_ _0436_ clknet_leaf_122_wb_clk_i net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput271 net271 custom_settings[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput260 net260 custom_settings[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_144_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput293 net293 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput282 net282 custom_settings[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_96_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold53_I wbs_adr_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__I _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__I _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ dffram.data\[38\]\[4\] _2311_ _2312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5781_ _2256_ _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4199__A2 _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4801_ _1431_ _1524_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2993_ net249 _2462_ _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4732_ _1565_ _1555_ _1566_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4663_ _1510_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6402_ _0359_ clknet_leaf_76_wb_clk_i dffram.data\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3614_ dffram.data\[19\]\[5\] _2950_ _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4594_ _1464_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6333_ _0290_ clknet_leaf_91_wb_clk_i dffram.data\[45\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3545_ dffram.data\[32\]\[6\] _2903_ _2906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3476_ dffram.data\[35\]\[7\] _2856_ _2860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6264_ _0221_ clknet_leaf_107_wb_clk_i dffram.data\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5320__A1 dffram.data\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4123__A2 _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5215_ dffram.data\[50\]\[6\] _1886_ _1891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6195_ _0152_ clknet_leaf_168_wb_clk_i dffram.data\[25\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5146_ _1830_ _1583_ _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input147_I qcpu_sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _1788_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4277__I3 _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ dffram.data\[20\]\[3\] dffram.data\[21\]\[3\] _0843_ _0974_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3634__A1 _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4582__I _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ net228 _2404_ _2407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__A2 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A1 _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output366_I net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3873__A1 _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__I _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4492__I _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3836__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ net227 _2750_ _2751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3261_ _2483_ _2691_ _2694_ _2466_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5000_ _1741_ _1743_ _1745_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3192_ _2619_ wb_counter\[22\] _2637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5902_ dffram.data\[62\]\[5\] _2345_ _2347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_81_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5833_ dffram.data\[13\]\[6\] _2298_ _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5369__A1 _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3947__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5764_ _2214_ _2249_ _2254_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5695_ _2210_ _2207_ _2211_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4715_ _1463_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4646_ _1503_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5541__A1 _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_112_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4577_ _1441_ _1449_ _1450_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _0273_ clknet_leaf_101_wb_clk_i dffram.data\[46\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3528_ _2847_ _2019_ _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3459_ _2848_ _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3481__I _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _0204_ clknet_leaf_165_wb_clk_i dffram.data\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6178_ _0135_ clknet_leaf_116_wb_clk_i dffram.data\[53\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5129_ _1802_ _1832_ _1834_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3607__A1 _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3083__A2 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_67_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5532__A1 dffram.data\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold70 wbs_dat_i[16] net488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold81 wbs_dat_i[8] net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold92 wbs_dat_i[24] net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ dffram.data\[45\]\[0\] _2065_ _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4500_ net190 _1381_ _1375_ net41 _1376_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_26_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5523__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _1252_ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5781__I _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4362_ _1282_ _1286_ net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6101_ _0058_ clknet_leaf_33_wb_clk_i dffram.data\[63\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4293_ dffram.data\[34\]\[7\] dffram.data\[35\]\[7\] _1189_ _1235_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3313_ _2723_ _2724_ _2719_ _2736_ _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_74_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ net243 _2437_ _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3244_ _2663_ wb_counter\[30\] _2681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3175_ net381 _2609_ _2602_ _2622_ _2623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5816_ _2276_ _2062_ _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5747_ dffram.data\[12\]\[0\] _2244_ _2245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5762__A1 _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4565__A2 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_144_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input75_I mc14500_sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _2194_ _2197_ _2199_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4629_ dffram.data\[31\]\[1\] _1492_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__S _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output329_I net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_114_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3851__I1 dffram.data\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__I _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4010__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__I _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput160 qcpu_sram_in[7] net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput171 sid_do[19] net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput182 sid_oeb net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput193 sn76489_do[19] net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4244__A1 _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _1683_ _1729_ _1732_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ dffram.data\[52\]\[1\] dffram.data\[53\]\[1\] _0878_ _0879_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6650_ _0607_ clknet_leaf_45_wb_clk_i dffram.data\[61\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3862_ _0781_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_117_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6581_ _0538_ clknet_leaf_35_wb_clk_i dffram.data\[36\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5601_ _2148_ _2145_ _2149_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ dffram.data\[10\]\[7\] _2099_ _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3793_ _0739_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5463_ _2007_ _2048_ _2053_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4414_ _1321_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5394_ _2007_ _2000_ _2008_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4345_ net115 _1272_ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4276_ dffram.data\[14\]\[7\] dffram.data\[15\]\[7\] _1216_ _1218_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3227_ net390 _2654_ _2647_ _2666_ _2667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6015_ _2399_ _2433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3158_ _2601_ _2608_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4086__I1 dffram.data\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3089_ net215 _2352_ _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5983__A1 net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4538__A2 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output279_I net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4474__A1 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__B2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__I _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3824__I1 dffram.data\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5974__A1 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_82_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_11_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3737__B1 _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3844__I _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_39_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ dffram.data\[40\]\[4\] dffram.data\[41\]\[4\] _0772_ _1075_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3780__S _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4465__A1 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4061_ _0774_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4465__B2 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3012_ _2475_ _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_48_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _1714_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3914_ _0733_ _0861_ _0750_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_74_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _0590_ clknet_leaf_48_wb_clk_i dffram.data\[60\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4894_ dffram.data\[55\]\[5\] _1673_ _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ dffram.data\[32\]\[0\] dffram.data\[33\]\[0\] _0793_ _0794_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3955__S _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ _0699_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6564_ _0521_ clknet_leaf_146_wb_clk_i wb_counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5515_ _2091_ _2093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3754__I _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ _0452_ clknet_leaf_142_wb_clk_i net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5446_ _2009_ _2041_ _2043_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input177_I sid_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5377_ _1951_ _1992_ _1996_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4328_ _1262_ _1264_ net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4585__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input38_I mc14500_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4259_ dffram.data\[16\]\[7\] dffram.data\[17\]\[7\] _1200_ _1201_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5956__A1 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_137_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5708__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3865__S _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output396_I net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3990__I0 _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4695__A1 _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ _2930_ _2956_ _2961_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3561_ _2908_ _2916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _1935_ _1946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6280_ _0237_ clknet_leaf_70_wb_clk_i dffram.data\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3492_ _2870_ _2863_ _2871_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5231_ _1894_ _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5162_ _1822_ _1851_ _1854_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4113_ dffram.data\[60\]\[4\] dffram.data\[61\]\[4\] _0868_ _1058_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5093_ _1802_ _1804_ _1806_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4289__I1 dffram.data\[55\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4044_ dffram.data\[10\]\[3\] dffram.data\[11\]\[3\] _0923_ _0990_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_88_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_56_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5995_ _2395_ _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4946_ dffram.data\[28\]\[5\] _1709_ _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4877_ _1429_ _0789_ _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3828_ _0658_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6616_ _0573_ clknet_leaf_1_wb_clk_i dffram.data\[32\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_65_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6547_ _0504_ clknet_leaf_157_wb_clk_i wb_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3759_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3484__I _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3972__I0 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _0435_ clknet_leaf_122_wb_clk_i net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ dffram.data\[0\]\[7\] _2028_ _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput261 net261 custom_settings[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput272 net272 custom_settings[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput283 net283 custom_settings[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput294 net294 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_96_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6626__CLK clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output311_I net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5929__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4204__I1 _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3168__A1 _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3891__A2 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5093__A1 _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4953__I _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__A1 _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4800_ _1538_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5780_ _2076_ _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2992_ _2457_ _2462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ dffram.data\[2\]\[7\] _1556_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4662_ _1460_ _1511_ _1516_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6401_ _0358_ clknet_leaf_77_wb_clk_i dffram.data\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3613_ _2932_ _2949_ _2951_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4593_ _1463_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6332_ _0289_ clknet_leaf_91_wb_clk_i dffram.data\[45\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3544_ _2876_ _2902_ _2905_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3475_ _2333_ _2855_ _2859_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6263_ _0220_ clknet_leaf_127_wb_clk_i dffram.data\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5214_ _1824_ _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_0_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6194_ _0151_ clknet_leaf_168_wb_clk_i dffram.data\[25\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5145_ _1828_ _1838_ _1843_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5084__A1 _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _1750_ _1789_ _1794_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4027_ dffram.data\[18\]\[3\] dffram.data\[19\]\[3\] _0972_ _0973_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ net262 _2400_ _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _1433_ _1507_ _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_139_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_139_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__A1 dffram.data\[55\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output261_I net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5075__A1 dffram.data\[39\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4822__A1 _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4214__S _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A1 _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3852__I _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3260_ net223 _2693_ _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3191_ _2624_ _2636_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5066__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5901_ _2327_ _2344_ _2346_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ _2270_ _2297_ _2300_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5763_ dffram.data\[12\]\[7\] _2250_ _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _1551_ _1541_ _1552_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_134_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ dffram.data\[11\]\[5\] _2208_ _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _1484_ _1067_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_86_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4576_ dffram.data\[5\]\[1\] _1445_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6315_ _0272_ clknet_leaf_105_wb_clk_i dffram.data\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3527_ _2880_ _2889_ _2894_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4858__I _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3762__I _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3458_ _2848_ _2849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6246_ _0203_ clknet_leaf_164_wb_clk_i dffram.data\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _0134_ clknet_leaf_115_wb_clk_i dffram.data\[53\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3389_ _2792_ _2798_ _2799_ _2785_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_23_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input20_I ay8913_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3855__A2 _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ dffram.data\[52\]\[0\] _1833_ _1834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4593__I _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _1752_ _1782_ _1784_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_173_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3002__I _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_36_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5599__I _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold82 wbs_dat_i[22] net500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold71 wbs_dat_i[13] net489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4209__S _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold93 wbs_dat_i[7] net511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XPHY_EDGE_ROW_11_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4559__B1 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5220__A1 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3909__I0 dffram.data\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4430_ _1332_ _1334_ _1336_ net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_123_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_78_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3534__A1 _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4177__I3 _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3582__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6100_ _0057_ clknet_4_4_0_wb_clk_i dffram.data\[63\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4361_ net120 _1284_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ dffram.data\[32\]\[7\] dffram.data\[33\]\[7\] _1194_ _1234_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3312_ wb_counter\[9\] wb_counter\[10\] _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ net277 _2368_ _2445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3243_ _2668_ _2680_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4495__C1 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3174_ _2620_ _2621_ _2622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4119__S _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3958__S _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _2274_ _2284_ _2289_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5746_ _2242_ _2244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5677_ dffram.data\[11\]\[0\] _2198_ _2199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _1444_ _1491_ _1493_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input68_I mc14500_sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4588__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__A1 _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4559_ wb_sram_we _0717_ _0643_ net71 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_25_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6229_ _0186_ clknet_leaf_125_wb_clk_i dffram.data\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_154_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_154_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5450__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4005__A2 _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__A1 _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3819__A2 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput172 sid_do[1] net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput161 sid_do[0] net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput150 qcpu_sram_addr[4] net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput183 sn76489_do[0] net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput194 sn76489_do[1] net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_19_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__S _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3930_ _0778_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ dffram.data\[42\]\[0\] dffram.data\[43\]\[0\] _0809_ _0810_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3792_ dffram.data\[12\]\[0\] dffram.data\[13\]\[0\] _0740_ _0741_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5744__A2 _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5600_ dffram.data\[43\]\[5\] _2146_ _2149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6580_ _0537_ clknet_leaf_121_wb_clk_i wb_sram_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5531_ _2085_ _2098_ _2102_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3507__A1 _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5462_ dffram.data\[1\]\[3\] _2049_ _2053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4413_ _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5393_ dffram.data\[20\]\[3\] _2001_ _2008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4344_ _1271_ _1274_ net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4275_ dffram.data\[12\]\[7\] dffram.data\[13\]\[7\] _1216_ _1217_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4468__C1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6014_ _2431_ _2432_ _2430_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3226_ _2664_ _2665_ _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3157_ net378 _2587_ _2602_ _2607_ _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_38_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input122_I qcpu_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_120_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5432__A1 _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3088_ _2546_ _2547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_120_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3487__I _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_119_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5729_ _2200_ _2230_ _2233_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__A1 _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5207__I _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A1 _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3737__B2 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__A1 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold76_I wbs_dat_i[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__S _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3860__I _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4060_ dffram.data\[48\]\[3\] dffram.data\[49\]\[3\] _0875_ _1006_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3011_ _0752_ _0821_ _2477_ _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5414__A1 _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _1687_ _1715_ _1720_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3913_ _0857_ _0858_ _0859_ _0860_ _0744_ _0746_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_4893_ _1621_ _1672_ _1674_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6632_ _0589_ clknet_leaf_46_wb_clk_i dffram.data\[60\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3844_ _0753_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3775_ _0700_ _0716_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _0520_ clknet_leaf_147_wb_clk_i wb_counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5514_ _2091_ _2092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _0451_ clknet_leaf_142_wb_clk_i net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5445_ dffram.data\[46\]\[4\] _2042_ _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5376_ dffram.data\[47\]\[6\] _1993_ _1996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4327_ net140 _1263_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4258_ _0826_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3209_ _2648_ _2651_ _2652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4189_ _1129_ _1130_ _1131_ _1132_ _0785_ _0787_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5956__A2 _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3010__I _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output291_I net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5644__A1 _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5400__I _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4016__I _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3560_ _2908_ _2915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3491_ dffram.data\[34\]\[3\] _2864_ _2871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5230_ _1882_ _1895_ _1900_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3590__I _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5161_ dffram.data\[51\]\[5\] _1852_ _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4686__I _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4112_ dffram.data\[58\]\[4\] dffram.data\[59\]\[4\] _0998_ _1057_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5092_ dffram.data\[24\]\[0\] _1805_ _1806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4043_ dffram.data\[8\]\[3\] dffram.data\[9\]\[3\] _0734_ _0989_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5994_ net232 _2415_ _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4945_ _1689_ _1708_ _1710_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _1629_ _1657_ _1662_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6615_ _0572_ clknet_leaf_1_wb_clk_i dffram.data\[32\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3827_ dffram.data\[50\]\[0\] dffram.data\[51\]\[0\] _0775_ _0776_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3758_ _0659_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6546_ _0503_ clknet_leaf_157_wb_clk_i wb_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3689_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3972__I1 _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _0434_ clknet_leaf_120_wb_clk_i net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input50_I mc14500_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _2015_ _2027_ _2031_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput262 net262 custom_settings[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5359_ _1984_ _1859_ _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput273 net273 custom_settings[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput295 net295 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput284 net284 custom_settings[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5626__A1 _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3101__A2 _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output304_I net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3675__I _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2991_ _0632_ _2458_ _2461_ _2454_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ _1564_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3585__I _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4661_ dffram.data\[58\]\[3\] _1512_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6400_ _0357_ clknet_leaf_76_wb_clk_i dffram.data\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3612_ dffram.data\[19\]\[4\] _2950_ _2951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ net249 _1451_ _1457_ net157 _1452_ net76 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_114_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _0288_ clknet_leaf_107_wb_clk_i dffram.data\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3543_ dffram.data\[32\]\[5\] _2903_ _2905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3474_ dffram.data\[35\]\[6\] _2856_ _2859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6100__CLK clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6262_ _0219_ clknet_leaf_127_wb_clk_i dffram.data\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5213_ _1888_ _1885_ _1889_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6193_ _0150_ clknet_leaf_167_wb_clk_i dffram.data\[25\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5144_ dffram.data\[52\]\[7\] _1839_ _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5608__A1 _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ dffram.data\[39\]\[3\] _1790_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4026_ _0702_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_163_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input202_I sn76489_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5977_ _2403_ _2405_ _2396_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ _1697_ _1690_ _1698_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3495__I _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input98_I qcpu_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4859_ dffram.data\[56\]\[0\] _1652_ _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_108_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6529_ _0486_ clknet_leaf_141_wb_clk_i net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3086__A1 _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6024__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4586__B2 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4189__I1 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3936__I1 _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_84_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3190_ net384 _2632_ _2625_ _2635_ _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4964__I _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__A2 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5900_ dffram.data\[62\]\[4\] _2345_ _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_93_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ dffram.data\[13\]\[5\] _2298_ _2300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5762_ _2212_ _2249_ _2253_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_17_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4713_ dffram.data\[2\]\[3\] _1542_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5693_ _2081_ _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _1478_ _1497_ _1502_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4575_ _1448_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6314_ _0271_ clknet_leaf_104_wb_clk_i dffram.data\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3526_ dffram.data\[33\]\[7\] _2890_ _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4140__S _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _0202_ clknet_leaf_166_wb_clk_i dffram.data\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3457_ _2847_ _2195_ _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input152_I qcpu_sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _0133_ clknet_leaf_165_wb_clk_i dffram.data\[53\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3388_ net238 _2790_ _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_127_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5127_ _1831_ _1833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_127_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5058_ dffram.data\[25\]\[4\] _1783_ _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input13_I ay8913_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4009_ dffram.data\[44\]\[2\] dffram.data\[45\]\[2\] _0811_ _0956_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_140_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6006__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3240__A1 net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3953__I _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output371_I net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold50 wbs_cyc_i net468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold72 wbs_dat_i[14] net490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold94 wbs_dat_i[9] net512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4559__A1 wb_sram_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4559__B2 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__S _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__A2 _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4360_ _1282_ _1285_ net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3311_ wb_counter\[9\] _2727_ wb_counter\[10\] _2735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4291_ _1199_ _1232_ _0789_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_91_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _2443_ _2444_ _2442_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3242_ net392 _2491_ _2669_ _2679_ _2680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input5_I ay8913_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3173_ net267 _2604_ _2605_ _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3103__I _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5814_ dffram.data\[15\]\[7\] _2285_ _2289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5745_ _2242_ _2243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4270__I0 _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5676_ _2196_ _2198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4627_ dffram.data\[31\]\[0\] _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4558_ _1432_ _1089_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4489_ net165 _1383_ _1378_ net84 net5 _1379_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_3509_ _2882_ _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _0185_ clknet_leaf_125_wb_clk_i dffram.data\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3289__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _0116_ clknet_leaf_173_wb_clk_i dffram.data\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4789__A1 _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3461__A1 _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_123_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__S _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput140 qcpu_oeb[4] net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput162 sid_do[10] net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput151 qcpu_sram_addr[5] net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput173 sid_do[20] net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput195 sn76489_do[20] net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput184 sn76489_do[10] net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_19_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3858__I _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _0774_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3794__S _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3791_ _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ dffram.data\[10\]\[6\] _2099_ _2102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5461_ _2005_ _2048_ _2052_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3593__I _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4412_ _0623_ _0620_ _1278_ _1252_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_93_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3507__A2 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _1813_ _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4343_ net114 _1272_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4274_ _0826_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4468__B1 _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ net238 _2426_ _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3225_ net276 _2649_ _2650_ _2665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3156_ _2603_ _2606_ _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3818__I0 _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3087_ _2362_ _2546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_120_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5432__A2 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input115_I qcpu_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3443__A1 _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5196__A1 _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ dffram.data\[40\]\[1\] _2231_ _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3989_ dffram.data\[62\]\[2\] dffram.data\[63\]\[2\] _0762_ _0936_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input80_I qcpu_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5659_ _2140_ _2182_ _2186_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output334_I net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3678__I design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4234__I0 dffram.data\[38\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3737__A2 _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold69_I wbs_dat_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_91_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_107_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_71_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5111__A1 _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _2476_ _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3789__S _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3425__A1 _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4961_ dffram.data\[27\]\[3\] _1716_ _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3912_ dffram.data\[14\]\[1\] dffram.data\[15\]\[1\] _0742_ _0860_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ dffram.data\[55\]\[4\] _1673_ _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6631_ _0588_ clknet_leaf_45_wb_clk_i dffram.data\[60\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3843_ _0699_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5178__A1 _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3728__A2 design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__A1 _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3774_ _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6562_ _0519_ clknet_leaf_153_wb_clk_i wb_counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5513_ _1956_ _2090_ _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _0450_ clknet_4_10_0_wb_clk_i net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5444_ _2034_ _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput400 net400 wbs_dat_o[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_113_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__A2 _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__A1 _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _1949_ _1992_ _1995_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4326_ _1257_ _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4257_ _0698_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4188_ dffram.data\[46\]\[5\] dffram.data\[47\]\[5\] _0957_ _1132_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3208_ net273 _2649_ _2650_ _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3139_ _2572_ wb_counter\[14\] _2592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3498__I _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3416__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__A2 _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4392__A2 _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output284_I net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3990__I2 _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4278__B _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3742__I2 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3655__A1 _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__I _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A1 _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A2 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ _1459_ _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _1817_ _1851_ _1853_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4111_ dffram.data\[56\]\[4\] dffram.data\[57\]\[4\] _0865_ _1056_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5091_ _1803_ _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4042_ _0725_ _0987_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_153_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__A1 _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ net266 _2411_ _2417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4944_ dffram.data\[28\]\[4\] _1709_ _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4875_ dffram.data\[56\]\[7\] _1658_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3826_ _0774_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6614_ _0571_ clknet_leaf_1_wb_clk_i dffram.data\[32\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4143__S _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__A1 _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3757_ dffram.data\[18\]\[0\] dffram.data\[19\]\[0\] _0705_ _0706_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_104_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _0502_ clknet_leaf_134_wb_clk_i net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input182_I sid_oeb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3688_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _0433_ clknet_leaf_122_wb_clk_i net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_113_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5323__A1 _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ dffram.data\[0\]\[6\] _2028_ _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input43_I mc14500_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5358_ _1983_ _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput274 net274 custom_settings[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput263 net263 custom_settings[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_7_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput285 net285 custom_settings[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4309_ _1249_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput296 net296 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5289_ _1934_ _1936_ _1938_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_113_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5501__I _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6522__CLK clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_122_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_131_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3628__A1 _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__I _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4228__S _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2990_ net248 _2459_ _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_140_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3866__I _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4660_ _1455_ _1511_ _1515_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5553__A1 _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3611_ _2942_ _2950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4591_ _1440_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6330_ _0287_ clknet_leaf_105_wb_clk_i dffram.data\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3542_ _2872_ _2902_ _2904_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3473_ _2331_ _2855_ _2858_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4697__I _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _0218_ clknet_leaf_127_wb_clk_i dffram.data\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ dffram.data\[50\]\[5\] _1886_ _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6192_ _0149_ clknet_leaf_166_wb_clk_i dffram.data\[25\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _1825_ _1838_ _1842_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A2 _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3619__A1 _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _1748_ _1789_ _1793_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4025_ dffram.data\[16\]\[3\] dffram.data\[17\]\[3\] _0840_ _0971_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3095__A2 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3977__S _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A2 _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5976_ net227 _2404_ _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5792__A1 dffram.data\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ dffram.data\[54\]\[7\] _1691_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4858_ _1650_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ dffram.data\[58\]\[0\] dffram.data\[59\]\[0\] _0757_ _0758_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4789_ _1551_ _1598_ _1603_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6528_ _0485_ clknet_leaf_141_wb_clk_i net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _0416_ clknet_leaf_60_wb_clk_i dffram.data\[38\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_148_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_148_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_50_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4189__I2 _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6011__B _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3077__A2 _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _2266_ _2297_ _2299_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5761_ dffram.data\[12\]\[6\] _2250_ _2253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3596__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4577__A2 _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4712_ _1550_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_44_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5692_ _2206_ _2207_ _2209_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4643_ dffram.data\[31\]\[7\] _1498_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4574_ net403 _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_112_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _0270_ clknet_leaf_104_wb_clk_i dffram.data\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3525_ _2878_ _2889_ _2893_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6244_ _0201_ clknet_leaf_164_wb_clk_i dffram.data\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3456_ _1567_ _2847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3387_ _2795_ _2797_ _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6175_ _0132_ clknet_leaf_162_wb_clk_i dffram.data\[53\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input145_I qcpu_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5126_ _1831_ _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_127_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5057_ _1775_ _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4008_ dffram.data\[42\]\[2\] dffram.data\[43\]\[2\] _0954_ _0955_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3068__A2 wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__I _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5959_ net254 _2391_ _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A1 _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output364_I net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 net507 net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 wbs_dat_i[3] net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold73 wbs_dat_i[15] net491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold51 _1483_ net469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold95 wbs_dat_i[1] net513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold84 net428 net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4559__A2 _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2990__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4040__I _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5136__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3310_ _2732_ _2733_ _2734_ _2718_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _1228_ _1229_ _1230_ _1231_ _0834_ _0882_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_10_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4495__A1 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__I _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3241_ _2677_ _2678_ _2679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4495__B2 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3172_ _2619_ wb_counter\[19\] _2620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _2272_ _2284_ _2288_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5744_ _1956_ _2118_ _2242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5675_ _2196_ _2197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _1490_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4557_ _0674_ net476 _0678_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_111_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4488_ _1330_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3508_ _2882_ _2883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _2316_ _2835_ _2837_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6227_ _0184_ clknet_leaf_118_wb_clk_i dffram.data\[51\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6158_ _0115_ clknet_leaf_174_wb_clk_i dffram.data\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5109_ _1803_ _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ _0046_ clknet_leaf_38_wb_clk_i dffram.data\[37\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5986__A1 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_163_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_163_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5910__A1 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4477__A1 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__B2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput130 qcpu_oeb[25] net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput141 qcpu_oeb[5] net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput163 sid_do[11] net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold14_I wbs_adr_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput152 qcpu_sram_gwe net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput174 sid_do[2] net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput196 sn76489_do[21] net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput185 sn76489_do[11] net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3204__I _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4088__S0 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ _0701_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3874__I _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__A2 _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5460_ dffram.data\[1\]\[2\] _2049_ _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4411_ net161 _1316_ _1317_ net80 net1 _1318_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_93_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5901__A1 _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2005_ _2000_ _2006_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4342_ _1271_ _1273_ net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_120_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4273_ dffram.data\[10\]\[7\] dffram.data\[11\]\[7\] _1209_ _1215_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4468__B2 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__A1 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6012_ net272 _2422_ _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3224_ _2663_ wb_counter\[27\] _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

