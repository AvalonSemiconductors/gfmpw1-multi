VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_pdp11
  CLASS BLOCK ;
  FOREIGN wrapped_pdp11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1700.000 BY 800.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 452.480 4.000 453.040 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 667.520 4.000 668.080 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 703.360 4.000 703.920 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.200 4.000 739.760 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 775.040 4.000 775.600 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.440 4.000 238.000 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.960 4.000 345.520 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END custom_settings[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 0.000 12.880 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 0.000 476.560 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 0.000 502.320 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 38.080 0.000 38.640 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 0.000 528.080 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 0.000 553.840 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 0.000 605.360 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 0.000 682.640 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 0.000 708.400 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 733.600 0.000 734.160 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 785.120 0.000 785.680 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 810.880 0.000 811.440 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 0.000 837.200 4.000 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 22.400 1700.000 22.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 257.600 1700.000 258.160 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 281.120 1700.000 281.680 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 304.640 1700.000 305.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 328.160 1700.000 328.720 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 351.680 1700.000 352.240 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 375.200 1700.000 375.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 398.720 1700.000 399.280 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 422.240 1700.000 422.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 445.760 1700.000 446.320 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 469.280 1700.000 469.840 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 45.920 1700.000 46.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 492.800 1700.000 493.360 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 516.320 1700.000 516.880 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 539.840 1700.000 540.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 563.360 1700.000 563.920 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 586.880 1700.000 587.440 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 610.400 1700.000 610.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 633.920 1700.000 634.480 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 657.440 1700.000 658.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 680.960 1700.000 681.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 704.480 1700.000 705.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 69.440 1700.000 70.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 728.000 1700.000 728.560 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 751.520 1700.000 752.080 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 775.040 1700.000 775.600 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 92.960 1700.000 93.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 116.480 1700.000 117.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 140.000 1700.000 140.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 163.520 1700.000 164.080 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 187.040 1700.000 187.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 210.560 1700.000 211.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 1696.000 234.080 1700.000 234.640 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1120.000 0.000 1120.560 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 0.000 1146.320 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1171.520 0.000 1172.080 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1197.280 0.000 1197.840 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1223.040 0.000 1223.600 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1248.800 0.000 1249.360 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 1274.560 0.000 1275.120 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 0.000 1300.880 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1326.080 0.000 1326.640 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 1351.840 0.000 1352.400 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 888.160 0.000 888.720 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1377.600 0.000 1378.160 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1403.360 0.000 1403.920 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1429.120 0.000 1429.680 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 1454.880 0.000 1455.440 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1480.640 0.000 1481.200 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 1506.400 0.000 1506.960 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1532.160 0.000 1532.720 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1557.920 0.000 1558.480 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1583.680 0.000 1584.240 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 0.000 1610.000 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 0.000 914.480 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1635.200 0.000 1635.760 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1660.960 0.000 1661.520 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1686.720 0.000 1687.280 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 0.000 940.240 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 0.000 966.000 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1016.960 0.000 1017.520 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 0.000 1043.280 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 0.000 1069.040 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1094.240 0.000 1094.800 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 4.000 58.800 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 4.000 22.960 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 15.250 1693.310 784.430 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1692.880 784.300 ;
      LAYER Metal2 ;
        RECT 0.140 4.300 1691.340 784.190 ;
        RECT 0.140 3.450 12.020 4.300 ;
        RECT 13.180 3.450 37.780 4.300 ;
        RECT 38.940 3.450 63.540 4.300 ;
        RECT 64.700 3.450 89.300 4.300 ;
        RECT 90.460 3.450 115.060 4.300 ;
        RECT 116.220 3.450 140.820 4.300 ;
        RECT 141.980 3.450 166.580 4.300 ;
        RECT 167.740 3.450 192.340 4.300 ;
        RECT 193.500 3.450 218.100 4.300 ;
        RECT 219.260 3.450 243.860 4.300 ;
        RECT 245.020 3.450 269.620 4.300 ;
        RECT 270.780 3.450 295.380 4.300 ;
        RECT 296.540 3.450 321.140 4.300 ;
        RECT 322.300 3.450 346.900 4.300 ;
        RECT 348.060 3.450 372.660 4.300 ;
        RECT 373.820 3.450 398.420 4.300 ;
        RECT 399.580 3.450 424.180 4.300 ;
        RECT 425.340 3.450 449.940 4.300 ;
        RECT 451.100 3.450 475.700 4.300 ;
        RECT 476.860 3.450 501.460 4.300 ;
        RECT 502.620 3.450 527.220 4.300 ;
        RECT 528.380 3.450 552.980 4.300 ;
        RECT 554.140 3.450 578.740 4.300 ;
        RECT 579.900 3.450 604.500 4.300 ;
        RECT 605.660 3.450 630.260 4.300 ;
        RECT 631.420 3.450 656.020 4.300 ;
        RECT 657.180 3.450 681.780 4.300 ;
        RECT 682.940 3.450 707.540 4.300 ;
        RECT 708.700 3.450 733.300 4.300 ;
        RECT 734.460 3.450 759.060 4.300 ;
        RECT 760.220 3.450 784.820 4.300 ;
        RECT 785.980 3.450 810.580 4.300 ;
        RECT 811.740 3.450 836.340 4.300 ;
        RECT 837.500 3.450 862.100 4.300 ;
        RECT 863.260 3.450 887.860 4.300 ;
        RECT 889.020 3.450 913.620 4.300 ;
        RECT 914.780 3.450 939.380 4.300 ;
        RECT 940.540 3.450 965.140 4.300 ;
        RECT 966.300 3.450 990.900 4.300 ;
        RECT 992.060 3.450 1016.660 4.300 ;
        RECT 1017.820 3.450 1042.420 4.300 ;
        RECT 1043.580 3.450 1068.180 4.300 ;
        RECT 1069.340 3.450 1093.940 4.300 ;
        RECT 1095.100 3.450 1119.700 4.300 ;
        RECT 1120.860 3.450 1145.460 4.300 ;
        RECT 1146.620 3.450 1171.220 4.300 ;
        RECT 1172.380 3.450 1196.980 4.300 ;
        RECT 1198.140 3.450 1222.740 4.300 ;
        RECT 1223.900 3.450 1248.500 4.300 ;
        RECT 1249.660 3.450 1274.260 4.300 ;
        RECT 1275.420 3.450 1300.020 4.300 ;
        RECT 1301.180 3.450 1325.780 4.300 ;
        RECT 1326.940 3.450 1351.540 4.300 ;
        RECT 1352.700 3.450 1377.300 4.300 ;
        RECT 1378.460 3.450 1403.060 4.300 ;
        RECT 1404.220 3.450 1428.820 4.300 ;
        RECT 1429.980 3.450 1454.580 4.300 ;
        RECT 1455.740 3.450 1480.340 4.300 ;
        RECT 1481.500 3.450 1506.100 4.300 ;
        RECT 1507.260 3.450 1531.860 4.300 ;
        RECT 1533.020 3.450 1557.620 4.300 ;
        RECT 1558.780 3.450 1583.380 4.300 ;
        RECT 1584.540 3.450 1609.140 4.300 ;
        RECT 1610.300 3.450 1634.900 4.300 ;
        RECT 1636.060 3.450 1660.660 4.300 ;
        RECT 1661.820 3.450 1686.420 4.300 ;
        RECT 1687.580 3.450 1691.340 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 775.900 1696.000 784.140 ;
        RECT 4.300 774.740 1695.700 775.900 ;
        RECT 0.090 752.380 1696.000 774.740 ;
        RECT 0.090 751.220 1695.700 752.380 ;
        RECT 0.090 740.060 1696.000 751.220 ;
        RECT 4.300 738.900 1696.000 740.060 ;
        RECT 0.090 728.860 1696.000 738.900 ;
        RECT 0.090 727.700 1695.700 728.860 ;
        RECT 0.090 705.340 1696.000 727.700 ;
        RECT 0.090 704.220 1695.700 705.340 ;
        RECT 4.300 704.180 1695.700 704.220 ;
        RECT 4.300 703.060 1696.000 704.180 ;
        RECT 0.090 681.820 1696.000 703.060 ;
        RECT 0.090 680.660 1695.700 681.820 ;
        RECT 0.090 668.380 1696.000 680.660 ;
        RECT 4.300 667.220 1696.000 668.380 ;
        RECT 0.090 658.300 1696.000 667.220 ;
        RECT 0.090 657.140 1695.700 658.300 ;
        RECT 0.090 634.780 1696.000 657.140 ;
        RECT 0.090 633.620 1695.700 634.780 ;
        RECT 0.090 632.540 1696.000 633.620 ;
        RECT 4.300 631.380 1696.000 632.540 ;
        RECT 0.090 611.260 1696.000 631.380 ;
        RECT 0.090 610.100 1695.700 611.260 ;
        RECT 0.090 596.700 1696.000 610.100 ;
        RECT 4.300 595.540 1696.000 596.700 ;
        RECT 0.090 587.740 1696.000 595.540 ;
        RECT 0.090 586.580 1695.700 587.740 ;
        RECT 0.090 564.220 1696.000 586.580 ;
        RECT 0.090 563.060 1695.700 564.220 ;
        RECT 0.090 560.860 1696.000 563.060 ;
        RECT 4.300 559.700 1696.000 560.860 ;
        RECT 0.090 540.700 1696.000 559.700 ;
        RECT 0.090 539.540 1695.700 540.700 ;
        RECT 0.090 525.020 1696.000 539.540 ;
        RECT 4.300 523.860 1696.000 525.020 ;
        RECT 0.090 517.180 1696.000 523.860 ;
        RECT 0.090 516.020 1695.700 517.180 ;
        RECT 0.090 493.660 1696.000 516.020 ;
        RECT 0.090 492.500 1695.700 493.660 ;
        RECT 0.090 489.180 1696.000 492.500 ;
        RECT 4.300 488.020 1696.000 489.180 ;
        RECT 0.090 470.140 1696.000 488.020 ;
        RECT 0.090 468.980 1695.700 470.140 ;
        RECT 0.090 453.340 1696.000 468.980 ;
        RECT 4.300 452.180 1696.000 453.340 ;
        RECT 0.090 446.620 1696.000 452.180 ;
        RECT 0.090 445.460 1695.700 446.620 ;
        RECT 0.090 423.100 1696.000 445.460 ;
        RECT 0.090 421.940 1695.700 423.100 ;
        RECT 0.090 417.500 1696.000 421.940 ;
        RECT 4.300 416.340 1696.000 417.500 ;
        RECT 0.090 399.580 1696.000 416.340 ;
        RECT 0.090 398.420 1695.700 399.580 ;
        RECT 0.090 381.660 1696.000 398.420 ;
        RECT 4.300 380.500 1696.000 381.660 ;
        RECT 0.090 376.060 1696.000 380.500 ;
        RECT 0.090 374.900 1695.700 376.060 ;
        RECT 0.090 352.540 1696.000 374.900 ;
        RECT 0.090 351.380 1695.700 352.540 ;
        RECT 0.090 345.820 1696.000 351.380 ;
        RECT 4.300 344.660 1696.000 345.820 ;
        RECT 0.090 329.020 1696.000 344.660 ;
        RECT 0.090 327.860 1695.700 329.020 ;
        RECT 0.090 309.980 1696.000 327.860 ;
        RECT 4.300 308.820 1696.000 309.980 ;
        RECT 0.090 305.500 1696.000 308.820 ;
        RECT 0.090 304.340 1695.700 305.500 ;
        RECT 0.090 281.980 1696.000 304.340 ;
        RECT 0.090 280.820 1695.700 281.980 ;
        RECT 0.090 274.140 1696.000 280.820 ;
        RECT 4.300 272.980 1696.000 274.140 ;
        RECT 0.090 258.460 1696.000 272.980 ;
        RECT 0.090 257.300 1695.700 258.460 ;
        RECT 0.090 238.300 1696.000 257.300 ;
        RECT 4.300 237.140 1696.000 238.300 ;
        RECT 0.090 234.940 1696.000 237.140 ;
        RECT 0.090 233.780 1695.700 234.940 ;
        RECT 0.090 211.420 1696.000 233.780 ;
        RECT 0.090 210.260 1695.700 211.420 ;
        RECT 0.090 202.460 1696.000 210.260 ;
        RECT 4.300 201.300 1696.000 202.460 ;
        RECT 0.090 187.900 1696.000 201.300 ;
        RECT 0.090 186.740 1695.700 187.900 ;
        RECT 0.090 166.620 1696.000 186.740 ;
        RECT 4.300 165.460 1696.000 166.620 ;
        RECT 0.090 164.380 1696.000 165.460 ;
        RECT 0.090 163.220 1695.700 164.380 ;
        RECT 0.090 140.860 1696.000 163.220 ;
        RECT 0.090 139.700 1695.700 140.860 ;
        RECT 0.090 130.780 1696.000 139.700 ;
        RECT 4.300 129.620 1696.000 130.780 ;
        RECT 0.090 117.340 1696.000 129.620 ;
        RECT 0.090 116.180 1695.700 117.340 ;
        RECT 0.090 94.940 1696.000 116.180 ;
        RECT 4.300 93.820 1696.000 94.940 ;
        RECT 4.300 93.780 1695.700 93.820 ;
        RECT 0.090 92.660 1695.700 93.780 ;
        RECT 0.090 70.300 1696.000 92.660 ;
        RECT 0.090 69.140 1695.700 70.300 ;
        RECT 0.090 59.100 1696.000 69.140 ;
        RECT 4.300 57.940 1696.000 59.100 ;
        RECT 0.090 46.780 1696.000 57.940 ;
        RECT 0.090 45.620 1695.700 46.780 ;
        RECT 0.090 23.260 1696.000 45.620 ;
        RECT 4.300 22.100 1695.700 23.260 ;
        RECT 0.090 3.500 1696.000 22.100 ;
      LAYER Metal4 ;
        RECT 68.460 15.080 98.740 782.230 ;
        RECT 100.940 15.080 175.540 782.230 ;
        RECT 177.740 15.080 252.340 782.230 ;
        RECT 254.540 15.080 329.140 782.230 ;
        RECT 331.340 15.080 405.940 782.230 ;
        RECT 408.140 15.080 482.740 782.230 ;
        RECT 484.940 15.080 559.540 782.230 ;
        RECT 561.740 15.080 636.340 782.230 ;
        RECT 638.540 15.080 713.140 782.230 ;
        RECT 715.340 15.080 789.940 782.230 ;
        RECT 792.140 15.080 866.740 782.230 ;
        RECT 868.940 15.080 943.540 782.230 ;
        RECT 945.740 15.080 1020.340 782.230 ;
        RECT 1022.540 15.080 1097.140 782.230 ;
        RECT 1099.340 15.080 1173.940 782.230 ;
        RECT 1176.140 15.080 1250.740 782.230 ;
        RECT 1252.940 15.080 1327.540 782.230 ;
        RECT 1329.740 15.080 1404.340 782.230 ;
        RECT 1406.540 15.080 1441.860 782.230 ;
        RECT 68.460 6.250 1441.860 15.080 ;
  END
END wrapped_pdp11
END LIBRARY

