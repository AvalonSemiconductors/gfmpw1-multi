magic
tech gf180mcuD
magscale 1 10
timestamp 1698874740
<< nwell >>
rect 1258 31712 34694 32230
rect 1258 30144 34694 31008
rect 1258 28601 34694 29440
rect 1258 28576 9149 28601
rect 1258 27847 11053 27872
rect 1258 27033 34694 27847
rect 1258 27008 2541 27033
rect 1258 26279 2541 26304
rect 1258 25465 34694 26279
rect 1258 25440 7805 25465
rect 1258 24711 20716 24736
rect 1258 23897 34694 24711
rect 1258 23872 7917 23897
rect 1258 23143 2877 23168
rect 1258 22329 34694 23143
rect 1258 22304 2541 22329
rect 1258 21575 28456 21600
rect 1258 20761 34694 21575
rect 1258 20736 23821 20761
rect 1258 20007 2653 20032
rect 1258 19193 34694 20007
rect 1258 19168 2541 19193
rect 1258 18439 14749 18464
rect 1258 17625 34694 18439
rect 1258 17600 2541 17625
rect 1258 16871 3997 16896
rect 1258 16057 34694 16871
rect 1258 16032 2989 16057
rect 1258 15303 6461 15328
rect 1258 14489 34694 15303
rect 1258 14464 2541 14489
rect 1258 13735 29688 13760
rect 1258 12921 34694 13735
rect 1258 12896 8701 12921
rect 1258 12167 18221 12192
rect 1258 11353 34694 12167
rect 1258 11328 14301 11353
rect 1258 10599 13069 10624
rect 1258 9785 34694 10599
rect 1258 9760 32109 9785
rect 1258 9031 12952 9056
rect 1258 8217 34694 9031
rect 1258 8192 12311 8217
rect 1258 7463 19565 7488
rect 1258 6649 34694 7463
rect 1258 6624 16093 6649
rect 1258 5895 23718 5920
rect 1258 5081 34694 5895
rect 1258 5056 25992 5081
rect 1258 4327 2541 4352
rect 1258 3513 34694 4327
rect 1258 3488 10269 3513
<< pwell >>
rect 1258 31008 34694 31712
rect 1258 29440 34694 30144
rect 1258 27872 34694 28576
rect 1258 26304 34694 27008
rect 1258 24736 34694 25440
rect 1258 23168 34694 23872
rect 1258 21600 34694 22304
rect 1258 20032 34694 20736
rect 1258 18464 34694 19168
rect 1258 16896 34694 17600
rect 1258 15328 34694 16032
rect 1258 13760 34694 14464
rect 1258 12192 34694 12896
rect 1258 10624 34694 11328
rect 1258 9056 34694 9760
rect 1258 7488 34694 8192
rect 1258 5920 34694 6624
rect 1258 4352 34694 5056
rect 1258 3050 34694 3488
<< obsm1 >>
rect 1344 3076 34768 32204
<< metal2 >>
rect 3584 0 3696 800
rect 10752 0 10864 800
rect 17920 0 18032 800
rect 25088 0 25200 800
rect 32256 0 32368 800
<< obsm2 >>
rect 1596 860 34740 32182
rect 1596 800 3524 860
rect 3756 800 10692 860
rect 10924 800 17860 860
rect 18092 800 25028 860
rect 25260 800 32196 860
rect 32428 800 34740 860
<< obsm3 >>
rect 1586 3108 34750 32172
<< metal4 >>
rect 5342 3076 5662 32204
rect 9500 3076 9820 32204
rect 13658 3076 13978 32204
rect 17816 3076 18136 32204
rect 21974 3076 22294 32204
rect 26132 3076 26452 32204
rect 30290 3076 30610 32204
rect 34448 3076 34768 32204
<< obsm4 >>
rect 4620 4498 5282 25294
rect 5722 4498 9440 25294
rect 9880 4498 13598 25294
rect 14038 4498 17756 25294
rect 18196 4498 21914 25294
rect 22354 4498 26072 25294
rect 26512 4498 26852 25294
<< labels >>
rlabel metal2 s 17920 0 18032 800 6 io_out[0]
port 1 nsew signal output
rlabel metal2 s 25088 0 25200 800 6 io_out[1]
port 2 nsew signal output
rlabel metal2 s 32256 0 32368 800 6 io_out[2]
port 3 nsew signal output
rlabel metal2 s 10752 0 10864 800 6 rst_n
port 4 nsew signal input
rlabel metal4 s 5342 3076 5662 32204 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 13658 3076 13978 32204 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 21974 3076 22294 32204 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 30290 3076 30610 32204 6 vdd
port 5 nsew power bidirectional
rlabel metal4 s 9500 3076 9820 32204 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 17816 3076 18136 32204 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 26132 3076 26452 32204 6 vss
port 6 nsew ground bidirectional
rlabel metal4 s 34448 3076 34768 32204 6 vss
port 6 nsew ground bidirectional
rlabel metal2 s 3584 0 3696 800 6 wb_clk_i
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 36000 36000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1086608
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1_group/openlane/blinker/runs/23_11_01_22_36/results/signoff/blinker.magic.gds
string GDS_START 255932
<< end >>

