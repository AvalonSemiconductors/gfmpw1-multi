magic
tech gf180mcuD
magscale 1 5
timestamp 1753965955
<< nwell >>
rect 629 20561 22331 20991
rect 629 19777 22331 20207
rect 629 18993 22331 19423
rect 629 18209 22331 18639
rect 629 17425 22331 17855
rect 629 16641 22331 17071
rect 629 15857 22331 16287
rect 629 15073 22331 15503
rect 629 14289 22331 14719
rect 629 13505 22331 13935
rect 629 12721 22331 13151
rect 629 11937 22331 12367
rect 629 11153 22331 11583
rect 629 10369 22331 10799
rect 629 9585 22331 10015
rect 629 8801 22331 9231
rect 629 8017 22331 8447
rect 629 7233 22331 7663
rect 629 6449 22331 6879
rect 629 5665 22331 6095
rect 629 4881 22331 5311
rect 629 4097 22331 4527
rect 629 3313 22331 3743
rect 629 2529 22331 2959
rect 629 1745 22331 2175
<< pwell >>
rect 629 20991 22331 21211
rect 629 20207 22331 20561
rect 629 19423 22331 19777
rect 629 18639 22331 18993
rect 629 17855 22331 18209
rect 629 17071 22331 17425
rect 629 16287 22331 16641
rect 629 15503 22331 15857
rect 629 14719 22331 15073
rect 629 13935 22331 14289
rect 629 13151 22331 13505
rect 629 12367 22331 12721
rect 629 11583 22331 11937
rect 629 10799 22331 11153
rect 629 10015 22331 10369
rect 629 9231 22331 9585
rect 629 8447 22331 8801
rect 629 7663 22331 8017
rect 629 6879 22331 7233
rect 629 6095 22331 6449
rect 629 5311 22331 5665
rect 629 4527 22331 4881
rect 629 3743 22331 4097
rect 629 2959 22331 3313
rect 629 2175 22331 2529
rect 629 1525 22331 1745
<< obsm1 >>
rect 672 1538 22288 21198
<< metal2 >>
rect 896 22600 952 23000
rect 2800 22600 2856 23000
rect 4704 22600 4760 23000
rect 6608 22600 6664 23000
rect 8512 22600 8568 23000
rect 10416 22600 10472 23000
rect 12320 22600 12376 23000
rect 14224 22600 14280 23000
rect 16128 22600 16184 23000
rect 18032 22600 18088 23000
rect 19936 22600 19992 23000
rect 21840 22600 21896 23000
<< obsm2 >>
rect 854 22570 866 22600
rect 982 22570 2770 22600
rect 2886 22570 4674 22600
rect 4790 22570 6578 22600
rect 6694 22570 8482 22600
rect 8598 22570 10386 22600
rect 10502 22570 12290 22600
rect 12406 22570 14194 22600
rect 14310 22570 16098 22600
rect 16214 22570 18002 22600
rect 18118 22570 19906 22600
rect 20022 22570 21810 22600
rect 21926 22570 21938 22600
rect 854 1549 21938 22570
<< obsm3 >>
rect 849 1554 21943 21182
<< metal4 >>
rect 2224 1538 2384 21198
rect 9904 1538 10064 21198
rect 17584 1538 17744 21198
<< obsm4 >>
rect 7462 12273 9874 17183
rect 10094 12273 17554 17183
rect 17774 12273 19922 17183
<< labels >>
rlabel metal2 s 4704 22600 4760 23000 6 io_in
port 1 nsew signal input
rlabel metal2 s 6608 22600 6664 23000 6 io_out[0]
port 2 nsew signal output
rlabel metal2 s 8512 22600 8568 23000 6 io_out[1]
port 3 nsew signal output
rlabel metal2 s 10416 22600 10472 23000 6 io_out[2]
port 4 nsew signal output
rlabel metal2 s 12320 22600 12376 23000 6 io_out[3]
port 5 nsew signal output
rlabel metal2 s 14224 22600 14280 23000 6 io_out[4]
port 6 nsew signal output
rlabel metal2 s 16128 22600 16184 23000 6 io_out[5]
port 7 nsew signal output
rlabel metal2 s 18032 22600 18088 23000 6 io_out[6]
port 8 nsew signal output
rlabel metal2 s 19936 22600 19992 23000 6 io_out[7]
port 9 nsew signal output
rlabel metal2 s 21840 22600 21896 23000 6 io_out[8]
port 10 nsew signal output
rlabel metal2 s 2800 22600 2856 23000 6 rst_n
port 11 nsew signal input
rlabel metal4 s 2224 1538 2384 21198 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 21198 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 21198 6 vss
port 13 nsew ground bidirectional
rlabel metal2 s 896 22600 952 23000 6 wb_clk_i
port 14 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 980604
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/diceroll/runs/25_07_31_14_44/results/signoff/diceroll.magic.gds
string GDS_START 163264
<< end >>

