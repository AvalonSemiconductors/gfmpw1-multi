VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_sid
  CLASS BLOCK ;
  FOREIGN wrapped_sid ;
  ORIGIN 0.000 0.000 ;
  SIZE 1150.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 13.440 1150.000 14.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 159.040 1150.000 159.600 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 173.600 1150.000 174.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 188.160 1150.000 188.720 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 202.720 1150.000 203.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 217.280 1150.000 217.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 231.840 1150.000 232.400 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 246.400 1150.000 246.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 260.960 1150.000 261.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 275.520 1150.000 276.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 290.080 1150.000 290.640 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 28.000 1150.000 28.560 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 304.640 1150.000 305.200 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 319.200 1150.000 319.760 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 333.760 1150.000 334.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 348.320 1150.000 348.880 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 362.880 1150.000 363.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 377.440 1150.000 378.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 392.000 1150.000 392.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 406.560 1150.000 407.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 421.120 1150.000 421.680 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 435.680 1150.000 436.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 42.560 1150.000 43.120 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 450.240 1150.000 450.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 464.800 1150.000 465.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 479.360 1150.000 479.920 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 57.120 1150.000 57.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 71.680 1150.000 72.240 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 86.240 1150.000 86.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 100.800 1150.000 101.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 115.360 1150.000 115.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 129.920 1150.000 130.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 144.480 1150.000 145.040 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 796.000 575.120 800.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 493.920 1150.000 494.480 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 639.520 1150.000 640.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 654.080 1150.000 654.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 668.640 1150.000 669.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 683.200 1150.000 683.760 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 697.760 1150.000 698.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 712.320 1150.000 712.880 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 726.880 1150.000 727.440 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 741.440 1150.000 742.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 756.000 1150.000 756.560 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 770.560 1150.000 771.120 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 508.480 1150.000 509.040 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 785.120 1150.000 785.680 ;
    END
  END io_out[20]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 523.040 1150.000 523.600 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 537.600 1150.000 538.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 552.160 1150.000 552.720 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 566.720 1150.000 567.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 581.280 1150.000 581.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 595.840 1150.000 596.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 610.400 1150.000 610.960 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1146.000 624.960 1150.000 625.520 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 0.000 861.840 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 782.240 1143.390 784.430 ;
      LAYER Nwell ;
        RECT 6.290 782.115 203.990 782.240 ;
        RECT 6.290 778.045 1143.390 782.115 ;
        RECT 6.290 777.920 173.820 778.045 ;
      LAYER Pwell ;
        RECT 6.290 774.400 1143.390 777.920 ;
      LAYER Nwell ;
        RECT 6.290 774.275 179.780 774.400 ;
        RECT 6.290 770.205 1143.390 774.275 ;
        RECT 6.290 770.080 128.600 770.205 ;
      LAYER Pwell ;
        RECT 6.290 766.560 1143.390 770.080 ;
      LAYER Nwell ;
        RECT 6.290 766.435 141.085 766.560 ;
        RECT 6.290 762.365 1143.390 766.435 ;
        RECT 6.290 762.240 123.910 762.365 ;
      LAYER Pwell ;
        RECT 6.290 758.720 1143.390 762.240 ;
      LAYER Nwell ;
        RECT 6.290 758.595 118.315 758.720 ;
        RECT 6.290 754.525 1143.390 758.595 ;
        RECT 6.290 754.400 69.905 754.525 ;
      LAYER Pwell ;
        RECT 6.290 750.880 1143.390 754.400 ;
      LAYER Nwell ;
        RECT 6.290 750.755 79.390 750.880 ;
        RECT 6.290 746.685 1143.390 750.755 ;
        RECT 6.290 746.560 76.125 746.685 ;
      LAYER Pwell ;
        RECT 6.290 743.040 1143.390 746.560 ;
      LAYER Nwell ;
        RECT 6.290 742.915 65.320 743.040 ;
        RECT 6.290 738.845 1143.390 742.915 ;
        RECT 6.290 738.720 54.540 738.845 ;
      LAYER Pwell ;
        RECT 6.290 735.200 1143.390 738.720 ;
      LAYER Nwell ;
        RECT 6.290 735.075 52.510 735.200 ;
        RECT 6.290 731.005 1143.390 735.075 ;
        RECT 6.290 730.880 39.115 731.005 ;
      LAYER Pwell ;
        RECT 6.290 727.360 1143.390 730.880 ;
      LAYER Nwell ;
        RECT 6.290 727.235 29.480 727.360 ;
        RECT 6.290 723.165 1143.390 727.235 ;
        RECT 6.290 723.040 40.120 723.165 ;
      LAYER Pwell ;
        RECT 6.290 719.520 1143.390 723.040 ;
      LAYER Nwell ;
        RECT 6.290 719.395 23.995 719.520 ;
        RECT 6.290 715.325 1143.390 719.395 ;
        RECT 6.290 715.200 75.515 715.325 ;
      LAYER Pwell ;
        RECT 6.290 711.680 1143.390 715.200 ;
      LAYER Nwell ;
        RECT 6.290 711.555 74.350 711.680 ;
        RECT 6.290 707.485 1143.390 711.555 ;
        RECT 6.290 707.360 13.800 707.485 ;
      LAYER Pwell ;
        RECT 6.290 703.840 1143.390 707.360 ;
      LAYER Nwell ;
        RECT 6.290 703.715 20.700 703.840 ;
        RECT 6.290 699.645 1143.390 703.715 ;
        RECT 6.290 699.520 33.400 699.645 ;
      LAYER Pwell ;
        RECT 6.290 696.000 1143.390 699.520 ;
      LAYER Nwell ;
        RECT 6.290 695.875 15.900 696.000 ;
        RECT 6.290 691.805 1143.390 695.875 ;
        RECT 6.290 691.680 31.790 691.805 ;
      LAYER Pwell ;
        RECT 6.290 688.160 1143.390 691.680 ;
      LAYER Nwell ;
        RECT 6.290 688.035 12.185 688.160 ;
        RECT 6.290 683.965 1143.390 688.035 ;
        RECT 6.290 683.840 35.150 683.965 ;
      LAYER Pwell ;
        RECT 6.290 680.320 1143.390 683.840 ;
      LAYER Nwell ;
        RECT 6.290 680.195 78.550 680.320 ;
        RECT 6.290 676.125 1143.390 680.195 ;
        RECT 6.290 676.000 76.030 676.125 ;
      LAYER Pwell ;
        RECT 6.290 672.480 1143.390 676.000 ;
      LAYER Nwell ;
        RECT 6.290 672.355 37.390 672.480 ;
        RECT 6.290 668.285 1143.390 672.355 ;
        RECT 6.290 668.160 91.710 668.285 ;
      LAYER Pwell ;
        RECT 6.290 664.640 1143.390 668.160 ;
      LAYER Nwell ;
        RECT 6.290 664.515 21.195 664.640 ;
        RECT 6.290 660.445 1143.390 664.515 ;
        RECT 6.290 660.320 13.310 660.445 ;
      LAYER Pwell ;
        RECT 6.290 656.800 1143.390 660.320 ;
      LAYER Nwell ;
        RECT 6.290 656.675 15.585 656.800 ;
        RECT 6.290 652.605 1143.390 656.675 ;
        RECT 6.290 652.480 15.830 652.605 ;
      LAYER Pwell ;
        RECT 6.290 648.960 1143.390 652.480 ;
      LAYER Nwell ;
        RECT 6.290 648.835 132.075 648.960 ;
        RECT 6.290 644.765 1143.390 648.835 ;
        RECT 6.290 644.640 23.670 644.765 ;
      LAYER Pwell ;
        RECT 6.290 641.120 1143.390 644.640 ;
      LAYER Nwell ;
        RECT 6.290 640.995 9.435 641.120 ;
        RECT 6.290 636.925 1143.390 640.995 ;
        RECT 6.290 636.800 56.465 636.925 ;
      LAYER Pwell ;
        RECT 6.290 633.280 1143.390 636.800 ;
      LAYER Nwell ;
        RECT 6.290 633.155 9.390 633.280 ;
        RECT 6.290 629.085 1143.390 633.155 ;
        RECT 6.290 628.960 17.275 629.085 ;
      LAYER Pwell ;
        RECT 6.290 625.440 1143.390 628.960 ;
      LAYER Nwell ;
        RECT 6.290 625.315 209.915 625.440 ;
        RECT 6.290 621.245 1143.390 625.315 ;
        RECT 6.290 621.120 38.230 621.245 ;
      LAYER Pwell ;
        RECT 6.290 617.600 1143.390 621.120 ;
      LAYER Nwell ;
        RECT 6.290 617.475 14.465 617.600 ;
        RECT 6.290 613.405 1143.390 617.475 ;
        RECT 6.290 613.280 86.715 613.405 ;
      LAYER Pwell ;
        RECT 6.290 609.760 1143.390 613.280 ;
      LAYER Nwell ;
        RECT 6.290 609.635 23.110 609.760 ;
        RECT 6.290 605.565 1143.390 609.635 ;
        RECT 6.290 605.440 14.475 605.565 ;
      LAYER Pwell ;
        RECT 6.290 601.920 1143.390 605.440 ;
      LAYER Nwell ;
        RECT 6.290 601.795 20.590 601.920 ;
        RECT 6.290 597.725 1143.390 601.795 ;
        RECT 6.290 597.600 70.985 597.725 ;
      LAYER Pwell ;
        RECT 6.290 594.080 1143.390 597.600 ;
      LAYER Nwell ;
        RECT 6.290 593.955 137.070 594.080 ;
        RECT 6.290 589.885 1143.390 593.955 ;
        RECT 6.290 589.760 68.190 589.885 ;
      LAYER Pwell ;
        RECT 6.290 586.240 1143.390 589.760 ;
      LAYER Nwell ;
        RECT 6.290 586.115 32.910 586.240 ;
        RECT 6.290 582.045 1143.390 586.115 ;
        RECT 6.290 581.920 165.065 582.045 ;
      LAYER Pwell ;
        RECT 6.290 578.400 1143.390 581.920 ;
      LAYER Nwell ;
        RECT 6.290 578.275 68.750 578.400 ;
        RECT 6.290 574.205 1143.390 578.275 ;
        RECT 6.290 574.080 49.710 574.205 ;
      LAYER Pwell ;
        RECT 6.290 570.560 1143.390 574.080 ;
      LAYER Nwell ;
        RECT 6.290 570.435 28.155 570.560 ;
        RECT 6.290 566.365 1143.390 570.435 ;
        RECT 6.290 566.240 39.350 566.365 ;
      LAYER Pwell ;
        RECT 6.290 562.720 1143.390 566.240 ;
      LAYER Nwell ;
        RECT 6.290 562.595 17.020 562.720 ;
        RECT 6.290 558.525 1143.390 562.595 ;
        RECT 6.290 558.400 57.270 558.525 ;
      LAYER Pwell ;
        RECT 6.290 554.880 1143.390 558.400 ;
      LAYER Nwell ;
        RECT 6.290 554.755 27.415 554.880 ;
        RECT 6.290 550.685 1143.390 554.755 ;
        RECT 6.290 550.560 29.635 550.685 ;
      LAYER Pwell ;
        RECT 6.290 547.040 1143.390 550.560 ;
      LAYER Nwell ;
        RECT 6.290 546.915 22.305 547.040 ;
        RECT 6.290 542.845 1143.390 546.915 ;
        RECT 6.290 542.720 20.870 542.845 ;
      LAYER Pwell ;
        RECT 6.290 539.200 1143.390 542.720 ;
      LAYER Nwell ;
        RECT 6.290 539.075 17.960 539.200 ;
        RECT 6.290 535.005 1143.390 539.075 ;
        RECT 6.290 534.880 52.465 535.005 ;
      LAYER Pwell ;
        RECT 6.290 531.360 1143.390 534.880 ;
      LAYER Nwell ;
        RECT 6.290 531.235 183.505 531.360 ;
        RECT 6.290 527.165 1143.390 531.235 ;
        RECT 6.290 527.040 126.385 527.165 ;
      LAYER Pwell ;
        RECT 6.290 523.520 1143.390 527.040 ;
      LAYER Nwell ;
        RECT 6.290 523.395 17.960 523.520 ;
        RECT 6.290 519.325 1143.390 523.395 ;
        RECT 6.290 519.200 92.200 519.325 ;
      LAYER Pwell ;
        RECT 6.290 515.680 1143.390 519.200 ;
      LAYER Nwell ;
        RECT 6.290 515.555 70.945 515.680 ;
        RECT 6.290 511.485 1143.390 515.555 ;
        RECT 6.290 511.360 32.945 511.485 ;
      LAYER Pwell ;
        RECT 6.290 507.840 1143.390 511.360 ;
      LAYER Nwell ;
        RECT 6.290 507.715 189.745 507.840 ;
        RECT 6.290 503.645 1143.390 507.715 ;
        RECT 6.290 503.520 17.825 503.645 ;
      LAYER Pwell ;
        RECT 6.290 500.000 1143.390 503.520 ;
      LAYER Nwell ;
        RECT 6.290 499.875 17.960 500.000 ;
        RECT 6.290 495.805 1143.390 499.875 ;
        RECT 6.290 495.680 83.265 495.805 ;
      LAYER Pwell ;
        RECT 6.290 492.160 1143.390 495.680 ;
      LAYER Nwell ;
        RECT 6.290 492.035 16.390 492.160 ;
        RECT 6.290 487.965 1143.390 492.035 ;
        RECT 6.290 487.840 152.705 487.965 ;
      LAYER Pwell ;
        RECT 6.290 484.320 1143.390 487.840 ;
      LAYER Nwell ;
        RECT 6.290 484.195 71.830 484.320 ;
        RECT 6.290 480.125 1143.390 484.195 ;
        RECT 6.290 480.000 33.260 480.125 ;
      LAYER Pwell ;
        RECT 6.290 476.480 1143.390 480.000 ;
      LAYER Nwell ;
        RECT 6.290 476.355 52.105 476.480 ;
        RECT 6.290 472.285 1143.390 476.355 ;
        RECT 6.290 472.160 71.340 472.285 ;
      LAYER Pwell ;
        RECT 6.290 468.640 1143.390 472.160 ;
      LAYER Nwell ;
        RECT 6.290 468.515 114.755 468.640 ;
        RECT 6.290 464.445 1143.390 468.515 ;
        RECT 6.290 464.320 228.070 464.445 ;
      LAYER Pwell ;
        RECT 6.290 460.800 1143.390 464.320 ;
      LAYER Nwell ;
        RECT 6.290 460.675 29.505 460.800 ;
        RECT 6.290 456.605 1143.390 460.675 ;
        RECT 6.290 456.480 275.345 456.605 ;
      LAYER Pwell ;
        RECT 6.290 452.960 1143.390 456.480 ;
      LAYER Nwell ;
        RECT 6.290 452.835 12.705 452.960 ;
        RECT 6.290 448.765 1143.390 452.835 ;
        RECT 6.290 448.640 125.825 448.765 ;
      LAYER Pwell ;
        RECT 6.290 445.120 1143.390 448.640 ;
      LAYER Nwell ;
        RECT 6.290 444.995 177.345 445.120 ;
        RECT 6.290 440.925 1143.390 444.995 ;
        RECT 6.290 440.800 13.825 440.925 ;
      LAYER Pwell ;
        RECT 6.290 437.280 1143.390 440.800 ;
      LAYER Nwell ;
        RECT 6.290 437.155 51.670 437.280 ;
        RECT 6.290 433.085 1143.390 437.155 ;
        RECT 6.290 432.960 85.160 433.085 ;
      LAYER Pwell ;
        RECT 6.290 429.440 1143.390 432.960 ;
      LAYER Nwell ;
        RECT 6.290 429.315 14.710 429.440 ;
        RECT 6.290 425.245 1143.390 429.315 ;
        RECT 6.290 425.120 35.710 425.245 ;
      LAYER Pwell ;
        RECT 6.290 421.600 1143.390 425.120 ;
      LAYER Nwell ;
        RECT 6.290 421.475 99.545 421.600 ;
        RECT 6.290 417.405 1143.390 421.475 ;
        RECT 6.290 417.280 92.915 417.405 ;
      LAYER Pwell ;
        RECT 6.290 413.760 1143.390 417.280 ;
      LAYER Nwell ;
        RECT 6.290 413.635 96.360 413.760 ;
        RECT 6.290 409.565 1143.390 413.635 ;
        RECT 6.290 409.440 247.390 409.565 ;
      LAYER Pwell ;
        RECT 6.290 405.920 1143.390 409.440 ;
      LAYER Nwell ;
        RECT 6.290 405.795 32.865 405.920 ;
        RECT 6.290 401.725 1143.390 405.795 ;
        RECT 6.290 401.600 50.225 401.725 ;
      LAYER Pwell ;
        RECT 6.290 398.080 1143.390 401.600 ;
      LAYER Nwell ;
        RECT 6.290 397.955 32.865 398.080 ;
        RECT 6.290 393.885 1143.390 397.955 ;
        RECT 6.290 393.760 14.945 393.885 ;
      LAYER Pwell ;
        RECT 6.290 390.240 1143.390 393.760 ;
      LAYER Nwell ;
        RECT 6.290 390.115 61.985 390.240 ;
        RECT 6.290 386.045 1143.390 390.115 ;
        RECT 6.290 385.920 12.705 386.045 ;
      LAYER Pwell ;
        RECT 6.290 382.400 1143.390 385.920 ;
      LAYER Nwell ;
        RECT 6.290 382.275 57.720 382.400 ;
        RECT 6.290 378.205 1143.390 382.275 ;
        RECT 6.290 378.080 96.360 378.205 ;
      LAYER Pwell ;
        RECT 6.290 374.560 1143.390 378.080 ;
      LAYER Nwell ;
        RECT 6.290 374.435 73.745 374.560 ;
        RECT 6.290 370.365 1143.390 374.435 ;
        RECT 6.290 370.240 41.355 370.365 ;
      LAYER Pwell ;
        RECT 6.290 366.720 1143.390 370.240 ;
      LAYER Nwell ;
        RECT 6.290 366.595 74.910 366.720 ;
        RECT 6.290 362.525 1143.390 366.595 ;
        RECT 6.290 362.400 95.070 362.525 ;
      LAYER Pwell ;
        RECT 6.290 358.880 1143.390 362.400 ;
      LAYER Nwell ;
        RECT 6.290 358.755 26.250 358.880 ;
        RECT 6.290 354.685 1143.390 358.755 ;
        RECT 6.290 354.560 59.510 354.685 ;
      LAYER Pwell ;
        RECT 6.290 351.040 1143.390 354.560 ;
      LAYER Nwell ;
        RECT 6.290 350.915 11.070 351.040 ;
        RECT 6.290 346.845 1143.390 350.915 ;
        RECT 6.290 346.720 130.070 346.845 ;
      LAYER Pwell ;
        RECT 6.290 343.200 1143.390 346.720 ;
      LAYER Nwell ;
        RECT 6.290 343.075 57.830 343.200 ;
        RECT 6.290 339.005 1143.390 343.075 ;
        RECT 6.290 338.880 85.595 339.005 ;
      LAYER Pwell ;
        RECT 6.290 335.360 1143.390 338.880 ;
      LAYER Nwell ;
        RECT 6.290 335.235 210.710 335.360 ;
        RECT 6.290 331.165 1143.390 335.235 ;
        RECT 6.290 331.040 71.270 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 1143.390 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 33.505 327.520 ;
        RECT 6.290 323.325 1143.390 327.395 ;
        RECT 6.290 323.200 11.070 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 1143.390 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 198.390 319.680 ;
        RECT 6.290 315.485 1143.390 319.555 ;
        RECT 6.290 315.360 11.070 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 1143.390 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 19.470 311.840 ;
        RECT 6.290 307.645 1143.390 311.715 ;
        RECT 6.290 307.520 197.505 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 1143.390 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 33.470 304.000 ;
        RECT 6.290 299.805 1143.390 303.875 ;
        RECT 6.290 299.680 252.600 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 1143.390 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 217.845 296.160 ;
        RECT 6.290 291.965 1143.390 296.035 ;
        RECT 6.290 291.840 31.790 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 1143.390 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 33.515 288.320 ;
        RECT 6.290 284.125 1143.390 288.195 ;
        RECT 6.290 284.000 109.180 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 1143.390 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 11.630 280.480 ;
        RECT 6.290 276.285 1143.390 280.355 ;
        RECT 6.290 276.160 16.755 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1143.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 208.705 272.640 ;
        RECT 6.290 268.445 1143.390 272.515 ;
        RECT 6.290 268.320 48.590 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1143.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 69.920 264.800 ;
        RECT 6.290 260.605 1143.390 264.675 ;
        RECT 6.290 260.480 129.885 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1143.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 38.790 256.960 ;
        RECT 6.290 252.765 1143.390 256.835 ;
        RECT 6.290 252.640 217.285 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1143.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 108.465 249.120 ;
        RECT 6.290 244.925 1143.390 248.995 ;
        RECT 6.290 244.800 17.960 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1143.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 32.305 241.280 ;
        RECT 6.290 237.085 1143.390 241.155 ;
        RECT 6.290 236.960 32.305 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1143.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 12.705 233.440 ;
        RECT 6.290 229.245 1143.390 233.315 ;
        RECT 6.290 229.120 32.305 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1143.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 191.560 225.600 ;
        RECT 6.290 221.405 1143.390 225.475 ;
        RECT 6.290 221.280 85.505 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1143.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 12.705 217.760 ;
        RECT 6.290 213.565 1143.390 217.635 ;
        RECT 6.290 213.440 32.305 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1143.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 384.140 209.920 ;
        RECT 6.290 205.725 1143.390 209.795 ;
        RECT 6.290 205.600 49.105 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1143.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 28.945 202.080 ;
        RECT 6.290 197.885 1143.390 201.955 ;
        RECT 6.290 197.760 47.985 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1143.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 65.345 194.240 ;
        RECT 6.290 190.045 1143.390 194.115 ;
        RECT 6.290 189.920 83.265 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1143.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 110.360 186.400 ;
        RECT 6.290 182.205 1143.390 186.275 ;
        RECT 6.290 182.080 54.145 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1143.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 181.480 178.560 ;
        RECT 6.290 174.365 1143.390 178.435 ;
        RECT 6.290 174.240 48.760 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1143.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 61.425 170.720 ;
        RECT 6.290 166.525 1143.390 170.595 ;
        RECT 6.290 166.400 198.625 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1143.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 57.505 162.880 ;
        RECT 6.290 158.685 1143.390 162.755 ;
        RECT 6.290 158.560 37.345 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1143.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 139.825 155.040 ;
        RECT 6.290 150.845 1143.390 154.915 ;
        RECT 6.290 150.720 46.305 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1143.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 137.070 147.200 ;
        RECT 6.290 143.005 1143.390 147.075 ;
        RECT 6.290 142.880 32.305 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1143.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 51.905 139.360 ;
        RECT 6.290 135.165 1143.390 139.235 ;
        RECT 6.290 135.040 177.000 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1143.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 138.705 131.520 ;
        RECT 6.290 127.325 1143.390 131.395 ;
        RECT 6.290 127.200 49.665 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1143.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 152.145 123.680 ;
        RECT 6.290 119.485 1143.390 123.555 ;
        RECT 6.290 119.360 38.680 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1143.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 91.105 115.840 ;
        RECT 6.290 111.645 1143.390 115.715 ;
        RECT 6.290 111.520 71.505 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1143.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 92.785 108.000 ;
        RECT 6.290 103.805 1143.390 107.875 ;
        RECT 6.290 103.680 72.625 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1143.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 63.105 100.160 ;
        RECT 6.290 95.965 1143.390 100.035 ;
        RECT 6.290 95.840 163.905 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1143.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 73.185 92.320 ;
        RECT 6.290 88.125 1143.390 92.195 ;
        RECT 6.290 88.000 126.600 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1143.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 314.200 84.480 ;
        RECT 6.290 80.285 1143.390 84.355 ;
        RECT 6.290 80.160 59.400 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1143.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 143.745 76.640 ;
        RECT 6.290 72.445 1143.390 76.515 ;
        RECT 6.290 72.320 115.285 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1143.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 70.945 68.800 ;
        RECT 6.290 64.605 1143.390 68.675 ;
        RECT 6.290 64.480 85.505 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1143.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 311.400 60.960 ;
        RECT 6.290 56.765 1143.390 60.835 ;
        RECT 6.290 56.640 83.265 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1143.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 101.185 53.120 ;
        RECT 6.290 48.925 1143.390 52.995 ;
        RECT 6.290 48.800 192.100 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1143.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 100.625 45.280 ;
        RECT 6.290 41.085 1143.390 45.155 ;
        RECT 6.290 40.960 163.345 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1143.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 139.825 37.440 ;
        RECT 6.290 33.245 1143.390 37.315 ;
        RECT 6.290 33.120 93.345 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1143.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 112.945 29.600 ;
        RECT 6.290 25.405 1143.390 29.475 ;
        RECT 6.290 25.280 196.385 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1143.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 181.825 21.760 ;
        RECT 6.290 17.565 1143.390 21.635 ;
        RECT 6.290 17.440 412.545 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1143.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1142.960 784.300 ;
      LAYER Metal2 ;
        RECT 7.420 795.700 574.260 796.000 ;
        RECT 575.420 795.700 1142.820 796.000 ;
        RECT 7.420 4.300 1142.820 795.700 ;
        RECT 7.420 3.500 286.420 4.300 ;
        RECT 287.580 3.500 860.980 4.300 ;
        RECT 862.140 3.500 1142.820 4.300 ;
      LAYER Metal3 ;
        RECT 7.370 785.980 1146.000 793.380 ;
        RECT 7.370 784.820 1145.700 785.980 ;
        RECT 7.370 771.420 1146.000 784.820 ;
        RECT 7.370 770.260 1145.700 771.420 ;
        RECT 7.370 756.860 1146.000 770.260 ;
        RECT 7.370 755.700 1145.700 756.860 ;
        RECT 7.370 742.300 1146.000 755.700 ;
        RECT 7.370 741.140 1145.700 742.300 ;
        RECT 7.370 727.740 1146.000 741.140 ;
        RECT 7.370 726.580 1145.700 727.740 ;
        RECT 7.370 713.180 1146.000 726.580 ;
        RECT 7.370 712.020 1145.700 713.180 ;
        RECT 7.370 698.620 1146.000 712.020 ;
        RECT 7.370 697.460 1145.700 698.620 ;
        RECT 7.370 684.060 1146.000 697.460 ;
        RECT 7.370 682.900 1145.700 684.060 ;
        RECT 7.370 669.500 1146.000 682.900 ;
        RECT 7.370 668.340 1145.700 669.500 ;
        RECT 7.370 654.940 1146.000 668.340 ;
        RECT 7.370 653.780 1145.700 654.940 ;
        RECT 7.370 640.380 1146.000 653.780 ;
        RECT 7.370 639.220 1145.700 640.380 ;
        RECT 7.370 625.820 1146.000 639.220 ;
        RECT 7.370 624.660 1145.700 625.820 ;
        RECT 7.370 611.260 1146.000 624.660 ;
        RECT 7.370 610.100 1145.700 611.260 ;
        RECT 7.370 596.700 1146.000 610.100 ;
        RECT 7.370 595.540 1145.700 596.700 ;
        RECT 7.370 582.140 1146.000 595.540 ;
        RECT 7.370 580.980 1145.700 582.140 ;
        RECT 7.370 567.580 1146.000 580.980 ;
        RECT 7.370 566.420 1145.700 567.580 ;
        RECT 7.370 553.020 1146.000 566.420 ;
        RECT 7.370 551.860 1145.700 553.020 ;
        RECT 7.370 538.460 1146.000 551.860 ;
        RECT 7.370 537.300 1145.700 538.460 ;
        RECT 7.370 523.900 1146.000 537.300 ;
        RECT 7.370 522.740 1145.700 523.900 ;
        RECT 7.370 509.340 1146.000 522.740 ;
        RECT 7.370 508.180 1145.700 509.340 ;
        RECT 7.370 494.780 1146.000 508.180 ;
        RECT 7.370 493.620 1145.700 494.780 ;
        RECT 7.370 480.220 1146.000 493.620 ;
        RECT 7.370 479.060 1145.700 480.220 ;
        RECT 7.370 465.660 1146.000 479.060 ;
        RECT 7.370 464.500 1145.700 465.660 ;
        RECT 7.370 451.100 1146.000 464.500 ;
        RECT 7.370 449.940 1145.700 451.100 ;
        RECT 7.370 436.540 1146.000 449.940 ;
        RECT 7.370 435.380 1145.700 436.540 ;
        RECT 7.370 421.980 1146.000 435.380 ;
        RECT 7.370 420.820 1145.700 421.980 ;
        RECT 7.370 407.420 1146.000 420.820 ;
        RECT 7.370 406.260 1145.700 407.420 ;
        RECT 7.370 392.860 1146.000 406.260 ;
        RECT 7.370 391.700 1145.700 392.860 ;
        RECT 7.370 378.300 1146.000 391.700 ;
        RECT 7.370 377.140 1145.700 378.300 ;
        RECT 7.370 363.740 1146.000 377.140 ;
        RECT 7.370 362.580 1145.700 363.740 ;
        RECT 7.370 349.180 1146.000 362.580 ;
        RECT 7.370 348.020 1145.700 349.180 ;
        RECT 7.370 334.620 1146.000 348.020 ;
        RECT 7.370 333.460 1145.700 334.620 ;
        RECT 7.370 320.060 1146.000 333.460 ;
        RECT 7.370 318.900 1145.700 320.060 ;
        RECT 7.370 305.500 1146.000 318.900 ;
        RECT 7.370 304.340 1145.700 305.500 ;
        RECT 7.370 290.940 1146.000 304.340 ;
        RECT 7.370 289.780 1145.700 290.940 ;
        RECT 7.370 276.380 1146.000 289.780 ;
        RECT 7.370 275.220 1145.700 276.380 ;
        RECT 7.370 261.820 1146.000 275.220 ;
        RECT 7.370 260.660 1145.700 261.820 ;
        RECT 7.370 247.260 1146.000 260.660 ;
        RECT 7.370 246.100 1145.700 247.260 ;
        RECT 7.370 232.700 1146.000 246.100 ;
        RECT 7.370 231.540 1145.700 232.700 ;
        RECT 7.370 218.140 1146.000 231.540 ;
        RECT 7.370 216.980 1145.700 218.140 ;
        RECT 7.370 203.580 1146.000 216.980 ;
        RECT 7.370 202.420 1145.700 203.580 ;
        RECT 7.370 189.020 1146.000 202.420 ;
        RECT 7.370 187.860 1145.700 189.020 ;
        RECT 7.370 174.460 1146.000 187.860 ;
        RECT 7.370 173.300 1145.700 174.460 ;
        RECT 7.370 159.900 1146.000 173.300 ;
        RECT 7.370 158.740 1145.700 159.900 ;
        RECT 7.370 145.340 1146.000 158.740 ;
        RECT 7.370 144.180 1145.700 145.340 ;
        RECT 7.370 130.780 1146.000 144.180 ;
        RECT 7.370 129.620 1145.700 130.780 ;
        RECT 7.370 116.220 1146.000 129.620 ;
        RECT 7.370 115.060 1145.700 116.220 ;
        RECT 7.370 101.660 1146.000 115.060 ;
        RECT 7.370 100.500 1145.700 101.660 ;
        RECT 7.370 87.100 1146.000 100.500 ;
        RECT 7.370 85.940 1145.700 87.100 ;
        RECT 7.370 72.540 1146.000 85.940 ;
        RECT 7.370 71.380 1145.700 72.540 ;
        RECT 7.370 57.980 1146.000 71.380 ;
        RECT 7.370 56.820 1145.700 57.980 ;
        RECT 7.370 43.420 1146.000 56.820 ;
        RECT 7.370 42.260 1145.700 43.420 ;
        RECT 7.370 28.860 1146.000 42.260 ;
        RECT 7.370 27.700 1145.700 28.860 ;
        RECT 7.370 14.300 1146.000 27.700 ;
        RECT 7.370 13.140 1145.700 14.300 ;
        RECT 7.370 4.060 1146.000 13.140 ;
      LAYER Metal4 ;
        RECT 21.420 784.600 1133.860 792.310 ;
        RECT 21.420 15.080 21.940 784.600 ;
        RECT 24.140 15.080 98.740 784.600 ;
        RECT 100.940 15.080 175.540 784.600 ;
        RECT 177.740 15.080 252.340 784.600 ;
        RECT 254.540 15.080 329.140 784.600 ;
        RECT 331.340 15.080 405.940 784.600 ;
        RECT 408.140 15.080 482.740 784.600 ;
        RECT 484.940 15.080 559.540 784.600 ;
        RECT 561.740 15.080 636.340 784.600 ;
        RECT 638.540 15.080 713.140 784.600 ;
        RECT 715.340 15.080 789.940 784.600 ;
        RECT 792.140 15.080 866.740 784.600 ;
        RECT 868.940 15.080 943.540 784.600 ;
        RECT 945.740 15.080 1020.340 784.600 ;
        RECT 1022.540 15.080 1097.140 784.600 ;
        RECT 1099.340 15.080 1133.860 784.600 ;
        RECT 21.420 5.130 1133.860 15.080 ;
  END
END wrapped_sid
END LIBRARY

