magic
tech gf180mcuD
magscale 1 10
timestamp 1702341871
<< nwell >>
rect 1258 33305 35702 33798
rect 1258 33280 13965 33305
rect 1258 32551 6909 32576
rect 1258 31737 35702 32551
rect 1258 31712 9373 31737
rect 1258 30983 5229 31008
rect 1258 30169 35702 30983
rect 1258 30144 24941 30169
rect 1258 29415 4669 29440
rect 1258 28576 35702 29415
rect 1258 27847 4333 27872
rect 1258 27033 35702 27847
rect 1258 27008 9382 27033
rect 1258 26279 4445 26304
rect 1258 25465 35702 26279
rect 1258 25440 24269 25465
rect 1258 24711 26061 24736
rect 1258 23897 35702 24711
rect 1258 23872 33117 23897
rect 1258 23143 4781 23168
rect 1258 22329 35702 23143
rect 1258 22304 8253 22329
rect 1258 21575 4445 21600
rect 1258 20761 35702 21575
rect 1258 20736 10717 20761
rect 1258 20007 5789 20032
rect 1258 19193 35702 20007
rect 1258 19168 6461 19193
rect 1258 18439 14749 18464
rect 1258 17625 35702 18439
rect 1258 17600 8141 17625
rect 1258 16871 12733 16896
rect 1258 16057 35702 16871
rect 1258 16032 10829 16057
rect 1258 15303 18701 15328
rect 1258 14489 35702 15303
rect 1258 14464 14525 14489
rect 1258 13735 10381 13760
rect 1258 12921 35702 13735
rect 1258 12896 26552 12921
rect 1258 12167 6728 12192
rect 1258 11353 35702 12167
rect 1258 11328 7512 11353
rect 1258 10599 13181 10624
rect 1258 9785 35702 10599
rect 1258 9760 7805 9785
rect 1258 9031 6056 9056
rect 1258 8217 35702 9031
rect 1258 8192 11656 8217
rect 1258 7463 12957 7488
rect 1258 6649 35702 7463
rect 1258 6624 16920 6649
rect 1258 5895 12509 5920
rect 1258 5081 35702 5895
rect 1258 5056 6909 5081
rect 1258 4327 6685 4352
rect 1258 3488 35702 4327
<< pwell >>
rect 1258 32576 35702 33280
rect 1258 31008 35702 31712
rect 1258 29440 35702 30144
rect 1258 27872 35702 28576
rect 1258 26304 35702 27008
rect 1258 24736 35702 25440
rect 1258 23168 35702 23872
rect 1258 21600 35702 22304
rect 1258 20032 35702 20736
rect 1258 18464 35702 19168
rect 1258 16896 35702 17600
rect 1258 15328 35702 16032
rect 1258 13760 35702 14464
rect 1258 12192 35702 12896
rect 1258 10624 35702 11328
rect 1258 9056 35702 9760
rect 1258 7488 35702 8192
rect 1258 5920 35702 6624
rect 1258 4352 35702 5056
rect 1258 3050 35702 3488
<< obsm1 >>
rect 1344 3076 35776 33772
<< metal2 >>
rect 1568 36200 1680 37000
rect 2688 36200 2800 37000
rect 3808 36200 3920 37000
rect 4928 36200 5040 37000
rect 6048 36200 6160 37000
rect 7168 36200 7280 37000
rect 8288 36200 8400 37000
rect 9408 36200 9520 37000
rect 10528 36200 10640 37000
rect 11648 36200 11760 37000
rect 12768 36200 12880 37000
rect 13888 36200 14000 37000
rect 15008 36200 15120 37000
rect 16128 36200 16240 37000
rect 17248 36200 17360 37000
rect 18368 36200 18480 37000
rect 19488 36200 19600 37000
rect 20608 36200 20720 37000
rect 21728 36200 21840 37000
rect 22848 36200 22960 37000
rect 23968 36200 24080 37000
rect 25088 36200 25200 37000
rect 26208 36200 26320 37000
rect 27328 36200 27440 37000
rect 28448 36200 28560 37000
rect 29568 36200 29680 37000
rect 30688 36200 30800 37000
rect 31808 36200 31920 37000
rect 32928 36200 33040 37000
rect 34048 36200 34160 37000
rect 35168 36200 35280 37000
rect 1792 0 1904 800
rect 3360 0 3472 800
rect 4928 0 5040 800
rect 6496 0 6608 800
rect 8064 0 8176 800
rect 9632 0 9744 800
rect 11200 0 11312 800
rect 12768 0 12880 800
rect 14336 0 14448 800
rect 15904 0 16016 800
rect 17472 0 17584 800
rect 19040 0 19152 800
rect 20608 0 20720 800
rect 22176 0 22288 800
rect 23744 0 23856 800
rect 25312 0 25424 800
rect 26880 0 26992 800
rect 28448 0 28560 800
rect 30016 0 30128 800
rect 31584 0 31696 800
rect 33152 0 33264 800
rect 34720 0 34832 800
<< obsm2 >>
rect 1740 36140 2628 36260
rect 2860 36140 3748 36260
rect 3980 36140 4868 36260
rect 5100 36140 5988 36260
rect 6220 36140 7108 36260
rect 7340 36140 8228 36260
rect 8460 36140 9348 36260
rect 9580 36140 10468 36260
rect 10700 36140 11588 36260
rect 11820 36140 12708 36260
rect 12940 36140 13828 36260
rect 14060 36140 14948 36260
rect 15180 36140 16068 36260
rect 16300 36140 17188 36260
rect 17420 36140 18308 36260
rect 18540 36140 19428 36260
rect 19660 36140 20548 36260
rect 20780 36140 21668 36260
rect 21900 36140 22788 36260
rect 23020 36140 23908 36260
rect 24140 36140 25028 36260
rect 25260 36140 26148 36260
rect 26380 36140 27268 36260
rect 27500 36140 28388 36260
rect 28620 36140 29508 36260
rect 29740 36140 30628 36260
rect 30860 36140 31748 36260
rect 31980 36140 32868 36260
rect 33100 36140 33988 36260
rect 34220 36140 35108 36260
rect 35340 36140 36260 36260
rect 1596 860 36260 36140
rect 1596 800 1732 860
rect 1964 800 3300 860
rect 3532 800 4868 860
rect 5100 800 6436 860
rect 6668 800 8004 860
rect 8236 800 9572 860
rect 9804 800 11140 860
rect 11372 800 12708 860
rect 12940 800 14276 860
rect 14508 800 15844 860
rect 16076 800 17412 860
rect 17644 800 18980 860
rect 19212 800 20548 860
rect 20780 800 22116 860
rect 22348 800 23684 860
rect 23916 800 25252 860
rect 25484 800 26820 860
rect 27052 800 28388 860
rect 28620 800 29956 860
rect 30188 800 31524 860
rect 31756 800 33092 860
rect 33324 800 34660 860
rect 34892 800 36260 860
<< metal3 >>
rect 36200 34496 37000 34608
rect 36200 31808 37000 31920
rect 36200 29120 37000 29232
rect 36200 26432 37000 26544
rect 36200 23744 37000 23856
rect 36200 21056 37000 21168
rect 36200 18368 37000 18480
rect 36200 15680 37000 15792
rect 36200 12992 37000 13104
rect 36200 10304 37000 10416
rect 36200 7616 37000 7728
rect 36200 4928 37000 5040
rect 36200 2240 37000 2352
<< obsm3 >>
rect 3602 34436 36140 34580
rect 3602 31980 36270 34436
rect 3602 31748 36140 31980
rect 3602 29292 36270 31748
rect 3602 29060 36140 29292
rect 3602 26604 36270 29060
rect 3602 26372 36140 26604
rect 3602 23916 36270 26372
rect 3602 23684 36140 23916
rect 3602 21228 36270 23684
rect 3602 20996 36140 21228
rect 3602 18540 36270 20996
rect 3602 18308 36140 18540
rect 3602 15852 36270 18308
rect 3602 15620 36140 15852
rect 3602 13164 36270 15620
rect 3602 12932 36140 13164
rect 3602 10476 36270 12932
rect 3602 10244 36140 10476
rect 3602 7788 36270 10244
rect 3602 7556 36140 7788
rect 3602 5100 36270 7556
rect 3602 4868 36140 5100
rect 3602 2412 36270 4868
rect 3602 2268 36140 2412
<< metal4 >>
rect 5468 3076 5788 33772
rect 9752 3076 10072 33772
rect 14036 3076 14356 33772
rect 18320 3076 18640 33772
rect 22604 3076 22924 33772
rect 26888 3076 27208 33772
rect 31172 3076 31492 33772
rect 35456 3076 35776 33772
<< obsm4 >>
rect 7644 5282 9692 31118
rect 10132 5282 13976 31118
rect 14416 5282 18260 31118
rect 18700 5282 22544 31118
rect 22984 5282 26828 31118
rect 27268 5282 31112 31118
rect 31552 5282 35140 31118
<< labels >>
rlabel metal3 s 36200 29120 37000 29232 6 SDI
port 1 nsew signal input
rlabel metal3 s 36200 2240 37000 2352 6 clk_i
port 2 nsew signal input
rlabel metal3 s 36200 34496 37000 34608 6 custom_setting
port 3 nsew signal input
rlabel metal3 s 36200 7616 37000 7728 6 io_in[0]
port 4 nsew signal input
rlabel metal3 s 36200 10304 37000 10416 6 io_in[1]
port 5 nsew signal input
rlabel metal3 s 36200 12992 37000 13104 6 io_in[2]
port 6 nsew signal input
rlabel metal3 s 36200 15680 37000 15792 6 io_in[3]
port 7 nsew signal input
rlabel metal3 s 36200 18368 37000 18480 6 io_in[4]
port 8 nsew signal input
rlabel metal3 s 36200 21056 37000 21168 6 io_in[5]
port 9 nsew signal input
rlabel metal3 s 36200 23744 37000 23856 6 io_in[6]
port 10 nsew signal input
rlabel metal3 s 36200 26432 37000 26544 6 io_in[7]
port 11 nsew signal input
rlabel metal2 s 1568 36200 1680 37000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 12768 36200 12880 37000 6 io_out[10]
port 13 nsew signal output
rlabel metal2 s 13888 36200 14000 37000 6 io_out[11]
port 14 nsew signal output
rlabel metal2 s 15008 36200 15120 37000 6 io_out[12]
port 15 nsew signal output
rlabel metal2 s 16128 36200 16240 37000 6 io_out[13]
port 16 nsew signal output
rlabel metal2 s 17248 36200 17360 37000 6 io_out[14]
port 17 nsew signal output
rlabel metal2 s 18368 36200 18480 37000 6 io_out[15]
port 18 nsew signal output
rlabel metal2 s 19488 36200 19600 37000 6 io_out[16]
port 19 nsew signal output
rlabel metal2 s 20608 36200 20720 37000 6 io_out[17]
port 20 nsew signal output
rlabel metal2 s 21728 36200 21840 37000 6 io_out[18]
port 21 nsew signal output
rlabel metal2 s 22848 36200 22960 37000 6 io_out[19]
port 22 nsew signal output
rlabel metal2 s 2688 36200 2800 37000 6 io_out[1]
port 23 nsew signal output
rlabel metal2 s 23968 36200 24080 37000 6 io_out[20]
port 24 nsew signal output
rlabel metal2 s 25088 36200 25200 37000 6 io_out[21]
port 25 nsew signal output
rlabel metal2 s 26208 36200 26320 37000 6 io_out[22]
port 26 nsew signal output
rlabel metal2 s 27328 36200 27440 37000 6 io_out[23]
port 27 nsew signal output
rlabel metal2 s 28448 36200 28560 37000 6 io_out[24]
port 28 nsew signal output
rlabel metal2 s 29568 36200 29680 37000 6 io_out[25]
port 29 nsew signal output
rlabel metal2 s 30688 36200 30800 37000 6 io_out[26]
port 30 nsew signal output
rlabel metal2 s 31808 36200 31920 37000 6 io_out[27]
port 31 nsew signal output
rlabel metal2 s 32928 36200 33040 37000 6 io_out[28]
port 32 nsew signal output
rlabel metal2 s 34048 36200 34160 37000 6 io_out[29]
port 33 nsew signal output
rlabel metal2 s 3808 36200 3920 37000 6 io_out[2]
port 34 nsew signal output
rlabel metal2 s 35168 36200 35280 37000 6 io_out[30]
port 35 nsew signal output
rlabel metal2 s 4928 36200 5040 37000 6 io_out[3]
port 36 nsew signal output
rlabel metal2 s 6048 36200 6160 37000 6 io_out[4]
port 37 nsew signal output
rlabel metal2 s 7168 36200 7280 37000 6 io_out[5]
port 38 nsew signal output
rlabel metal2 s 8288 36200 8400 37000 6 io_out[6]
port 39 nsew signal output
rlabel metal2 s 9408 36200 9520 37000 6 io_out[7]
port 40 nsew signal output
rlabel metal2 s 10528 36200 10640 37000 6 io_out[8]
port 41 nsew signal output
rlabel metal2 s 11648 36200 11760 37000 6 io_out[9]
port 42 nsew signal output
rlabel metal3 s 36200 4928 37000 5040 6 rst_n
port 43 nsew signal input
rlabel metal2 s 1792 0 1904 800 6 sram_addr[0]
port 44 nsew signal output
rlabel metal2 s 3360 0 3472 800 6 sram_addr[1]
port 45 nsew signal output
rlabel metal2 s 4928 0 5040 800 6 sram_addr[2]
port 46 nsew signal output
rlabel metal2 s 6496 0 6608 800 6 sram_addr[3]
port 47 nsew signal output
rlabel metal2 s 8064 0 8176 800 6 sram_addr[4]
port 48 nsew signal output
rlabel metal2 s 9632 0 9744 800 6 sram_addr[5]
port 49 nsew signal output
rlabel metal3 s 36200 31808 37000 31920 6 sram_gwe
port 50 nsew signal output
rlabel metal2 s 11200 0 11312 800 6 sram_in[0]
port 51 nsew signal output
rlabel metal2 s 12768 0 12880 800 6 sram_in[1]
port 52 nsew signal output
rlabel metal2 s 14336 0 14448 800 6 sram_in[2]
port 53 nsew signal output
rlabel metal2 s 15904 0 16016 800 6 sram_in[3]
port 54 nsew signal output
rlabel metal2 s 17472 0 17584 800 6 sram_in[4]
port 55 nsew signal output
rlabel metal2 s 19040 0 19152 800 6 sram_in[5]
port 56 nsew signal output
rlabel metal2 s 20608 0 20720 800 6 sram_in[6]
port 57 nsew signal output
rlabel metal2 s 22176 0 22288 800 6 sram_in[7]
port 58 nsew signal output
rlabel metal2 s 23744 0 23856 800 6 sram_out[0]
port 59 nsew signal input
rlabel metal2 s 25312 0 25424 800 6 sram_out[1]
port 60 nsew signal input
rlabel metal2 s 26880 0 26992 800 6 sram_out[2]
port 61 nsew signal input
rlabel metal2 s 28448 0 28560 800 6 sram_out[3]
port 62 nsew signal input
rlabel metal2 s 30016 0 30128 800 6 sram_out[4]
port 63 nsew signal input
rlabel metal2 s 31584 0 31696 800 6 sram_out[5]
port 64 nsew signal input
rlabel metal2 s 33152 0 33264 800 6 sram_out[6]
port 65 nsew signal input
rlabel metal2 s 34720 0 34832 800 6 sram_out[7]
port 66 nsew signal input
rlabel metal4 s 5468 3076 5788 33772 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 14036 3076 14356 33772 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 22604 3076 22924 33772 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 31172 3076 31492 33772 6 vdd
port 67 nsew power bidirectional
rlabel metal4 s 9752 3076 10072 33772 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 18320 3076 18640 33772 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 26888 3076 27208 33772 6 vss
port 68 nsew ground bidirectional
rlabel metal4 s 35456 3076 35776 33772 6 vss
port 68 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 37000 37000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1370914
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_mc14500/runs/23_12_12_01_41/results/signoff/wrapped_mc14500.magic.gds
string GDS_START 268356
<< end >>

