magic
tech gf180mcuD
magscale 1 10
timestamp 1702341366
<< metal1 >>
rect 13570 44830 13582 44882
rect 13634 44879 13646 44882
rect 14466 44879 14478 44882
rect 13634 44833 14478 44879
rect 13634 44830 13646 44833
rect 14466 44830 14478 44833
rect 14530 44830 14542 44882
rect 1344 44714 46592 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 46592 44714
rect 1344 44628 46592 44662
rect 31278 44546 31330 44558
rect 31278 44482 31330 44494
rect 14478 44434 14530 44446
rect 10098 44382 10110 44434
rect 10162 44382 10174 44434
rect 14478 44370 14530 44382
rect 14590 44434 14642 44446
rect 14590 44370 14642 44382
rect 15598 44434 15650 44446
rect 20078 44434 20130 44446
rect 23550 44434 23602 44446
rect 29150 44434 29202 44446
rect 15810 44382 15822 44434
rect 15874 44382 15886 44434
rect 23090 44382 23102 44434
rect 23154 44382 23166 44434
rect 27794 44382 27806 44434
rect 27858 44382 27870 44434
rect 32498 44382 32510 44434
rect 32562 44382 32574 44434
rect 39218 44382 39230 44434
rect 39282 44382 39294 44434
rect 43026 44382 43038 44434
rect 43090 44382 43102 44434
rect 15598 44370 15650 44382
rect 20078 44370 20130 44382
rect 23550 44370 23602 44382
rect 29150 44370 29202 44382
rect 13582 44322 13634 44334
rect 13582 44258 13634 44270
rect 14142 44322 14194 44334
rect 14142 44258 14194 44270
rect 17502 44322 17554 44334
rect 17502 44258 17554 44270
rect 18174 44322 18226 44334
rect 18174 44258 18226 44270
rect 18734 44322 18786 44334
rect 18734 44258 18786 44270
rect 21758 44322 21810 44334
rect 21758 44258 21810 44270
rect 22766 44322 22818 44334
rect 30046 44322 30098 44334
rect 24994 44270 25006 44322
rect 25058 44270 25070 44322
rect 22766 44258 22818 44270
rect 30046 44258 30098 44270
rect 30606 44322 30658 44334
rect 30606 44258 30658 44270
rect 34526 44322 34578 44334
rect 34850 44270 34862 44322
rect 34914 44270 34926 44322
rect 36418 44270 36430 44322
rect 36482 44270 36494 44322
rect 40114 44270 40126 44322
rect 40178 44270 40190 44322
rect 45154 44270 45166 44322
rect 45218 44270 45230 44322
rect 34526 44258 34578 44270
rect 9774 44210 9826 44222
rect 9774 44146 9826 44158
rect 13694 44210 13746 44222
rect 13694 44146 13746 44158
rect 16158 44210 16210 44222
rect 16158 44146 16210 44158
rect 20190 44210 20242 44222
rect 20190 44146 20242 44158
rect 20750 44210 20802 44222
rect 20750 44146 20802 44158
rect 21534 44210 21586 44222
rect 21534 44146 21586 44158
rect 21870 44210 21922 44222
rect 21870 44146 21922 44158
rect 22542 44210 22594 44222
rect 29710 44210 29762 44222
rect 25666 44158 25678 44210
rect 25730 44158 25742 44210
rect 22542 44146 22594 44158
rect 29710 44146 29762 44158
rect 30942 44210 30994 44222
rect 30942 44146 30994 44158
rect 32174 44210 32226 44222
rect 32174 44146 32226 44158
rect 33406 44210 33458 44222
rect 33406 44146 33458 44158
rect 33518 44210 33570 44222
rect 33518 44146 33570 44158
rect 33854 44210 33906 44222
rect 33854 44146 33906 44158
rect 35422 44210 35474 44222
rect 43598 44210 43650 44222
rect 37090 44158 37102 44210
rect 37154 44158 37166 44210
rect 40898 44158 40910 44210
rect 40962 44158 40974 44210
rect 35422 44146 35474 44158
rect 43598 44146 43650 44158
rect 44270 44210 44322 44222
rect 44930 44158 44942 44210
rect 44994 44158 45006 44210
rect 44270 44146 44322 44158
rect 9550 44098 9602 44110
rect 9550 44034 9602 44046
rect 9998 44098 10050 44110
rect 9998 44034 10050 44046
rect 13806 44098 13858 44110
rect 13806 44034 13858 44046
rect 15150 44098 15202 44110
rect 15150 44034 15202 44046
rect 15934 44098 15986 44110
rect 15934 44034 15986 44046
rect 17950 44098 18002 44110
rect 17950 44034 18002 44046
rect 19294 44098 19346 44110
rect 19294 44034 19346 44046
rect 19854 44098 19906 44110
rect 19854 44034 19906 44046
rect 20862 44098 20914 44110
rect 20862 44034 20914 44046
rect 21086 44098 21138 44110
rect 21086 44034 21138 44046
rect 21982 44098 22034 44110
rect 21982 44034 22034 44046
rect 22094 44098 22146 44110
rect 22094 44034 22146 44046
rect 22990 44098 23042 44110
rect 22990 44034 23042 44046
rect 23102 44098 23154 44110
rect 23102 44034 23154 44046
rect 23662 44098 23714 44110
rect 23662 44034 23714 44046
rect 28702 44098 28754 44110
rect 28702 44034 28754 44046
rect 29486 44098 29538 44110
rect 29486 44034 29538 44046
rect 29598 44098 29650 44110
rect 29598 44034 29650 44046
rect 31166 44098 31218 44110
rect 31166 44034 31218 44046
rect 32398 44098 32450 44110
rect 32398 44034 32450 44046
rect 33182 44098 33234 44110
rect 33182 44034 33234 44046
rect 33966 44098 34018 44110
rect 33966 44034 34018 44046
rect 34190 44098 34242 44110
rect 34190 44034 34242 44046
rect 43710 44098 43762 44110
rect 43710 44034 43762 44046
rect 44382 44098 44434 44110
rect 44382 44034 44434 44046
rect 44494 44098 44546 44110
rect 45950 44098 46002 44110
rect 45602 44046 45614 44098
rect 45666 44046 45678 44098
rect 44494 44034 44546 44046
rect 45950 44034 46002 44046
rect 1344 43930 46592 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 46592 43930
rect 1344 43844 46592 43878
rect 8866 43710 8878 43762
rect 8930 43710 8942 43762
rect 29474 43710 29486 43762
rect 29538 43710 29550 43762
rect 29150 43650 29202 43662
rect 19058 43598 19070 43650
rect 19122 43598 19134 43650
rect 23874 43598 23886 43650
rect 23938 43598 23950 43650
rect 29150 43586 29202 43598
rect 30158 43650 30210 43662
rect 32622 43650 32674 43662
rect 31042 43598 31054 43650
rect 31106 43598 31118 43650
rect 30158 43586 30210 43598
rect 32622 43586 32674 43598
rect 39902 43650 39954 43662
rect 39902 43586 39954 43598
rect 10110 43538 10162 43550
rect 25230 43538 25282 43550
rect 29822 43538 29874 43550
rect 5954 43486 5966 43538
rect 6018 43486 6030 43538
rect 10770 43486 10782 43538
rect 10834 43486 10846 43538
rect 14018 43486 14030 43538
rect 14082 43486 14094 43538
rect 17602 43486 17614 43538
rect 17666 43486 17678 43538
rect 18386 43486 18398 43538
rect 18450 43486 18462 43538
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 25666 43486 25678 43538
rect 25730 43486 25742 43538
rect 10110 43474 10162 43486
rect 25230 43474 25282 43486
rect 29822 43474 29874 43486
rect 30718 43538 30770 43550
rect 30718 43474 30770 43486
rect 31726 43538 31778 43550
rect 31726 43474 31778 43486
rect 31838 43538 31890 43550
rect 39454 43538 39506 43550
rect 35970 43486 35982 43538
rect 36034 43486 36046 43538
rect 36418 43486 36430 43538
rect 36482 43486 36494 43538
rect 31838 43474 31890 43486
rect 39454 43474 39506 43486
rect 40014 43538 40066 43550
rect 40014 43474 40066 43486
rect 41022 43538 41074 43550
rect 41022 43474 41074 43486
rect 41134 43538 41186 43550
rect 41134 43474 41186 43486
rect 41246 43538 41298 43550
rect 41246 43474 41298 43486
rect 42142 43538 42194 43550
rect 42142 43474 42194 43486
rect 42366 43538 42418 43550
rect 43250 43486 43262 43538
rect 43314 43486 43326 43538
rect 42366 43474 42418 43486
rect 17838 43426 17890 43438
rect 30494 43426 30546 43438
rect 6626 43374 6638 43426
rect 6690 43374 6702 43426
rect 11442 43374 11454 43426
rect 11506 43374 11518 43426
rect 13570 43374 13582 43426
rect 13634 43374 13646 43426
rect 14690 43374 14702 43426
rect 14754 43374 14766 43426
rect 16818 43374 16830 43426
rect 16882 43374 16894 43426
rect 21186 43374 21198 43426
rect 21250 43374 21262 43426
rect 21634 43374 21646 43426
rect 21698 43374 21710 43426
rect 26450 43374 26462 43426
rect 26514 43374 26526 43426
rect 28578 43374 28590 43426
rect 28642 43374 28654 43426
rect 17838 43362 17890 43374
rect 30494 43362 30546 43374
rect 31390 43426 31442 43438
rect 39678 43426 39730 43438
rect 33058 43374 33070 43426
rect 33122 43374 33134 43426
rect 35186 43374 35198 43426
rect 35250 43374 35262 43426
rect 37090 43374 37102 43426
rect 37154 43374 37166 43426
rect 39218 43374 39230 43426
rect 39282 43374 39294 43426
rect 44034 43374 44046 43426
rect 44098 43374 44110 43426
rect 46162 43374 46174 43426
rect 46226 43374 46238 43426
rect 31390 43362 31442 43374
rect 39678 43362 39730 43374
rect 9886 43314 9938 43326
rect 9538 43262 9550 43314
rect 9602 43262 9614 43314
rect 9886 43250 9938 43262
rect 17950 43314 18002 43326
rect 17950 43250 18002 43262
rect 25342 43314 25394 43326
rect 25342 43250 25394 43262
rect 31502 43314 31554 43326
rect 42030 43314 42082 43326
rect 41682 43262 41694 43314
rect 41746 43262 41758 43314
rect 31502 43250 31554 43262
rect 42030 43250 42082 43262
rect 42478 43314 42530 43326
rect 42478 43250 42530 43262
rect 1344 43146 46592 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 46592 43146
rect 1344 43060 46592 43094
rect 9998 42978 10050 42990
rect 9998 42914 10050 42926
rect 10670 42978 10722 42990
rect 10670 42914 10722 42926
rect 11006 42978 11058 42990
rect 11006 42914 11058 42926
rect 11342 42978 11394 42990
rect 11342 42914 11394 42926
rect 11678 42978 11730 42990
rect 14814 42978 14866 42990
rect 32510 42978 32562 42990
rect 13458 42926 13470 42978
rect 13522 42926 13534 42978
rect 20066 42926 20078 42978
rect 20130 42926 20142 42978
rect 31042 42926 31054 42978
rect 31106 42926 31118 42978
rect 11678 42914 11730 42926
rect 14814 42914 14866 42926
rect 32510 42914 32562 42926
rect 32846 42978 32898 42990
rect 32846 42914 32898 42926
rect 35310 42978 35362 42990
rect 35310 42914 35362 42926
rect 35646 42978 35698 42990
rect 35646 42914 35698 42926
rect 38446 42978 38498 42990
rect 38446 42914 38498 42926
rect 39118 42978 39170 42990
rect 39118 42914 39170 42926
rect 9214 42866 9266 42878
rect 26462 42866 26514 42878
rect 18610 42814 18622 42866
rect 18674 42814 18686 42866
rect 19282 42814 19294 42866
rect 19346 42814 19358 42866
rect 21746 42814 21758 42866
rect 21810 42814 21822 42866
rect 24770 42814 24782 42866
rect 24834 42814 24846 42866
rect 9214 42802 9266 42814
rect 26462 42802 26514 42814
rect 29262 42866 29314 42878
rect 29262 42802 29314 42814
rect 30494 42866 30546 42878
rect 33506 42814 33518 42866
rect 33570 42814 33582 42866
rect 39442 42814 39454 42866
rect 39506 42814 39518 42866
rect 41570 42814 41582 42866
rect 41634 42814 41646 42866
rect 42802 42814 42814 42866
rect 42866 42814 42878 42866
rect 30494 42802 30546 42814
rect 9662 42754 9714 42766
rect 9662 42690 9714 42702
rect 9886 42754 9938 42766
rect 9886 42690 9938 42702
rect 10558 42754 10610 42766
rect 10558 42690 10610 42702
rect 10894 42754 10946 42766
rect 10894 42690 10946 42702
rect 11454 42754 11506 42766
rect 13918 42754 13970 42766
rect 11890 42702 11902 42754
rect 11954 42702 11966 42754
rect 11454 42690 11506 42702
rect 13918 42690 13970 42702
rect 14142 42754 14194 42766
rect 14142 42690 14194 42702
rect 14926 42754 14978 42766
rect 14926 42690 14978 42702
rect 15150 42754 15202 42766
rect 20638 42754 20690 42766
rect 26350 42754 26402 42766
rect 15362 42702 15374 42754
rect 15426 42702 15438 42754
rect 15810 42702 15822 42754
rect 15874 42702 15886 42754
rect 19170 42702 19182 42754
rect 19234 42702 19246 42754
rect 20402 42702 20414 42754
rect 20466 42702 20478 42754
rect 21858 42702 21870 42754
rect 21922 42702 21934 42754
rect 22866 42702 22878 42754
rect 22930 42702 22942 42754
rect 23538 42702 23550 42754
rect 23602 42702 23614 42754
rect 24322 42702 24334 42754
rect 24386 42702 24398 42754
rect 15150 42690 15202 42702
rect 20638 42690 20690 42702
rect 26350 42690 26402 42702
rect 26686 42754 26738 42766
rect 26686 42690 26738 42702
rect 29486 42754 29538 42766
rect 29486 42690 29538 42702
rect 30046 42754 30098 42766
rect 30046 42690 30098 42702
rect 30718 42754 30770 42766
rect 30718 42690 30770 42702
rect 32398 42754 32450 42766
rect 32398 42690 32450 42702
rect 32734 42754 32786 42766
rect 37550 42754 37602 42766
rect 35634 42702 35646 42754
rect 35698 42702 35710 42754
rect 36082 42702 36094 42754
rect 36146 42702 36158 42754
rect 32734 42690 32786 42702
rect 37550 42690 37602 42702
rect 37774 42754 37826 42766
rect 38558 42754 38610 42766
rect 37986 42702 37998 42754
rect 38050 42702 38062 42754
rect 37774 42690 37826 42702
rect 38558 42690 38610 42702
rect 38782 42754 38834 42766
rect 38782 42690 38834 42702
rect 39006 42754 39058 42766
rect 45278 42754 45330 42766
rect 42354 42702 42366 42754
rect 42418 42702 42430 42754
rect 43026 42702 43038 42754
rect 43090 42702 43102 42754
rect 39006 42690 39058 42702
rect 45278 42690 45330 42702
rect 9550 42642 9602 42654
rect 9550 42578 9602 42590
rect 12910 42642 12962 42654
rect 12910 42578 12962 42590
rect 14030 42642 14082 42654
rect 26126 42642 26178 42654
rect 16482 42590 16494 42642
rect 16546 42590 16558 42642
rect 14030 42578 14082 42590
rect 26126 42578 26178 42590
rect 29598 42642 29650 42654
rect 29598 42578 29650 42590
rect 33182 42642 33234 42654
rect 33182 42578 33234 42590
rect 33406 42642 33458 42654
rect 33406 42578 33458 42590
rect 34414 42642 34466 42654
rect 43710 42642 43762 42654
rect 34626 42590 34638 42642
rect 34690 42590 34702 42642
rect 34414 42578 34466 42590
rect 43710 42578 43762 42590
rect 44270 42642 44322 42654
rect 45390 42642 45442 42654
rect 44818 42590 44830 42642
rect 44882 42590 44894 42642
rect 44270 42578 44322 42590
rect 45390 42578 45442 42590
rect 45502 42642 45554 42654
rect 45502 42578 45554 42590
rect 46062 42642 46114 42654
rect 46062 42578 46114 42590
rect 12798 42530 12850 42542
rect 12798 42466 12850 42478
rect 26574 42530 26626 42542
rect 26574 42466 26626 42478
rect 27358 42530 27410 42542
rect 27358 42466 27410 42478
rect 27806 42530 27858 42542
rect 27806 42466 27858 42478
rect 28142 42530 28194 42542
rect 28142 42466 28194 42478
rect 28702 42530 28754 42542
rect 28702 42466 28754 42478
rect 30270 42530 30322 42542
rect 30270 42466 30322 42478
rect 31502 42530 31554 42542
rect 31502 42466 31554 42478
rect 31950 42530 32002 42542
rect 31950 42466 32002 42478
rect 34974 42530 35026 42542
rect 37214 42530 37266 42542
rect 36306 42478 36318 42530
rect 36370 42478 36382 42530
rect 34974 42466 35026 42478
rect 37214 42466 37266 42478
rect 37886 42530 37938 42542
rect 37886 42466 37938 42478
rect 43934 42530 43986 42542
rect 43934 42466 43986 42478
rect 44158 42530 44210 42542
rect 44158 42466 44210 42478
rect 45950 42530 46002 42542
rect 45950 42466 46002 42478
rect 1344 42362 46592 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 46592 42362
rect 1344 42276 46592 42310
rect 15822 42194 15874 42206
rect 15822 42130 15874 42142
rect 16382 42194 16434 42206
rect 31054 42194 31106 42206
rect 18834 42142 18846 42194
rect 18898 42142 18910 42194
rect 36642 42142 36654 42194
rect 36706 42142 36718 42194
rect 16382 42130 16434 42142
rect 31054 42130 31106 42142
rect 32174 42082 32226 42094
rect 17490 42030 17502 42082
rect 17554 42030 17566 42082
rect 32174 42018 32226 42030
rect 15486 41970 15538 41982
rect 5954 41918 5966 41970
rect 6018 41918 6030 41970
rect 6626 41918 6638 41970
rect 6690 41918 6702 41970
rect 13682 41918 13694 41970
rect 13746 41918 13758 41970
rect 15486 41906 15538 41918
rect 15710 41970 15762 41982
rect 15710 41906 15762 41918
rect 15934 41970 15986 41982
rect 15934 41906 15986 41918
rect 16494 41970 16546 41982
rect 31166 41970 31218 41982
rect 18050 41918 18062 41970
rect 18114 41918 18126 41970
rect 18386 41918 18398 41970
rect 18450 41918 18462 41970
rect 19394 41918 19406 41970
rect 19458 41918 19470 41970
rect 30146 41918 30158 41970
rect 30210 41918 30222 41970
rect 30930 41918 30942 41970
rect 30994 41918 31006 41970
rect 16494 41906 16546 41918
rect 31166 41906 31218 41918
rect 31838 41970 31890 41982
rect 36318 41970 36370 41982
rect 35970 41918 35982 41970
rect 36034 41918 36046 41970
rect 31838 41906 31890 41918
rect 36318 41906 36370 41918
rect 37102 41970 37154 41982
rect 37426 41918 37438 41970
rect 37490 41918 37502 41970
rect 44706 41918 44718 41970
rect 44770 41918 44782 41970
rect 37102 41906 37154 41918
rect 36990 41858 37042 41870
rect 8754 41806 8766 41858
rect 8818 41806 8830 41858
rect 10098 41806 10110 41858
rect 10162 41806 10174 41858
rect 18162 41806 18174 41858
rect 18226 41806 18238 41858
rect 21970 41806 21982 41858
rect 22034 41806 22046 41858
rect 28018 41806 28030 41858
rect 28082 41806 28094 41858
rect 33058 41806 33070 41858
rect 33122 41806 33134 41858
rect 35186 41806 35198 41858
rect 35250 41806 35262 41858
rect 38210 41806 38222 41858
rect 38274 41806 38286 41858
rect 40338 41806 40350 41858
rect 40402 41806 40414 41858
rect 42690 41806 42702 41858
rect 42754 41806 42766 41858
rect 36990 41794 37042 41806
rect 16382 41746 16434 41758
rect 16382 41682 16434 41694
rect 16718 41746 16770 41758
rect 16718 41682 16770 41694
rect 31390 41746 31442 41758
rect 31390 41682 31442 41694
rect 1344 41578 46592 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 46592 41578
rect 1344 41492 46592 41526
rect 9326 41410 9378 41422
rect 33182 41410 33234 41422
rect 9650 41358 9662 41410
rect 9714 41358 9726 41410
rect 30818 41358 30830 41410
rect 30882 41358 30894 41410
rect 9326 41346 9378 41358
rect 33182 41346 33234 41358
rect 33294 41410 33346 41422
rect 33294 41346 33346 41358
rect 33630 41410 33682 41422
rect 33630 41346 33682 41358
rect 35310 41410 35362 41422
rect 36094 41410 36146 41422
rect 35634 41358 35646 41410
rect 35698 41358 35710 41410
rect 35310 41346 35362 41358
rect 36094 41346 36146 41358
rect 45166 41410 45218 41422
rect 45166 41346 45218 41358
rect 15262 41298 15314 41310
rect 12898 41246 12910 41298
rect 12962 41246 12974 41298
rect 14914 41246 14926 41298
rect 14978 41246 14990 41298
rect 15262 41234 15314 41246
rect 16270 41298 16322 41310
rect 24670 41298 24722 41310
rect 30270 41298 30322 41310
rect 21298 41246 21310 41298
rect 21362 41246 21374 41298
rect 28130 41246 28142 41298
rect 28194 41246 28206 41298
rect 16270 41234 16322 41246
rect 24670 41234 24722 41246
rect 30270 41234 30322 41246
rect 32398 41298 32450 41310
rect 32398 41234 32450 41246
rect 35086 41298 35138 41310
rect 43934 41298 43986 41310
rect 37202 41246 37214 41298
rect 37266 41246 37278 41298
rect 35086 41234 35138 41246
rect 43934 41234 43986 41246
rect 45838 41298 45890 41310
rect 45838 41234 45890 41246
rect 9102 41186 9154 41198
rect 18062 41186 18114 41198
rect 30046 41186 30098 41198
rect 10098 41134 10110 41186
rect 10162 41134 10174 41186
rect 14690 41134 14702 41186
rect 14754 41134 14766 41186
rect 15586 41134 15598 41186
rect 15650 41134 15662 41186
rect 17266 41134 17278 41186
rect 17330 41134 17342 41186
rect 18386 41134 18398 41186
rect 18450 41134 18462 41186
rect 20402 41134 20414 41186
rect 20466 41134 20478 41186
rect 24210 41134 24222 41186
rect 24274 41134 24286 41186
rect 25330 41134 25342 41186
rect 25394 41134 25406 41186
rect 9102 41122 9154 41134
rect 18062 41122 18114 41134
rect 30046 41122 30098 41134
rect 30494 41186 30546 41198
rect 30494 41122 30546 41134
rect 33518 41186 33570 41198
rect 42590 41186 42642 41198
rect 36418 41134 36430 41186
rect 36482 41134 36494 41186
rect 41906 41134 41918 41186
rect 41970 41134 41982 41186
rect 33518 41122 33570 41134
rect 42590 41122 42642 41134
rect 43486 41186 43538 41198
rect 43486 41122 43538 41134
rect 43710 41186 43762 41198
rect 43710 41122 43762 41134
rect 44830 41186 44882 41198
rect 44830 41122 44882 41134
rect 44942 41186 44994 41198
rect 44942 41122 44994 41134
rect 45278 41186 45330 41198
rect 45278 41122 45330 41134
rect 14030 41074 14082 41086
rect 28590 41074 28642 41086
rect 10770 41022 10782 41074
rect 10834 41022 10846 41074
rect 15810 41022 15822 41074
rect 15874 41022 15886 41074
rect 16146 41022 16158 41074
rect 16210 41022 16222 41074
rect 20626 41022 20638 41074
rect 20690 41022 20702 41074
rect 23426 41022 23438 41074
rect 23490 41022 23502 41074
rect 26002 41022 26014 41074
rect 26066 41022 26078 41074
rect 14030 41010 14082 41022
rect 28590 41010 28642 41022
rect 31166 41074 31218 41086
rect 31166 41010 31218 41022
rect 31950 41074 32002 41086
rect 31950 41010 32002 41022
rect 44046 41074 44098 41086
rect 44046 41010 44098 41022
rect 45726 41074 45778 41086
rect 45726 41010 45778 41022
rect 13694 40962 13746 40974
rect 13694 40898 13746 40910
rect 20862 40962 20914 40974
rect 20862 40898 20914 40910
rect 24558 40962 24610 40974
rect 24558 40898 24610 40910
rect 28478 40962 28530 40974
rect 28478 40898 28530 40910
rect 29374 40962 29426 40974
rect 29374 40898 29426 40910
rect 29486 40962 29538 40974
rect 29486 40898 29538 40910
rect 29598 40962 29650 40974
rect 29598 40898 29650 40910
rect 31278 40962 31330 40974
rect 31278 40898 31330 40910
rect 31390 40962 31442 40974
rect 31390 40898 31442 40910
rect 31838 40962 31890 40974
rect 31838 40898 31890 40910
rect 32286 40962 32338 40974
rect 32286 40898 32338 40910
rect 32846 40962 32898 40974
rect 32846 40898 32898 40910
rect 34190 40962 34242 40974
rect 34190 40898 34242 40910
rect 34750 40962 34802 40974
rect 34750 40898 34802 40910
rect 36206 40962 36258 40974
rect 36206 40898 36258 40910
rect 43150 40962 43202 40974
rect 43150 40898 43202 40910
rect 45950 40962 46002 40974
rect 45950 40898 46002 40910
rect 1344 40794 46592 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 46592 40794
rect 1344 40708 46592 40742
rect 16718 40626 16770 40638
rect 24446 40626 24498 40638
rect 16258 40574 16270 40626
rect 16322 40574 16334 40626
rect 22194 40574 22206 40626
rect 22258 40574 22270 40626
rect 23538 40574 23550 40626
rect 23602 40574 23614 40626
rect 16718 40562 16770 40574
rect 24446 40562 24498 40574
rect 28590 40626 28642 40638
rect 28590 40562 28642 40574
rect 30606 40626 30658 40638
rect 30606 40562 30658 40574
rect 32174 40626 32226 40638
rect 32174 40562 32226 40574
rect 33182 40626 33234 40638
rect 33182 40562 33234 40574
rect 33854 40626 33906 40638
rect 33854 40562 33906 40574
rect 35198 40626 35250 40638
rect 35198 40562 35250 40574
rect 36766 40626 36818 40638
rect 36766 40562 36818 40574
rect 40350 40626 40402 40638
rect 40350 40562 40402 40574
rect 45614 40626 45666 40638
rect 45614 40562 45666 40574
rect 11230 40514 11282 40526
rect 11230 40450 11282 40462
rect 15038 40514 15090 40526
rect 15038 40450 15090 40462
rect 15710 40514 15762 40526
rect 15710 40450 15762 40462
rect 15822 40514 15874 40526
rect 15822 40450 15874 40462
rect 17502 40514 17554 40526
rect 29374 40514 29426 40526
rect 18946 40462 18958 40514
rect 19010 40462 19022 40514
rect 21634 40462 21646 40514
rect 21698 40462 21710 40514
rect 22866 40462 22878 40514
rect 22930 40462 22942 40514
rect 23202 40462 23214 40514
rect 23266 40462 23278 40514
rect 17502 40450 17554 40462
rect 29374 40450 29426 40462
rect 30494 40514 30546 40526
rect 30494 40450 30546 40462
rect 30718 40514 30770 40526
rect 30718 40450 30770 40462
rect 35086 40514 35138 40526
rect 35086 40450 35138 40462
rect 35534 40514 35586 40526
rect 45838 40514 45890 40526
rect 35858 40462 35870 40514
rect 35922 40462 35934 40514
rect 41682 40462 41694 40514
rect 41746 40462 41758 40514
rect 35534 40450 35586 40462
rect 45838 40450 45890 40462
rect 9774 40402 9826 40414
rect 16830 40402 16882 40414
rect 30382 40402 30434 40414
rect 31278 40402 31330 40414
rect 6066 40350 6078 40402
rect 6130 40350 6142 40402
rect 10098 40350 10110 40402
rect 10162 40350 10174 40402
rect 11778 40350 11790 40402
rect 11842 40350 11854 40402
rect 15474 40350 15486 40402
rect 15538 40350 15550 40402
rect 18722 40350 18734 40402
rect 18786 40350 18798 40402
rect 20178 40350 20190 40402
rect 20242 40350 20254 40402
rect 21858 40350 21870 40402
rect 21922 40350 21934 40402
rect 23650 40350 23662 40402
rect 23714 40350 23726 40402
rect 24098 40350 24110 40402
rect 24162 40350 24174 40402
rect 27346 40350 27358 40402
rect 27410 40350 27422 40402
rect 28018 40350 28030 40402
rect 28082 40350 28094 40402
rect 30930 40350 30942 40402
rect 30994 40350 31006 40402
rect 9774 40338 9826 40350
rect 16830 40338 16882 40350
rect 30382 40338 30434 40350
rect 31278 40338 31330 40350
rect 31838 40402 31890 40414
rect 31838 40338 31890 40350
rect 31950 40402 32002 40414
rect 33406 40402 33458 40414
rect 32386 40350 32398 40402
rect 32450 40350 32462 40402
rect 31950 40338 32002 40350
rect 33406 40338 33458 40350
rect 34302 40402 34354 40414
rect 39118 40402 39170 40414
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 38882 40350 38894 40402
rect 38946 40350 38958 40402
rect 34302 40338 34354 40350
rect 39118 40338 39170 40350
rect 39342 40402 39394 40414
rect 39342 40338 39394 40350
rect 39454 40402 39506 40414
rect 45054 40402 45106 40414
rect 40114 40350 40126 40402
rect 40178 40350 40190 40402
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 44706 40350 44718 40402
rect 44770 40350 44782 40402
rect 39454 40338 39506 40350
rect 45054 40338 45106 40350
rect 45166 40402 45218 40414
rect 45166 40338 45218 40350
rect 45390 40402 45442 40414
rect 45390 40338 45442 40350
rect 45950 40402 46002 40414
rect 45950 40338 46002 40350
rect 10670 40290 10722 40302
rect 11454 40290 11506 40302
rect 17614 40290 17666 40302
rect 6850 40238 6862 40290
rect 6914 40238 6926 40290
rect 8978 40238 8990 40290
rect 9042 40238 9054 40290
rect 11106 40238 11118 40290
rect 11170 40238 11182 40290
rect 12562 40238 12574 40290
rect 12626 40238 12638 40290
rect 14690 40238 14702 40290
rect 14754 40238 14766 40290
rect 10670 40226 10722 40238
rect 11454 40226 11506 40238
rect 17614 40226 17666 40238
rect 22542 40290 22594 40302
rect 29710 40290 29762 40302
rect 25218 40238 25230 40290
rect 25282 40238 25294 40290
rect 22542 40226 22594 40238
rect 29710 40226 29762 40238
rect 29822 40290 29874 40302
rect 29822 40226 29874 40238
rect 31390 40290 31442 40302
rect 34862 40290 34914 40302
rect 32274 40238 32286 40290
rect 32338 40238 32350 40290
rect 31390 40226 31442 40238
rect 34862 40226 34914 40238
rect 36878 40290 36930 40302
rect 36878 40226 36930 40238
rect 37214 40290 37266 40302
rect 38098 40238 38110 40290
rect 38162 40238 38174 40290
rect 43810 40238 43822 40290
rect 43874 40238 43886 40290
rect 37214 40226 37266 40238
rect 15150 40178 15202 40190
rect 15150 40114 15202 40126
rect 16718 40178 16770 40190
rect 16718 40114 16770 40126
rect 17726 40178 17778 40190
rect 17726 40114 17778 40126
rect 28590 40178 28642 40190
rect 28590 40114 28642 40126
rect 28702 40178 28754 40190
rect 28702 40114 28754 40126
rect 28926 40178 28978 40190
rect 28926 40114 28978 40126
rect 29486 40178 29538 40190
rect 29486 40114 29538 40126
rect 33070 40178 33122 40190
rect 39006 40178 39058 40190
rect 33618 40126 33630 40178
rect 33682 40175 33694 40178
rect 34178 40175 34190 40178
rect 33682 40129 34190 40175
rect 33682 40126 33694 40129
rect 34178 40126 34190 40129
rect 34242 40126 34254 40178
rect 33070 40114 33122 40126
rect 39006 40114 39058 40126
rect 1344 40010 46592 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 46592 40010
rect 1344 39924 46592 39958
rect 10222 39842 10274 39854
rect 10222 39778 10274 39790
rect 10558 39842 10610 39854
rect 10558 39778 10610 39790
rect 11006 39842 11058 39854
rect 11006 39778 11058 39790
rect 11790 39842 11842 39854
rect 11790 39778 11842 39790
rect 13470 39842 13522 39854
rect 21422 39842 21474 39854
rect 18274 39790 18286 39842
rect 18338 39790 18350 39842
rect 13470 39778 13522 39790
rect 21422 39778 21474 39790
rect 30270 39842 30322 39854
rect 30270 39778 30322 39790
rect 31166 39842 31218 39854
rect 31166 39778 31218 39790
rect 34078 39842 34130 39854
rect 34078 39778 34130 39790
rect 36990 39842 37042 39854
rect 36990 39778 37042 39790
rect 37326 39842 37378 39854
rect 37326 39778 37378 39790
rect 11118 39730 11170 39742
rect 29710 39730 29762 39742
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 15698 39678 15710 39730
rect 15762 39678 15774 39730
rect 17266 39678 17278 39730
rect 17330 39678 17342 39730
rect 18386 39678 18398 39730
rect 18450 39678 18462 39730
rect 24658 39678 24670 39730
rect 24722 39678 24734 39730
rect 24994 39678 25006 39730
rect 25058 39678 25070 39730
rect 27122 39678 27134 39730
rect 27186 39678 27198 39730
rect 11118 39666 11170 39678
rect 29710 39666 29762 39678
rect 32958 39730 33010 39742
rect 32958 39666 33010 39678
rect 34190 39730 34242 39742
rect 34190 39666 34242 39678
rect 37774 39730 37826 39742
rect 41906 39678 41918 39730
rect 41970 39678 41982 39730
rect 37774 39666 37826 39678
rect 8094 39618 8146 39630
rect 9662 39618 9714 39630
rect 12910 39618 12962 39630
rect 14142 39618 14194 39630
rect 19070 39618 19122 39630
rect 28254 39618 28306 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 8306 39566 8318 39618
rect 8370 39566 8382 39618
rect 11890 39566 11902 39618
rect 11954 39566 11966 39618
rect 13458 39566 13470 39618
rect 13522 39566 13534 39618
rect 15474 39566 15486 39618
rect 15538 39566 15550 39618
rect 17154 39566 17166 39618
rect 17218 39566 17230 39618
rect 18162 39566 18174 39618
rect 18226 39566 18238 39618
rect 19282 39566 19294 39618
rect 19346 39566 19358 39618
rect 20066 39566 20078 39618
rect 20130 39566 20142 39618
rect 20514 39566 20526 39618
rect 20578 39566 20590 39618
rect 21858 39566 21870 39618
rect 21922 39566 21934 39618
rect 27906 39566 27918 39618
rect 27970 39566 27982 39618
rect 8094 39554 8146 39566
rect 9662 39554 9714 39566
rect 12910 39554 12962 39566
rect 14142 39554 14194 39566
rect 19070 39554 19122 39566
rect 28254 39554 28306 39566
rect 29822 39618 29874 39630
rect 31166 39618 31218 39630
rect 29922 39566 29934 39618
rect 29986 39566 29998 39618
rect 29822 39554 29874 39566
rect 31166 39554 31218 39566
rect 31614 39618 31666 39630
rect 32734 39618 32786 39630
rect 32498 39566 32510 39618
rect 32562 39566 32574 39618
rect 31614 39554 31666 39566
rect 32734 39554 32786 39566
rect 33070 39618 33122 39630
rect 33070 39554 33122 39566
rect 33518 39618 33570 39630
rect 33518 39554 33570 39566
rect 34974 39618 35026 39630
rect 34974 39554 35026 39566
rect 35758 39618 35810 39630
rect 44830 39618 44882 39630
rect 38658 39566 38670 39618
rect 38722 39566 38734 39618
rect 40674 39566 40686 39618
rect 40738 39566 40750 39618
rect 43026 39566 43038 39618
rect 43090 39566 43102 39618
rect 43362 39566 43374 39618
rect 43426 39566 43438 39618
rect 44258 39566 44270 39618
rect 44322 39566 44334 39618
rect 35758 39554 35810 39566
rect 44830 39554 44882 39566
rect 45614 39618 45666 39630
rect 45614 39554 45666 39566
rect 7758 39506 7810 39518
rect 2482 39454 2494 39506
rect 2546 39454 2558 39506
rect 7758 39442 7810 39454
rect 10334 39506 10386 39518
rect 10334 39442 10386 39454
rect 11230 39506 11282 39518
rect 11230 39442 11282 39454
rect 13806 39506 13858 39518
rect 13806 39442 13858 39454
rect 14814 39506 14866 39518
rect 21310 39506 21362 39518
rect 30606 39506 30658 39518
rect 16146 39454 16158 39506
rect 16210 39454 16222 39506
rect 19618 39454 19630 39506
rect 19682 39454 19694 39506
rect 22530 39454 22542 39506
rect 22594 39454 22606 39506
rect 14814 39442 14866 39454
rect 21310 39442 21362 39454
rect 30606 39442 30658 39454
rect 31726 39506 31778 39518
rect 31726 39442 31778 39454
rect 32286 39506 32338 39518
rect 32286 39442 32338 39454
rect 33182 39506 33234 39518
rect 33182 39442 33234 39454
rect 33630 39506 33682 39518
rect 33630 39442 33682 39454
rect 35198 39506 35250 39518
rect 35198 39442 35250 39454
rect 35534 39506 35586 39518
rect 41246 39506 41298 39518
rect 44046 39506 44098 39518
rect 38770 39454 38782 39506
rect 38834 39454 38846 39506
rect 42802 39454 42814 39506
rect 42866 39454 42878 39506
rect 35534 39442 35586 39454
rect 41246 39442 41298 39454
rect 44046 39442 44098 39454
rect 7086 39394 7138 39406
rect 7086 39330 7138 39342
rect 7422 39394 7474 39406
rect 7422 39330 7474 39342
rect 7870 39394 7922 39406
rect 7870 39330 7922 39342
rect 8654 39394 8706 39406
rect 8654 39330 8706 39342
rect 8766 39394 8818 39406
rect 8766 39330 8818 39342
rect 8878 39394 8930 39406
rect 8878 39330 8930 39342
rect 9438 39394 9490 39406
rect 9438 39330 9490 39342
rect 9774 39394 9826 39406
rect 9774 39330 9826 39342
rect 9998 39394 10050 39406
rect 9998 39330 10050 39342
rect 12574 39394 12626 39406
rect 16494 39394 16546 39406
rect 29598 39394 29650 39406
rect 14466 39342 14478 39394
rect 14530 39342 14542 39394
rect 28578 39342 28590 39394
rect 28642 39342 28654 39394
rect 12574 39330 12626 39342
rect 16494 39330 16546 39342
rect 29598 39330 29650 39342
rect 30830 39394 30882 39406
rect 30830 39330 30882 39342
rect 31054 39394 31106 39406
rect 31054 39330 31106 39342
rect 31950 39394 32002 39406
rect 31950 39330 32002 39342
rect 33854 39394 33906 39406
rect 37102 39394 37154 39406
rect 34626 39342 34638 39394
rect 34690 39342 34702 39394
rect 36082 39342 36094 39394
rect 36146 39342 36158 39394
rect 33854 39330 33906 39342
rect 37102 39330 37154 39342
rect 38334 39394 38386 39406
rect 46174 39394 46226 39406
rect 45154 39342 45166 39394
rect 45218 39342 45230 39394
rect 38334 39330 38386 39342
rect 46174 39330 46226 39342
rect 1344 39226 46592 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 46592 39226
rect 1344 39140 46592 39174
rect 13134 39058 13186 39070
rect 23102 39058 23154 39070
rect 14130 39006 14142 39058
rect 14194 39006 14206 39058
rect 17378 39006 17390 39058
rect 17442 39006 17454 39058
rect 13134 38994 13186 39006
rect 23102 38994 23154 39006
rect 23214 39058 23266 39070
rect 23214 38994 23266 39006
rect 23438 39058 23490 39070
rect 23438 38994 23490 39006
rect 24334 39058 24386 39070
rect 24334 38994 24386 39006
rect 26686 39058 26738 39070
rect 26686 38994 26738 39006
rect 27358 39058 27410 39070
rect 27358 38994 27410 39006
rect 27470 39058 27522 39070
rect 27470 38994 27522 39006
rect 27582 39058 27634 39070
rect 27582 38994 27634 39006
rect 29822 39058 29874 39070
rect 29822 38994 29874 39006
rect 32174 39058 32226 39070
rect 32174 38994 32226 39006
rect 33070 39058 33122 39070
rect 33070 38994 33122 39006
rect 33630 39058 33682 39070
rect 33630 38994 33682 39006
rect 35086 39058 35138 39070
rect 35086 38994 35138 39006
rect 40014 39058 40066 39070
rect 40014 38994 40066 39006
rect 41022 39058 41074 39070
rect 45042 39006 45054 39058
rect 45106 39006 45118 39058
rect 41022 38994 41074 39006
rect 2830 38946 2882 38958
rect 2830 38882 2882 38894
rect 3502 38946 3554 38958
rect 3502 38882 3554 38894
rect 4174 38946 4226 38958
rect 8990 38946 9042 38958
rect 6066 38894 6078 38946
rect 6130 38894 6142 38946
rect 4174 38882 4226 38894
rect 8990 38882 9042 38894
rect 13806 38946 13858 38958
rect 13806 38882 13858 38894
rect 16606 38946 16658 38958
rect 16606 38882 16658 38894
rect 22878 38946 22930 38958
rect 22878 38882 22930 38894
rect 23326 38946 23378 38958
rect 23326 38882 23378 38894
rect 24110 38946 24162 38958
rect 24110 38882 24162 38894
rect 24670 38946 24722 38958
rect 24670 38882 24722 38894
rect 28030 38946 28082 38958
rect 28030 38882 28082 38894
rect 29374 38946 29426 38958
rect 29374 38882 29426 38894
rect 31726 38946 31778 38958
rect 31726 38882 31778 38894
rect 34302 38946 34354 38958
rect 40238 38946 40290 38958
rect 36530 38894 36542 38946
rect 36594 38894 36606 38946
rect 34302 38882 34354 38894
rect 40238 38882 40290 38894
rect 40350 38946 40402 38958
rect 45950 38946 46002 38958
rect 43474 38894 43486 38946
rect 43538 38894 43550 38946
rect 44930 38894 44942 38946
rect 44994 38894 45006 38946
rect 40350 38882 40402 38894
rect 45950 38882 46002 38894
rect 3950 38834 4002 38846
rect 3714 38782 3726 38834
rect 3778 38782 3790 38834
rect 3950 38770 4002 38782
rect 4286 38834 4338 38846
rect 8654 38834 8706 38846
rect 13022 38834 13074 38846
rect 5282 38782 5294 38834
rect 5346 38782 5358 38834
rect 9874 38782 9886 38834
rect 9938 38782 9950 38834
rect 4286 38770 4338 38782
rect 8654 38770 8706 38782
rect 13022 38770 13074 38782
rect 13470 38834 13522 38846
rect 13470 38770 13522 38782
rect 14478 38834 14530 38846
rect 16046 38834 16098 38846
rect 15698 38782 15710 38834
rect 15762 38782 15774 38834
rect 14478 38770 14530 38782
rect 16046 38770 16098 38782
rect 17726 38834 17778 38846
rect 24446 38834 24498 38846
rect 27246 38834 27298 38846
rect 19170 38782 19182 38834
rect 19234 38782 19246 38834
rect 20178 38782 20190 38834
rect 20242 38782 20254 38834
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 21298 38782 21310 38834
rect 21362 38782 21374 38834
rect 25890 38782 25902 38834
rect 25954 38782 25966 38834
rect 27010 38782 27022 38834
rect 27074 38782 27086 38834
rect 17726 38770 17778 38782
rect 24446 38770 24498 38782
rect 27246 38770 27298 38782
rect 28366 38834 28418 38846
rect 28926 38834 28978 38846
rect 28690 38782 28702 38834
rect 28754 38782 28766 38834
rect 28366 38770 28418 38782
rect 28926 38770 28978 38782
rect 29262 38834 29314 38846
rect 29262 38770 29314 38782
rect 30494 38834 30546 38846
rect 30494 38770 30546 38782
rect 30718 38834 30770 38846
rect 30718 38770 30770 38782
rect 30942 38834 30994 38846
rect 30942 38770 30994 38782
rect 33854 38834 33906 38846
rect 33854 38770 33906 38782
rect 34414 38834 34466 38846
rect 34414 38770 34466 38782
rect 34638 38834 34690 38846
rect 34638 38770 34690 38782
rect 34974 38834 35026 38846
rect 39118 38834 39170 38846
rect 35746 38782 35758 38834
rect 35810 38782 35822 38834
rect 34974 38770 35026 38782
rect 39118 38770 39170 38782
rect 39342 38834 39394 38846
rect 39342 38770 39394 38782
rect 40910 38834 40962 38846
rect 44146 38782 44158 38834
rect 44210 38782 44222 38834
rect 45154 38782 45166 38834
rect 45218 38782 45230 38834
rect 45602 38782 45614 38834
rect 45666 38782 45678 38834
rect 40910 38770 40962 38782
rect 3054 38722 3106 38734
rect 15150 38722 15202 38734
rect 2706 38670 2718 38722
rect 2770 38670 2782 38722
rect 8194 38670 8206 38722
rect 8258 38670 8270 38722
rect 10546 38670 10558 38722
rect 10610 38670 10622 38722
rect 12674 38670 12686 38722
rect 12738 38670 12750 38722
rect 3054 38658 3106 38670
rect 15150 38658 15202 38670
rect 15262 38722 15314 38734
rect 15262 38658 15314 38670
rect 15486 38722 15538 38734
rect 16830 38722 16882 38734
rect 25230 38722 25282 38734
rect 29150 38722 29202 38734
rect 16482 38670 16494 38722
rect 16546 38670 16558 38722
rect 18722 38670 18734 38722
rect 18786 38670 18798 38722
rect 20626 38670 20638 38722
rect 20690 38670 20702 38722
rect 26114 38670 26126 38722
rect 26178 38670 26190 38722
rect 15486 38658 15538 38670
rect 16830 38658 16882 38670
rect 25230 38658 25282 38670
rect 29150 38658 29202 38670
rect 33182 38722 33234 38734
rect 39230 38722 39282 38734
rect 38658 38670 38670 38722
rect 38722 38670 38734 38722
rect 33182 38658 33234 38670
rect 39230 38658 39282 38670
rect 39566 38722 39618 38734
rect 39566 38658 39618 38670
rect 39790 38722 39842 38734
rect 41346 38670 41358 38722
rect 41410 38670 41422 38722
rect 39790 38658 39842 38670
rect 3390 38610 3442 38622
rect 3390 38546 3442 38558
rect 16158 38610 16210 38622
rect 16158 38546 16210 38558
rect 28142 38610 28194 38622
rect 28142 38546 28194 38558
rect 31390 38610 31442 38622
rect 31390 38546 31442 38558
rect 1344 38442 46592 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 46592 38442
rect 1344 38356 46592 38390
rect 4398 38274 4450 38286
rect 27246 38274 27298 38286
rect 21746 38222 21758 38274
rect 21810 38222 21822 38274
rect 4398 38210 4450 38222
rect 27246 38210 27298 38222
rect 32510 38274 32562 38286
rect 32510 38210 32562 38222
rect 35198 38274 35250 38286
rect 35198 38210 35250 38222
rect 11342 38162 11394 38174
rect 25118 38162 25170 38174
rect 27358 38162 27410 38174
rect 3602 38110 3614 38162
rect 3666 38110 3678 38162
rect 20066 38110 20078 38162
rect 20130 38110 20142 38162
rect 25442 38110 25454 38162
rect 25506 38110 25518 38162
rect 11342 38098 11394 38110
rect 25118 38098 25170 38110
rect 27358 38098 27410 38110
rect 29486 38162 29538 38174
rect 43374 38162 43426 38174
rect 45950 38162 46002 38174
rect 34514 38110 34526 38162
rect 34578 38110 34590 38162
rect 39778 38110 39790 38162
rect 39842 38110 39854 38162
rect 41906 38110 41918 38162
rect 41970 38110 41982 38162
rect 44930 38110 44942 38162
rect 44994 38110 45006 38162
rect 29486 38098 29538 38110
rect 43374 38098 43426 38110
rect 45950 38098 46002 38110
rect 4286 38050 4338 38062
rect 11118 38050 11170 38062
rect 3378 37998 3390 38050
rect 3442 37998 3454 38050
rect 10098 37998 10110 38050
rect 10162 37998 10174 38050
rect 4286 37986 4338 37998
rect 11118 37986 11170 37998
rect 11566 38050 11618 38062
rect 11566 37986 11618 37998
rect 11790 38050 11842 38062
rect 27694 38050 27746 38062
rect 29374 38050 29426 38062
rect 18050 37998 18062 38050
rect 18114 37998 18126 38050
rect 19058 37998 19070 38050
rect 19122 37998 19134 38050
rect 20290 37998 20302 38050
rect 20354 37998 20366 38050
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 22530 37998 22542 38050
rect 22594 37998 22606 38050
rect 24434 37998 24446 38050
rect 24498 37998 24510 38050
rect 25778 37998 25790 38050
rect 25842 37998 25854 38050
rect 26674 37998 26686 38050
rect 26738 37998 26750 38050
rect 28018 37998 28030 38050
rect 28082 37998 28094 38050
rect 11790 37986 11842 37998
rect 27694 37986 27746 37998
rect 29374 37986 29426 37998
rect 29598 38050 29650 38062
rect 30158 38050 30210 38062
rect 29810 37998 29822 38050
rect 29874 37998 29886 38050
rect 29598 37986 29650 37998
rect 30158 37986 30210 37998
rect 30494 38050 30546 38062
rect 30494 37986 30546 37998
rect 30718 38050 30770 38062
rect 30718 37986 30770 37998
rect 31054 38050 31106 38062
rect 34414 38050 34466 38062
rect 31378 37998 31390 38050
rect 31442 37998 31454 38050
rect 31826 37998 31838 38050
rect 31890 37998 31902 38050
rect 32722 37998 32734 38050
rect 32786 37998 32798 38050
rect 31054 37986 31106 37998
rect 34414 37986 34466 37998
rect 34974 38050 35026 38062
rect 34974 37986 35026 37998
rect 35982 38050 36034 38062
rect 35982 37986 36034 37998
rect 36094 38050 36146 38062
rect 39342 38050 39394 38062
rect 43486 38050 43538 38062
rect 45054 38050 45106 38062
rect 37874 37998 37886 38050
rect 37938 37998 37950 38050
rect 38322 37998 38334 38050
rect 38386 37998 38398 38050
rect 38882 37998 38894 38050
rect 38946 37998 38958 38050
rect 42690 37998 42702 38050
rect 42754 37998 42766 38050
rect 43026 37998 43038 38050
rect 43090 37998 43102 38050
rect 43698 37998 43710 38050
rect 43762 37998 43774 38050
rect 36094 37986 36146 37998
rect 39342 37986 39394 37998
rect 43486 37986 43538 37998
rect 45054 37986 45106 37998
rect 45278 38050 45330 38062
rect 45278 37986 45330 37998
rect 45390 38050 45442 38062
rect 45390 37986 45442 37998
rect 3950 37938 4002 37950
rect 12574 37938 12626 37950
rect 5842 37886 5854 37938
rect 5906 37886 5918 37938
rect 3950 37874 4002 37886
rect 12574 37874 12626 37886
rect 12798 37938 12850 37950
rect 28254 37938 28306 37950
rect 13682 37886 13694 37938
rect 13746 37886 13758 37938
rect 20402 37886 20414 37938
rect 20466 37886 20478 37938
rect 23874 37886 23886 37938
rect 23938 37886 23950 37938
rect 26786 37886 26798 37938
rect 26850 37886 26862 37938
rect 12798 37874 12850 37886
rect 28254 37874 28306 37886
rect 29150 37938 29202 37950
rect 29150 37874 29202 37886
rect 33966 37938 34018 37950
rect 35870 37938 35922 37950
rect 35522 37886 35534 37938
rect 35586 37886 35598 37938
rect 33966 37874 34018 37886
rect 35870 37874 35922 37886
rect 36430 37938 36482 37950
rect 36430 37874 36482 37886
rect 37326 37938 37378 37950
rect 44046 37938 44098 37950
rect 38546 37886 38558 37938
rect 38610 37886 38622 37938
rect 37326 37874 37378 37886
rect 44046 37874 44098 37886
rect 44158 37938 44210 37950
rect 44158 37874 44210 37886
rect 45838 37938 45890 37950
rect 45838 37874 45890 37886
rect 46062 37938 46114 37950
rect 46062 37874 46114 37886
rect 4398 37826 4450 37838
rect 4398 37762 4450 37774
rect 12350 37826 12402 37838
rect 12350 37762 12402 37774
rect 12686 37826 12738 37838
rect 12686 37762 12738 37774
rect 19294 37826 19346 37838
rect 28142 37826 28194 37838
rect 26002 37774 26014 37826
rect 26066 37774 26078 37826
rect 19294 37762 19346 37774
rect 28142 37762 28194 37774
rect 28366 37826 28418 37838
rect 28366 37762 28418 37774
rect 30270 37826 30322 37838
rect 30270 37762 30322 37774
rect 30830 37826 30882 37838
rect 30830 37762 30882 37774
rect 33182 37826 33234 37838
rect 33182 37762 33234 37774
rect 33518 37826 33570 37838
rect 33518 37762 33570 37774
rect 34190 37826 34242 37838
rect 34190 37762 34242 37774
rect 34526 37826 34578 37838
rect 34526 37762 34578 37774
rect 37214 37826 37266 37838
rect 37214 37762 37266 37774
rect 43262 37826 43314 37838
rect 43262 37762 43314 37774
rect 44382 37826 44434 37838
rect 44382 37762 44434 37774
rect 44942 37826 44994 37838
rect 44942 37762 44994 37774
rect 1344 37658 46592 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 46592 37658
rect 1344 37572 46592 37606
rect 5070 37490 5122 37502
rect 5070 37426 5122 37438
rect 5182 37490 5234 37502
rect 5182 37426 5234 37438
rect 8990 37490 9042 37502
rect 17502 37490 17554 37502
rect 30830 37490 30882 37502
rect 12898 37438 12910 37490
rect 12962 37438 12974 37490
rect 22866 37438 22878 37490
rect 22930 37438 22942 37490
rect 23650 37438 23662 37490
rect 23714 37438 23726 37490
rect 27794 37438 27806 37490
rect 27858 37438 27870 37490
rect 8990 37426 9042 37438
rect 17502 37426 17554 37438
rect 30830 37426 30882 37438
rect 31390 37490 31442 37502
rect 31390 37426 31442 37438
rect 38894 37490 38946 37502
rect 38894 37426 38946 37438
rect 8878 37378 8930 37390
rect 24110 37378 24162 37390
rect 6402 37326 6414 37378
rect 6466 37326 6478 37378
rect 9538 37326 9550 37378
rect 9602 37326 9614 37378
rect 10434 37326 10446 37378
rect 10498 37326 10510 37378
rect 14242 37326 14254 37378
rect 14306 37326 14318 37378
rect 18386 37326 18398 37378
rect 18450 37326 18462 37378
rect 8878 37314 8930 37326
rect 24110 37314 24162 37326
rect 24222 37378 24274 37390
rect 24222 37314 24274 37326
rect 26686 37378 26738 37390
rect 29922 37326 29934 37378
rect 29986 37326 29998 37378
rect 39778 37326 39790 37378
rect 39842 37326 39854 37378
rect 26686 37314 26738 37326
rect 9886 37266 9938 37278
rect 4610 37214 4622 37266
rect 4674 37214 4686 37266
rect 5730 37214 5742 37266
rect 5794 37214 5806 37266
rect 9886 37202 9938 37214
rect 10782 37266 10834 37278
rect 10782 37202 10834 37214
rect 11790 37266 11842 37278
rect 11790 37202 11842 37214
rect 12574 37266 12626 37278
rect 16942 37266 16994 37278
rect 13458 37214 13470 37266
rect 13522 37214 13534 37266
rect 12574 37202 12626 37214
rect 16942 37202 16994 37214
rect 17726 37266 17778 37278
rect 17726 37202 17778 37214
rect 18174 37266 18226 37278
rect 23326 37266 23378 37278
rect 21970 37214 21982 37266
rect 22034 37214 22046 37266
rect 22642 37214 22654 37266
rect 22706 37214 22718 37266
rect 18174 37202 18226 37214
rect 23326 37202 23378 37214
rect 24670 37266 24722 37278
rect 31278 37266 31330 37278
rect 26114 37214 26126 37266
rect 26178 37214 26190 37266
rect 28130 37214 28142 37266
rect 28194 37214 28206 37266
rect 35298 37214 35310 37266
rect 35362 37214 35374 37266
rect 38994 37214 39006 37266
rect 39058 37214 39070 37266
rect 39554 37214 39566 37266
rect 39618 37214 39630 37266
rect 41794 37214 41806 37266
rect 41858 37214 41870 37266
rect 24670 37202 24722 37214
rect 31278 37202 31330 37214
rect 10110 37154 10162 37166
rect 1698 37102 1710 37154
rect 1762 37102 1774 37154
rect 3826 37102 3838 37154
rect 3890 37102 3902 37154
rect 8530 37102 8542 37154
rect 8594 37102 8606 37154
rect 10110 37090 10162 37102
rect 12014 37154 12066 37166
rect 12014 37090 12066 37102
rect 12350 37154 12402 37166
rect 18510 37154 18562 37166
rect 25454 37154 25506 37166
rect 16370 37102 16382 37154
rect 16434 37102 16446 37154
rect 19170 37102 19182 37154
rect 19234 37102 19246 37154
rect 21298 37102 21310 37154
rect 21362 37102 21374 37154
rect 12350 37090 12402 37102
rect 18510 37090 18562 37102
rect 25454 37090 25506 37102
rect 30270 37154 30322 37166
rect 30270 37090 30322 37102
rect 30382 37154 30434 37166
rect 30382 37090 30434 37102
rect 31838 37154 31890 37166
rect 31838 37090 31890 37102
rect 32398 37154 32450 37166
rect 32398 37090 32450 37102
rect 33294 37154 33346 37166
rect 33294 37090 33346 37102
rect 33742 37154 33794 37166
rect 33742 37090 33794 37102
rect 34078 37154 34130 37166
rect 34078 37090 34130 37102
rect 34526 37154 34578 37166
rect 35970 37102 35982 37154
rect 36034 37102 36046 37154
rect 38098 37102 38110 37154
rect 38162 37102 38174 37154
rect 39442 37102 39454 37154
rect 39506 37102 39518 37154
rect 43362 37102 43374 37154
rect 43426 37102 43438 37154
rect 34526 37090 34578 37102
rect 4958 37042 5010 37054
rect 4958 36978 5010 36990
rect 11454 37042 11506 37054
rect 11454 36978 11506 36990
rect 24110 37042 24162 37054
rect 24110 36978 24162 36990
rect 31726 37042 31778 37054
rect 31726 36978 31778 36990
rect 32510 37042 32562 37054
rect 32510 36978 32562 36990
rect 33966 37042 34018 37054
rect 33966 36978 34018 36990
rect 1344 36874 46592 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 46592 36874
rect 1344 36788 46592 36822
rect 3614 36706 3666 36718
rect 3614 36642 3666 36654
rect 8878 36706 8930 36718
rect 8878 36642 8930 36654
rect 20190 36594 20242 36606
rect 3826 36542 3838 36594
rect 3890 36542 3902 36594
rect 5618 36542 5630 36594
rect 5682 36542 5694 36594
rect 12450 36542 12462 36594
rect 12514 36542 12526 36594
rect 14242 36542 14254 36594
rect 14306 36542 14318 36594
rect 16370 36542 16382 36594
rect 16434 36542 16446 36594
rect 19842 36542 19854 36594
rect 19906 36542 19918 36594
rect 20190 36530 20242 36542
rect 21422 36594 21474 36606
rect 27246 36594 27298 36606
rect 45502 36594 45554 36606
rect 21858 36542 21870 36594
rect 21922 36591 21934 36594
rect 22082 36591 22094 36594
rect 21922 36545 22094 36591
rect 21922 36542 21934 36545
rect 22082 36542 22094 36545
rect 22146 36542 22158 36594
rect 29250 36542 29262 36594
rect 29314 36542 29326 36594
rect 31490 36542 31502 36594
rect 31554 36542 31566 36594
rect 33618 36542 33630 36594
rect 33682 36542 33694 36594
rect 36194 36542 36206 36594
rect 36258 36542 36270 36594
rect 37986 36542 37998 36594
rect 38050 36542 38062 36594
rect 40226 36542 40238 36594
rect 40290 36542 40302 36594
rect 42354 36542 42366 36594
rect 42418 36591 42430 36594
rect 42418 36545 42639 36591
rect 42418 36542 42430 36545
rect 21422 36530 21474 36542
rect 27246 36530 27298 36542
rect 2830 36482 2882 36494
rect 2830 36418 2882 36430
rect 3054 36482 3106 36494
rect 16718 36482 16770 36494
rect 17390 36482 17442 36494
rect 3266 36430 3278 36482
rect 3330 36430 3342 36482
rect 4946 36430 4958 36482
rect 5010 36430 5022 36482
rect 8530 36430 8542 36482
rect 8594 36430 8606 36482
rect 9650 36430 9662 36482
rect 9714 36430 9726 36482
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 17042 36430 17054 36482
rect 17106 36430 17118 36482
rect 3054 36418 3106 36430
rect 16718 36418 16770 36430
rect 17390 36418 17442 36430
rect 18286 36482 18338 36494
rect 18286 36418 18338 36430
rect 20750 36482 20802 36494
rect 22318 36482 22370 36494
rect 21858 36430 21870 36482
rect 21922 36430 21934 36482
rect 20750 36418 20802 36430
rect 22318 36418 22370 36430
rect 23214 36482 23266 36494
rect 23214 36418 23266 36430
rect 23550 36482 23602 36494
rect 23550 36418 23602 36430
rect 23886 36482 23938 36494
rect 23886 36418 23938 36430
rect 26910 36482 26962 36494
rect 34974 36482 35026 36494
rect 42478 36482 42530 36494
rect 30818 36430 30830 36482
rect 30882 36430 30894 36482
rect 38434 36430 38446 36482
rect 38498 36430 38510 36482
rect 39442 36430 39454 36482
rect 39506 36430 39518 36482
rect 40562 36430 40574 36482
rect 40626 36430 40638 36482
rect 41458 36430 41470 36482
rect 41522 36430 41534 36482
rect 26910 36418 26962 36430
rect 34974 36418 35026 36430
rect 42478 36418 42530 36430
rect 2718 36370 2770 36382
rect 9102 36370 9154 36382
rect 18398 36370 18450 36382
rect 7746 36318 7758 36370
rect 7810 36318 7822 36370
rect 10322 36318 10334 36370
rect 10386 36318 10398 36370
rect 2718 36306 2770 36318
rect 9102 36306 9154 36318
rect 18398 36306 18450 36318
rect 18510 36370 18562 36382
rect 18510 36306 18562 36318
rect 18958 36370 19010 36382
rect 18958 36306 19010 36318
rect 19182 36370 19234 36382
rect 19182 36306 19234 36318
rect 19518 36370 19570 36382
rect 19518 36306 19570 36318
rect 20638 36370 20690 36382
rect 20638 36306 20690 36318
rect 22654 36370 22706 36382
rect 22654 36306 22706 36318
rect 23662 36370 23714 36382
rect 23662 36306 23714 36318
rect 26014 36370 26066 36382
rect 26014 36306 26066 36318
rect 29598 36370 29650 36382
rect 29598 36306 29650 36318
rect 29822 36370 29874 36382
rect 29822 36306 29874 36318
rect 30270 36370 30322 36382
rect 30270 36306 30322 36318
rect 34414 36370 34466 36382
rect 34414 36306 34466 36318
rect 35310 36370 35362 36382
rect 35310 36306 35362 36318
rect 36430 36370 36482 36382
rect 36430 36306 36482 36318
rect 41918 36370 41970 36382
rect 42593 36367 42639 36545
rect 43586 36542 43598 36594
rect 43650 36542 43662 36594
rect 45502 36530 45554 36542
rect 45166 36482 45218 36494
rect 42802 36430 42814 36482
rect 42866 36430 42878 36482
rect 43922 36430 43934 36482
rect 43986 36430 43998 36482
rect 45166 36418 45218 36430
rect 44830 36370 44882 36382
rect 42802 36367 42814 36370
rect 42593 36321 42814 36367
rect 42802 36318 42814 36321
rect 42866 36318 42878 36370
rect 43810 36318 43822 36370
rect 43874 36318 43886 36370
rect 41918 36306 41970 36318
rect 44830 36306 44882 36318
rect 46174 36370 46226 36382
rect 46174 36306 46226 36318
rect 3838 36258 3890 36270
rect 3838 36194 3890 36206
rect 4734 36258 4786 36270
rect 4734 36194 4786 36206
rect 8990 36258 9042 36270
rect 8990 36194 9042 36206
rect 13022 36258 13074 36270
rect 13022 36194 13074 36206
rect 17166 36258 17218 36270
rect 17166 36194 17218 36206
rect 17278 36258 17330 36270
rect 19406 36258 19458 36270
rect 17826 36206 17838 36258
rect 17890 36206 17902 36258
rect 17278 36194 17330 36206
rect 19406 36194 19458 36206
rect 20414 36258 20466 36270
rect 20414 36194 20466 36206
rect 21310 36258 21362 36270
rect 21310 36194 21362 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 22878 36258 22930 36270
rect 22878 36194 22930 36206
rect 23102 36258 23154 36270
rect 23102 36194 23154 36206
rect 24446 36258 24498 36270
rect 24446 36194 24498 36206
rect 25230 36258 25282 36270
rect 25230 36194 25282 36206
rect 26910 36258 26962 36270
rect 26910 36194 26962 36206
rect 28702 36258 28754 36270
rect 28702 36194 28754 36206
rect 29262 36258 29314 36270
rect 29262 36194 29314 36206
rect 29374 36258 29426 36270
rect 29374 36194 29426 36206
rect 30158 36258 30210 36270
rect 30158 36194 30210 36206
rect 34302 36258 34354 36270
rect 34302 36194 34354 36206
rect 34638 36258 34690 36270
rect 34638 36194 34690 36206
rect 34862 36258 34914 36270
rect 34862 36194 34914 36206
rect 35422 36258 35474 36270
rect 35422 36194 35474 36206
rect 35646 36258 35698 36270
rect 35646 36194 35698 36206
rect 41806 36258 41858 36270
rect 41806 36194 41858 36206
rect 42030 36258 42082 36270
rect 42030 36194 42082 36206
rect 43038 36258 43090 36270
rect 43038 36194 43090 36206
rect 44942 36258 44994 36270
rect 44942 36194 44994 36206
rect 45390 36258 45442 36270
rect 45390 36194 45442 36206
rect 45838 36258 45890 36270
rect 45838 36194 45890 36206
rect 1344 36090 46592 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 46592 36090
rect 1344 36004 46592 36038
rect 5854 35922 5906 35934
rect 5854 35858 5906 35870
rect 6974 35922 7026 35934
rect 6974 35858 7026 35870
rect 15710 35922 15762 35934
rect 15710 35858 15762 35870
rect 16494 35922 16546 35934
rect 16494 35858 16546 35870
rect 25230 35922 25282 35934
rect 25230 35858 25282 35870
rect 27134 35922 27186 35934
rect 27134 35858 27186 35870
rect 31054 35922 31106 35934
rect 31054 35858 31106 35870
rect 31278 35922 31330 35934
rect 31278 35858 31330 35870
rect 32174 35922 32226 35934
rect 32174 35858 32226 35870
rect 36990 35922 37042 35934
rect 36990 35858 37042 35870
rect 41022 35922 41074 35934
rect 41022 35858 41074 35870
rect 5742 35810 5794 35822
rect 17502 35810 17554 35822
rect 30718 35810 30770 35822
rect 2482 35758 2494 35810
rect 2546 35758 2558 35810
rect 7858 35758 7870 35810
rect 7922 35758 7934 35810
rect 16818 35758 16830 35810
rect 16882 35758 16894 35810
rect 28242 35758 28254 35810
rect 28306 35758 28318 35810
rect 5742 35746 5794 35758
rect 17502 35746 17554 35758
rect 30718 35746 30770 35758
rect 31166 35810 31218 35822
rect 31166 35746 31218 35758
rect 32510 35810 32562 35822
rect 40910 35810 40962 35822
rect 33842 35758 33854 35810
rect 33906 35758 33918 35810
rect 32510 35746 32562 35758
rect 40910 35746 40962 35758
rect 6750 35698 6802 35710
rect 15374 35698 15426 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 7746 35646 7758 35698
rect 7810 35646 7822 35698
rect 8418 35646 8430 35698
rect 8482 35646 8494 35698
rect 8978 35646 8990 35698
rect 9042 35646 9054 35698
rect 14690 35646 14702 35698
rect 14754 35646 14766 35698
rect 6750 35634 6802 35646
rect 15374 35634 15426 35646
rect 15598 35698 15650 35710
rect 15598 35634 15650 35646
rect 15710 35698 15762 35710
rect 15710 35634 15762 35646
rect 17614 35698 17666 35710
rect 25342 35698 25394 35710
rect 17938 35646 17950 35698
rect 18002 35646 18014 35698
rect 20402 35646 20414 35698
rect 20466 35646 20478 35698
rect 17614 35634 17666 35646
rect 25342 35634 25394 35646
rect 26238 35698 26290 35710
rect 26238 35634 26290 35646
rect 26686 35698 26738 35710
rect 30942 35698 30994 35710
rect 32062 35698 32114 35710
rect 27458 35646 27470 35698
rect 27522 35646 27534 35698
rect 31826 35646 31838 35698
rect 31890 35646 31902 35698
rect 26686 35634 26738 35646
rect 30942 35634 30994 35646
rect 32062 35634 32114 35646
rect 32286 35698 32338 35710
rect 36654 35698 36706 35710
rect 33058 35646 33070 35698
rect 33122 35646 33134 35698
rect 32286 35634 32338 35646
rect 36654 35634 36706 35646
rect 36878 35698 36930 35710
rect 36878 35634 36930 35646
rect 37214 35698 37266 35710
rect 41246 35698 41298 35710
rect 37538 35646 37550 35698
rect 37602 35646 37614 35698
rect 42242 35646 42254 35698
rect 42306 35646 42318 35698
rect 42914 35646 42926 35698
rect 42978 35646 42990 35698
rect 43362 35646 43374 35698
rect 43426 35646 43438 35698
rect 37214 35634 37266 35646
rect 41246 35634 41298 35646
rect 5294 35586 5346 35598
rect 4610 35534 4622 35586
rect 4674 35534 4686 35586
rect 5294 35522 5346 35534
rect 5966 35586 6018 35598
rect 5966 35522 6018 35534
rect 6526 35586 6578 35598
rect 6526 35522 6578 35534
rect 6862 35586 6914 35598
rect 25902 35586 25954 35598
rect 7634 35534 7646 35586
rect 7698 35534 7710 35586
rect 9762 35534 9774 35586
rect 9826 35534 9838 35586
rect 21858 35534 21870 35586
rect 21922 35534 21934 35586
rect 30370 35534 30382 35586
rect 30434 35534 30446 35586
rect 35970 35534 35982 35586
rect 36034 35534 36046 35586
rect 38210 35534 38222 35586
rect 38274 35534 38286 35586
rect 40338 35534 40350 35586
rect 40402 35534 40414 35586
rect 42130 35534 42142 35586
rect 42194 35534 42206 35586
rect 44034 35534 44046 35586
rect 44098 35534 44110 35586
rect 46162 35534 46174 35586
rect 46226 35534 46238 35586
rect 6862 35522 6914 35534
rect 25902 35522 25954 35534
rect 5182 35474 5234 35486
rect 5182 35410 5234 35422
rect 6302 35474 6354 35486
rect 42018 35422 42030 35474
rect 42082 35422 42094 35474
rect 6302 35410 6354 35422
rect 1344 35306 46592 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 46592 35306
rect 1344 35220 46592 35254
rect 7198 35138 7250 35150
rect 7198 35074 7250 35086
rect 29374 35138 29426 35150
rect 29374 35074 29426 35086
rect 35534 35138 35586 35150
rect 35534 35074 35586 35086
rect 36094 35138 36146 35150
rect 36094 35074 36146 35086
rect 37550 35138 37602 35150
rect 37550 35074 37602 35086
rect 43150 35138 43202 35150
rect 43150 35074 43202 35086
rect 44942 35138 44994 35150
rect 44942 35074 44994 35086
rect 3054 35026 3106 35038
rect 3054 34962 3106 34974
rect 4846 35026 4898 35038
rect 17838 35026 17890 35038
rect 36318 35026 36370 35038
rect 46174 35026 46226 35038
rect 8082 34974 8094 35026
rect 8146 34974 8158 35026
rect 9650 34974 9662 35026
rect 9714 34974 9726 35026
rect 13682 34974 13694 35026
rect 13746 34974 13758 35026
rect 15810 34974 15822 35026
rect 15874 34974 15886 35026
rect 24658 34974 24670 35026
rect 24722 34974 24734 35026
rect 27906 34974 27918 35026
rect 27970 34974 27982 35026
rect 30258 34974 30270 35026
rect 30322 34974 30334 35026
rect 35858 34974 35870 35026
rect 35922 34974 35934 35026
rect 38434 34974 38446 35026
rect 38498 34974 38510 35026
rect 39554 34974 39566 35026
rect 39618 34974 39630 35026
rect 4846 34962 4898 34974
rect 17838 34962 17890 34974
rect 36318 34962 36370 34974
rect 46174 34962 46226 34974
rect 3278 34914 3330 34926
rect 3278 34850 3330 34862
rect 3950 34914 4002 34926
rect 3950 34850 4002 34862
rect 4062 34914 4114 34926
rect 7646 34914 7698 34926
rect 16942 34914 16994 34926
rect 35646 34914 35698 34926
rect 4386 34862 4398 34914
rect 4450 34862 4462 34914
rect 7858 34862 7870 34914
rect 7922 34862 7934 34914
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 12562 34862 12574 34914
rect 12626 34862 12638 34914
rect 16594 34862 16606 34914
rect 16658 34862 16670 34914
rect 20626 34862 20638 34914
rect 20690 34862 20702 34914
rect 21858 34862 21870 34914
rect 21922 34862 21934 34914
rect 25106 34862 25118 34914
rect 25170 34862 25182 34914
rect 34738 34862 34750 34914
rect 34802 34862 34814 34914
rect 4062 34850 4114 34862
rect 7646 34850 7698 34862
rect 16942 34850 16994 34862
rect 35646 34850 35698 34862
rect 37214 34914 37266 34926
rect 37214 34850 37266 34862
rect 37774 34914 37826 34926
rect 41134 34914 41186 34926
rect 38994 34862 39006 34914
rect 39058 34862 39070 34914
rect 37774 34850 37826 34862
rect 41134 34850 41186 34862
rect 43710 34914 43762 34926
rect 43710 34850 43762 34862
rect 43934 34914 43986 34926
rect 43934 34850 43986 34862
rect 45390 34914 45442 34926
rect 45390 34850 45442 34862
rect 45614 34914 45666 34926
rect 45614 34850 45666 34862
rect 2942 34802 2994 34814
rect 2942 34738 2994 34750
rect 3502 34802 3554 34814
rect 7198 34802 7250 34814
rect 4274 34750 4286 34802
rect 4338 34750 4350 34802
rect 3502 34738 3554 34750
rect 7198 34738 7250 34750
rect 7310 34802 7362 34814
rect 7310 34738 7362 34750
rect 9326 34802 9378 34814
rect 29262 34802 29314 34814
rect 11778 34750 11790 34802
rect 11842 34750 11854 34802
rect 19954 34750 19966 34802
rect 20018 34750 20030 34802
rect 22530 34750 22542 34802
rect 22594 34750 22606 34802
rect 25778 34750 25790 34802
rect 25842 34750 25854 34802
rect 9326 34738 9378 34750
rect 29262 34738 29314 34750
rect 36990 34802 37042 34814
rect 36990 34738 37042 34750
rect 37326 34802 37378 34814
rect 37326 34738 37378 34750
rect 38670 34802 38722 34814
rect 38670 34738 38722 34750
rect 39678 34802 39730 34814
rect 43374 34802 43426 34814
rect 42690 34750 42702 34802
rect 42754 34750 42766 34802
rect 39678 34738 39730 34750
rect 43374 34738 43426 34750
rect 43486 34802 43538 34814
rect 43486 34738 43538 34750
rect 44830 34802 44882 34814
rect 44830 34738 44882 34750
rect 45054 34802 45106 34814
rect 45054 34738 45106 34750
rect 17278 34690 17330 34702
rect 17278 34626 17330 34638
rect 21534 34690 21586 34702
rect 21534 34626 21586 34638
rect 28590 34690 28642 34702
rect 28590 34626 28642 34638
rect 46062 34690 46114 34702
rect 46062 34626 46114 34638
rect 1344 34522 46592 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 46592 34522
rect 1344 34436 46592 34470
rect 2830 34354 2882 34366
rect 2830 34290 2882 34302
rect 2942 34354 2994 34366
rect 5070 34354 5122 34366
rect 3938 34302 3950 34354
rect 4002 34302 4014 34354
rect 2942 34290 2994 34302
rect 5070 34290 5122 34302
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 9102 34354 9154 34366
rect 9102 34290 9154 34302
rect 9886 34354 9938 34366
rect 9886 34290 9938 34302
rect 9998 34354 10050 34366
rect 9998 34290 10050 34302
rect 10446 34354 10498 34366
rect 10446 34290 10498 34302
rect 11118 34354 11170 34366
rect 11118 34290 11170 34302
rect 11902 34354 11954 34366
rect 11902 34290 11954 34302
rect 12014 34354 12066 34366
rect 12014 34290 12066 34302
rect 12574 34354 12626 34366
rect 12574 34290 12626 34302
rect 13022 34354 13074 34366
rect 13022 34290 13074 34302
rect 13806 34354 13858 34366
rect 13806 34290 13858 34302
rect 14926 34354 14978 34366
rect 14926 34290 14978 34302
rect 16494 34354 16546 34366
rect 16494 34290 16546 34302
rect 17390 34354 17442 34366
rect 17390 34290 17442 34302
rect 19070 34354 19122 34366
rect 19070 34290 19122 34302
rect 19294 34354 19346 34366
rect 19294 34290 19346 34302
rect 20414 34354 20466 34366
rect 20414 34290 20466 34302
rect 21422 34354 21474 34366
rect 22990 34354 23042 34366
rect 22642 34302 22654 34354
rect 22706 34302 22718 34354
rect 21422 34290 21474 34302
rect 22990 34290 23042 34302
rect 25342 34354 25394 34366
rect 25342 34290 25394 34302
rect 26350 34354 26402 34366
rect 26350 34290 26402 34302
rect 26910 34354 26962 34366
rect 26910 34290 26962 34302
rect 27358 34354 27410 34366
rect 27358 34290 27410 34302
rect 27806 34354 27858 34366
rect 27806 34290 27858 34302
rect 32174 34354 32226 34366
rect 32174 34290 32226 34302
rect 33294 34354 33346 34366
rect 33294 34290 33346 34302
rect 33406 34354 33458 34366
rect 33406 34290 33458 34302
rect 35534 34354 35586 34366
rect 35534 34290 35586 34302
rect 40238 34354 40290 34366
rect 44818 34302 44830 34354
rect 44882 34302 44894 34354
rect 40238 34290 40290 34302
rect 4398 34242 4450 34254
rect 4398 34178 4450 34190
rect 4622 34242 4674 34254
rect 4622 34178 4674 34190
rect 6302 34242 6354 34254
rect 6302 34178 6354 34190
rect 6862 34242 6914 34254
rect 6862 34178 6914 34190
rect 7422 34242 7474 34254
rect 7422 34178 7474 34190
rect 8206 34242 8258 34254
rect 8206 34178 8258 34190
rect 11454 34242 11506 34254
rect 11454 34178 11506 34190
rect 11678 34242 11730 34254
rect 11678 34178 11730 34190
rect 18958 34242 19010 34254
rect 18958 34178 19010 34190
rect 20750 34242 20802 34254
rect 20750 34178 20802 34190
rect 20862 34242 20914 34254
rect 20862 34178 20914 34190
rect 24334 34242 24386 34254
rect 24334 34178 24386 34190
rect 24446 34242 24498 34254
rect 24446 34178 24498 34190
rect 25230 34242 25282 34254
rect 25230 34178 25282 34190
rect 26462 34242 26514 34254
rect 26462 34178 26514 34190
rect 32510 34242 32562 34254
rect 32510 34178 32562 34190
rect 33518 34242 33570 34254
rect 34862 34242 34914 34254
rect 34066 34190 34078 34242
rect 34130 34190 34142 34242
rect 33518 34178 33570 34190
rect 34862 34178 34914 34190
rect 35198 34242 35250 34254
rect 35198 34178 35250 34190
rect 35310 34242 35362 34254
rect 39006 34242 39058 34254
rect 36530 34190 36542 34242
rect 36594 34190 36606 34242
rect 35310 34178 35362 34190
rect 39006 34178 39058 34190
rect 39342 34242 39394 34254
rect 39342 34178 39394 34190
rect 40350 34242 40402 34254
rect 44270 34242 44322 34254
rect 41682 34190 41694 34242
rect 41746 34190 41758 34242
rect 46162 34190 46174 34242
rect 46226 34190 46238 34242
rect 40350 34178 40402 34190
rect 44270 34178 44322 34190
rect 1934 34130 1986 34142
rect 1934 34066 1986 34078
rect 2158 34130 2210 34142
rect 2158 34066 2210 34078
rect 2494 34130 2546 34142
rect 2494 34066 2546 34078
rect 2718 34130 2770 34142
rect 4510 34130 4562 34142
rect 5854 34130 5906 34142
rect 3266 34078 3278 34130
rect 3330 34078 3342 34130
rect 5282 34078 5294 34130
rect 5346 34078 5358 34130
rect 2718 34066 2770 34078
rect 4510 34066 4562 34078
rect 5854 34066 5906 34078
rect 6414 34130 6466 34142
rect 6414 34066 6466 34078
rect 6974 34130 7026 34142
rect 6974 34066 7026 34078
rect 7198 34130 7250 34142
rect 7198 34066 7250 34078
rect 7758 34130 7810 34142
rect 7758 34066 7810 34078
rect 7982 34130 8034 34142
rect 7982 34066 8034 34078
rect 9438 34130 9490 34142
rect 9438 34066 9490 34078
rect 10110 34130 10162 34142
rect 10110 34066 10162 34078
rect 10558 34130 10610 34142
rect 13582 34130 13634 34142
rect 13346 34078 13358 34130
rect 13410 34078 13422 34130
rect 10558 34066 10610 34078
rect 13582 34066 13634 34078
rect 13918 34130 13970 34142
rect 13918 34066 13970 34078
rect 21086 34130 21138 34142
rect 21086 34066 21138 34078
rect 21310 34130 21362 34142
rect 21310 34066 21362 34078
rect 21534 34130 21586 34142
rect 21534 34066 21586 34078
rect 21982 34130 22034 34142
rect 21982 34066 22034 34078
rect 22318 34130 22370 34142
rect 22318 34066 22370 34078
rect 23326 34130 23378 34142
rect 23326 34066 23378 34078
rect 23774 34130 23826 34142
rect 23774 34066 23826 34078
rect 24110 34130 24162 34142
rect 32062 34130 32114 34142
rect 31154 34078 31166 34130
rect 31218 34078 31230 34130
rect 31826 34078 31838 34130
rect 31890 34078 31902 34130
rect 24110 34066 24162 34078
rect 32062 34066 32114 34078
rect 32286 34130 32338 34142
rect 33630 34130 33682 34142
rect 33058 34078 33070 34130
rect 33122 34078 33134 34130
rect 32286 34066 32338 34078
rect 33630 34066 33682 34078
rect 34414 34130 34466 34142
rect 39118 34130 39170 34142
rect 35858 34078 35870 34130
rect 35922 34078 35934 34130
rect 34414 34066 34466 34078
rect 39118 34066 39170 34078
rect 39566 34130 39618 34142
rect 44158 34130 44210 34142
rect 40898 34078 40910 34130
rect 40962 34078 40974 34130
rect 39566 34066 39618 34078
rect 44158 34066 44210 34078
rect 44494 34130 44546 34142
rect 45154 34078 45166 34130
rect 45218 34078 45230 34130
rect 45602 34078 45614 34130
rect 45666 34078 45678 34130
rect 44494 34066 44546 34078
rect 2270 34018 2322 34030
rect 2270 33954 2322 33966
rect 6078 34018 6130 34030
rect 6078 33954 6130 33966
rect 11006 34018 11058 34030
rect 11006 33954 11058 33966
rect 11790 34018 11842 34030
rect 11790 33954 11842 33966
rect 13694 34018 13746 34030
rect 13694 33954 13746 33966
rect 14590 34018 14642 34030
rect 14590 33954 14642 33966
rect 15486 34018 15538 34030
rect 15486 33954 15538 33966
rect 15934 34018 15986 34030
rect 15934 33954 15986 33966
rect 16942 34018 16994 34030
rect 16942 33954 16994 33966
rect 17502 34018 17554 34030
rect 17502 33954 17554 33966
rect 18062 34018 18114 34030
rect 18062 33954 18114 33966
rect 18622 34018 18674 34030
rect 18622 33954 18674 33966
rect 19966 34018 20018 34030
rect 19966 33954 20018 33966
rect 26014 34018 26066 34030
rect 28354 33966 28366 34018
rect 28418 33966 28430 34018
rect 30482 33966 30494 34018
rect 30546 33966 30558 34018
rect 38658 33966 38670 34018
rect 38722 33966 38734 34018
rect 43810 33966 43822 34018
rect 43874 33966 43886 34018
rect 45490 33966 45502 34018
rect 45554 33966 45566 34018
rect 26014 33954 26066 33966
rect 17950 33906 18002 33918
rect 17950 33842 18002 33854
rect 23102 33906 23154 33918
rect 23102 33842 23154 33854
rect 23886 33906 23938 33918
rect 23886 33842 23938 33854
rect 25342 33906 25394 33918
rect 25342 33842 25394 33854
rect 25902 33906 25954 33918
rect 25902 33842 25954 33854
rect 34750 33906 34802 33918
rect 34750 33842 34802 33854
rect 39790 33906 39842 33918
rect 39790 33842 39842 33854
rect 1344 33738 46592 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 46592 33738
rect 1344 33652 46592 33686
rect 21646 33570 21698 33582
rect 10770 33518 10782 33570
rect 10834 33518 10846 33570
rect 9438 33458 9490 33470
rect 2482 33406 2494 33458
rect 2546 33406 2558 33458
rect 4610 33406 4622 33458
rect 4674 33406 4686 33458
rect 6402 33406 6414 33458
rect 6466 33406 6478 33458
rect 8530 33406 8542 33458
rect 8594 33406 8606 33458
rect 9438 33394 9490 33406
rect 10334 33346 10386 33358
rect 1810 33294 1822 33346
rect 1874 33294 1886 33346
rect 5618 33294 5630 33346
rect 5682 33294 5694 33346
rect 9986 33294 9998 33346
rect 10050 33294 10062 33346
rect 10334 33282 10386 33294
rect 10785 33119 10831 33518
rect 21646 33506 21698 33518
rect 21982 33570 22034 33582
rect 21982 33506 22034 33518
rect 44830 33570 44882 33582
rect 44830 33506 44882 33518
rect 44942 33570 44994 33582
rect 44942 33506 44994 33518
rect 45390 33570 45442 33582
rect 45390 33506 45442 33518
rect 45614 33570 45666 33582
rect 45614 33506 45666 33518
rect 46062 33570 46114 33582
rect 46062 33506 46114 33518
rect 11790 33458 11842 33470
rect 11790 33394 11842 33406
rect 12798 33458 12850 33470
rect 28254 33458 28306 33470
rect 46174 33458 46226 33470
rect 16370 33406 16382 33458
rect 16434 33406 16446 33458
rect 17490 33406 17502 33458
rect 17554 33406 17566 33458
rect 19618 33406 19630 33458
rect 19682 33406 19694 33458
rect 25442 33406 25454 33458
rect 25506 33406 25518 33458
rect 27570 33406 27582 33458
rect 27634 33406 27646 33458
rect 30034 33406 30046 33458
rect 30098 33406 30110 33458
rect 32722 33406 32734 33458
rect 32786 33406 32798 33458
rect 34850 33406 34862 33458
rect 34914 33406 34926 33458
rect 40450 33406 40462 33458
rect 40514 33406 40526 33458
rect 12798 33394 12850 33406
rect 28254 33394 28306 33406
rect 46174 33394 46226 33406
rect 22430 33346 22482 33358
rect 13458 33294 13470 33346
rect 13522 33294 13534 33346
rect 16818 33294 16830 33346
rect 16882 33294 16894 33346
rect 21970 33294 21982 33346
rect 22034 33294 22046 33346
rect 22430 33282 22482 33294
rect 22990 33346 23042 33358
rect 28366 33346 28418 33358
rect 31502 33346 31554 33358
rect 24770 33294 24782 33346
rect 24834 33294 24846 33346
rect 27906 33294 27918 33346
rect 27970 33294 27982 33346
rect 28578 33294 28590 33346
rect 28642 33294 28654 33346
rect 29474 33294 29486 33346
rect 29538 33294 29550 33346
rect 30146 33294 30158 33346
rect 30210 33294 30222 33346
rect 31938 33294 31950 33346
rect 32002 33294 32014 33346
rect 35410 33294 35422 33346
rect 35474 33294 35486 33346
rect 37202 33294 37214 33346
rect 37266 33294 37278 33346
rect 42802 33294 42814 33346
rect 42866 33294 42878 33346
rect 22990 33282 23042 33294
rect 28366 33282 28418 33294
rect 31502 33282 31554 33294
rect 20414 33234 20466 33246
rect 14242 33182 14254 33234
rect 14306 33182 14318 33234
rect 20414 33170 20466 33182
rect 22766 33234 22818 33246
rect 24222 33234 24274 33246
rect 23314 33182 23326 33234
rect 23378 33182 23390 33234
rect 22766 33170 22818 33182
rect 24222 33170 24274 33182
rect 28142 33234 28194 33246
rect 28142 33170 28194 33182
rect 29710 33234 29762 33246
rect 36206 33234 36258 33246
rect 45054 33234 45106 33246
rect 30482 33182 30494 33234
rect 30546 33182 30558 33234
rect 31154 33182 31166 33234
rect 31218 33182 31230 33234
rect 35186 33182 35198 33234
rect 35250 33182 35262 33234
rect 36978 33182 36990 33234
rect 37042 33182 37054 33234
rect 38658 33182 38670 33234
rect 38722 33182 38734 33234
rect 29710 33170 29762 33182
rect 36206 33170 36258 33182
rect 45054 33170 45106 33182
rect 11118 33122 11170 33134
rect 10882 33119 10894 33122
rect 10785 33073 10894 33119
rect 10882 33070 10894 33073
rect 10946 33070 10958 33122
rect 11118 33058 11170 33070
rect 12238 33122 12290 33134
rect 12238 33058 12290 33070
rect 12910 33122 12962 33134
rect 12910 33058 12962 33070
rect 20862 33122 20914 33134
rect 20862 33058 20914 33070
rect 22542 33122 22594 33134
rect 22542 33058 22594 33070
rect 23662 33122 23714 33134
rect 23662 33058 23714 33070
rect 23886 33122 23938 33134
rect 23886 33058 23938 33070
rect 24110 33122 24162 33134
rect 24110 33058 24162 33070
rect 29934 33122 29986 33134
rect 29934 33058 29986 33070
rect 30830 33122 30882 33134
rect 30830 33058 30882 33070
rect 36094 33122 36146 33134
rect 37998 33122 38050 33134
rect 37650 33070 37662 33122
rect 37714 33070 37726 33122
rect 36094 33058 36146 33070
rect 37998 33058 38050 33070
rect 38334 33122 38386 33134
rect 38334 33058 38386 33070
rect 1344 32954 46592 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 46592 32954
rect 1344 32868 46592 32902
rect 11342 32786 11394 32798
rect 11342 32722 11394 32734
rect 15374 32786 15426 32798
rect 15374 32722 15426 32734
rect 16494 32786 16546 32798
rect 16494 32722 16546 32734
rect 17502 32786 17554 32798
rect 17502 32722 17554 32734
rect 18286 32786 18338 32798
rect 18286 32722 18338 32734
rect 19406 32786 19458 32798
rect 19406 32722 19458 32734
rect 23326 32786 23378 32798
rect 29150 32786 29202 32798
rect 23874 32734 23886 32786
rect 23938 32734 23950 32786
rect 23326 32722 23378 32734
rect 29150 32722 29202 32734
rect 30382 32786 30434 32798
rect 31950 32786 32002 32798
rect 31266 32734 31278 32786
rect 31330 32734 31342 32786
rect 30382 32722 30434 32734
rect 31950 32722 32002 32734
rect 39790 32786 39842 32798
rect 39790 32722 39842 32734
rect 41918 32786 41970 32798
rect 41918 32722 41970 32734
rect 42142 32786 42194 32798
rect 42142 32722 42194 32734
rect 17390 32674 17442 32686
rect 14018 32622 14030 32674
rect 14082 32622 14094 32674
rect 15586 32622 15598 32674
rect 15650 32671 15662 32674
rect 16034 32671 16046 32674
rect 15650 32625 16046 32671
rect 15650 32622 15662 32625
rect 16034 32622 16046 32625
rect 16098 32622 16110 32674
rect 17390 32610 17442 32622
rect 18622 32674 18674 32686
rect 29598 32674 29650 32686
rect 37886 32674 37938 32686
rect 19058 32622 19070 32674
rect 19122 32622 19134 32674
rect 26338 32622 26350 32674
rect 26402 32622 26414 32674
rect 33730 32622 33742 32674
rect 33794 32622 33806 32674
rect 18622 32610 18674 32622
rect 29598 32610 29650 32622
rect 37886 32610 37938 32622
rect 41806 32674 41858 32686
rect 41806 32610 41858 32622
rect 11118 32562 11170 32574
rect 15486 32562 15538 32574
rect 7522 32510 7534 32562
rect 7586 32510 7598 32562
rect 10882 32510 10894 32562
rect 10946 32510 10958 32562
rect 11554 32510 11566 32562
rect 11618 32510 11630 32562
rect 14802 32510 14814 32562
rect 14866 32510 14878 32562
rect 11118 32498 11170 32510
rect 15486 32498 15538 32510
rect 16270 32562 16322 32574
rect 16270 32498 16322 32510
rect 16382 32562 16434 32574
rect 16382 32498 16434 32510
rect 16606 32562 16658 32574
rect 16606 32498 16658 32510
rect 16718 32562 16770 32574
rect 18174 32562 18226 32574
rect 17938 32510 17950 32562
rect 18002 32510 18014 32562
rect 16718 32498 16770 32510
rect 18174 32498 18226 32510
rect 18398 32562 18450 32574
rect 22990 32562 23042 32574
rect 19730 32510 19742 32562
rect 19794 32510 19806 32562
rect 18398 32498 18450 32510
rect 22990 32498 23042 32510
rect 23326 32562 23378 32574
rect 23326 32498 23378 32510
rect 23550 32562 23602 32574
rect 23550 32498 23602 32510
rect 24222 32562 24274 32574
rect 24222 32498 24274 32510
rect 24558 32562 24610 32574
rect 24558 32498 24610 32510
rect 25454 32562 25506 32574
rect 27358 32562 27410 32574
rect 26562 32510 26574 32562
rect 26626 32510 26638 32562
rect 25454 32498 25506 32510
rect 27358 32498 27410 32510
rect 27582 32562 27634 32574
rect 27582 32498 27634 32510
rect 27806 32562 27858 32574
rect 27806 32498 27858 32510
rect 30942 32562 30994 32574
rect 32174 32562 32226 32574
rect 34078 32562 34130 32574
rect 38110 32562 38162 32574
rect 31714 32510 31726 32562
rect 31778 32510 31790 32562
rect 32386 32510 32398 32562
rect 32450 32510 32462 32562
rect 33394 32510 33406 32562
rect 33458 32510 33470 32562
rect 34738 32510 34750 32562
rect 34802 32510 34814 32562
rect 30942 32498 30994 32510
rect 32174 32498 32226 32510
rect 34078 32498 34130 32510
rect 38110 32498 38162 32510
rect 38446 32562 38498 32574
rect 38446 32498 38498 32510
rect 38894 32562 38946 32574
rect 38894 32498 38946 32510
rect 39006 32562 39058 32574
rect 39006 32498 39058 32510
rect 39454 32562 39506 32574
rect 42466 32510 42478 32562
rect 42530 32510 42542 32562
rect 43362 32510 43374 32562
rect 43426 32510 43438 32562
rect 39454 32498 39506 32510
rect 10558 32450 10610 32462
rect 27694 32450 27746 32462
rect 7970 32398 7982 32450
rect 8034 32398 8046 32450
rect 10994 32398 11006 32450
rect 11058 32398 11070 32450
rect 11890 32398 11902 32450
rect 11954 32398 11966 32450
rect 20514 32398 20526 32450
rect 20578 32398 20590 32450
rect 22642 32398 22654 32450
rect 22706 32398 22718 32450
rect 25890 32398 25902 32450
rect 25954 32398 25966 32450
rect 10558 32386 10610 32398
rect 27694 32386 27746 32398
rect 28254 32450 28306 32462
rect 28254 32386 28306 32398
rect 28814 32450 28866 32462
rect 37998 32450 38050 32462
rect 30482 32398 30494 32450
rect 30546 32398 30558 32450
rect 32274 32398 32286 32450
rect 32338 32398 32350 32450
rect 35410 32398 35422 32450
rect 35474 32398 35486 32450
rect 37538 32398 37550 32450
rect 37602 32398 37614 32450
rect 28814 32386 28866 32398
rect 37998 32386 38050 32398
rect 39230 32450 39282 32462
rect 39230 32386 39282 32398
rect 40238 32450 40290 32462
rect 40238 32386 40290 32398
rect 41022 32450 41074 32462
rect 41022 32386 41074 32398
rect 41470 32450 41522 32462
rect 42802 32398 42814 32450
rect 42866 32398 42878 32450
rect 44034 32398 44046 32450
rect 44098 32398 44110 32450
rect 46162 32398 46174 32450
rect 46226 32398 46238 32450
rect 41470 32386 41522 32398
rect 8766 32338 8818 32350
rect 8766 32274 8818 32286
rect 10446 32338 10498 32350
rect 10446 32274 10498 32286
rect 24670 32338 24722 32350
rect 24670 32274 24722 32286
rect 30158 32338 30210 32350
rect 30158 32274 30210 32286
rect 33070 32338 33122 32350
rect 33070 32274 33122 32286
rect 33406 32338 33458 32350
rect 33406 32274 33458 32286
rect 1344 32170 46592 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 46592 32170
rect 1344 32084 46592 32118
rect 28030 32002 28082 32014
rect 16818 31950 16830 32002
rect 16882 31999 16894 32002
rect 18274 31999 18286 32002
rect 16882 31953 18286 31999
rect 16882 31950 16894 31953
rect 18274 31950 18286 31953
rect 18338 31950 18350 32002
rect 28030 31938 28082 31950
rect 16270 31890 16322 31902
rect 4610 31838 4622 31890
rect 4674 31838 4686 31890
rect 9538 31838 9550 31890
rect 9602 31838 9614 31890
rect 11666 31838 11678 31890
rect 11730 31838 11742 31890
rect 16270 31826 16322 31838
rect 16830 31890 16882 31902
rect 16830 31826 16882 31838
rect 19854 31890 19906 31902
rect 19854 31826 19906 31838
rect 27358 31890 27410 31902
rect 27358 31826 27410 31838
rect 29262 31890 29314 31902
rect 29262 31826 29314 31838
rect 29710 31890 29762 31902
rect 35646 31890 35698 31902
rect 31042 31838 31054 31890
rect 31106 31838 31118 31890
rect 33170 31838 33182 31890
rect 33234 31838 33246 31890
rect 29710 31826 29762 31838
rect 35646 31826 35698 31838
rect 37102 31890 37154 31902
rect 44942 31890 44994 31902
rect 42130 31838 42142 31890
rect 42194 31838 42206 31890
rect 43810 31838 43822 31890
rect 43874 31838 43886 31890
rect 37102 31826 37154 31838
rect 44942 31826 44994 31838
rect 45390 31890 45442 31902
rect 45390 31826 45442 31838
rect 8430 31778 8482 31790
rect 13918 31778 13970 31790
rect 17278 31778 17330 31790
rect 1810 31726 1822 31778
rect 1874 31726 1886 31778
rect 8866 31726 8878 31778
rect 8930 31726 8942 31778
rect 14130 31726 14142 31778
rect 14194 31726 14206 31778
rect 8430 31714 8482 31726
rect 13918 31714 13970 31726
rect 17278 31714 17330 31726
rect 20190 31778 20242 31790
rect 20190 31714 20242 31726
rect 20862 31778 20914 31790
rect 27246 31778 27298 31790
rect 21298 31726 21310 31778
rect 21362 31726 21374 31778
rect 20862 31714 20914 31726
rect 27246 31714 27298 31726
rect 27470 31778 27522 31790
rect 34302 31778 34354 31790
rect 33954 31726 33966 31778
rect 34018 31726 34030 31778
rect 27470 31714 27522 31726
rect 34302 31714 34354 31726
rect 34862 31778 34914 31790
rect 34862 31714 34914 31726
rect 35534 31778 35586 31790
rect 35534 31714 35586 31726
rect 36094 31778 36146 31790
rect 36094 31714 36146 31726
rect 37326 31778 37378 31790
rect 37326 31714 37378 31726
rect 37662 31778 37714 31790
rect 37662 31714 37714 31726
rect 37886 31778 37938 31790
rect 42478 31778 42530 31790
rect 39330 31726 39342 31778
rect 39394 31726 39406 31778
rect 37886 31714 37938 31726
rect 42478 31714 42530 31726
rect 43038 31778 43090 31790
rect 43038 31714 43090 31726
rect 5854 31666 5906 31678
rect 2482 31614 2494 31666
rect 2546 31614 2558 31666
rect 5854 31602 5906 31614
rect 6302 31666 6354 31678
rect 6302 31602 6354 31614
rect 6638 31666 6690 31678
rect 6638 31602 6690 31614
rect 6862 31666 6914 31678
rect 6862 31602 6914 31614
rect 7198 31666 7250 31678
rect 7198 31602 7250 31614
rect 7422 31666 7474 31678
rect 7422 31602 7474 31614
rect 7758 31666 7810 31678
rect 7758 31602 7810 31614
rect 13470 31666 13522 31678
rect 15822 31666 15874 31678
rect 14466 31614 14478 31666
rect 14530 31614 14542 31666
rect 13470 31602 13522 31614
rect 15822 31602 15874 31614
rect 18510 31666 18562 31678
rect 18510 31602 18562 31614
rect 19406 31666 19458 31678
rect 19406 31602 19458 31614
rect 20414 31666 20466 31678
rect 27022 31666 27074 31678
rect 23314 31614 23326 31666
rect 23378 31614 23390 31666
rect 20414 31602 20466 31614
rect 27022 31602 27074 31614
rect 28142 31666 28194 31678
rect 28142 31602 28194 31614
rect 28590 31666 28642 31678
rect 30718 31666 30770 31678
rect 30370 31614 30382 31666
rect 30434 31614 30446 31666
rect 28590 31602 28642 31614
rect 30718 31602 30770 31614
rect 35870 31666 35922 31678
rect 35870 31602 35922 31614
rect 37550 31666 37602 31678
rect 38658 31614 38670 31666
rect 38722 31614 38734 31666
rect 40002 31614 40014 31666
rect 40066 31614 40078 31666
rect 37550 31602 37602 31614
rect 5518 31554 5570 31566
rect 5518 31490 5570 31502
rect 5742 31554 5794 31566
rect 5742 31490 5794 31502
rect 6414 31554 6466 31566
rect 6414 31490 6466 31502
rect 6974 31554 7026 31566
rect 6974 31490 7026 31502
rect 7870 31554 7922 31566
rect 7870 31490 7922 31502
rect 8094 31554 8146 31566
rect 8094 31490 8146 31502
rect 12574 31554 12626 31566
rect 12574 31490 12626 31502
rect 13022 31554 13074 31566
rect 13022 31490 13074 31502
rect 13694 31554 13746 31566
rect 13694 31490 13746 31502
rect 13806 31554 13858 31566
rect 13806 31490 13858 31502
rect 14814 31554 14866 31566
rect 14814 31490 14866 31502
rect 15486 31554 15538 31566
rect 15486 31490 15538 31502
rect 15710 31554 15762 31566
rect 15710 31490 15762 31502
rect 17838 31554 17890 31566
rect 17838 31490 17890 31502
rect 18174 31554 18226 31566
rect 18174 31490 18226 31502
rect 18622 31554 18674 31566
rect 18622 31490 18674 31502
rect 20526 31554 20578 31566
rect 20526 31490 20578 31502
rect 28366 31554 28418 31566
rect 28366 31490 28418 31502
rect 38334 31554 38386 31566
rect 38334 31490 38386 31502
rect 43374 31554 43426 31566
rect 43374 31490 43426 31502
rect 45950 31554 46002 31566
rect 45950 31490 46002 31502
rect 1344 31386 46592 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 46592 31386
rect 1344 31300 46592 31334
rect 9550 31218 9602 31230
rect 34078 31218 34130 31230
rect 21410 31166 21422 31218
rect 21474 31166 21486 31218
rect 9550 31154 9602 31166
rect 34078 31154 34130 31166
rect 41022 31218 41074 31230
rect 41022 31154 41074 31166
rect 41806 31218 41858 31230
rect 44494 31218 44546 31230
rect 42578 31166 42590 31218
rect 42642 31166 42654 31218
rect 41806 31154 41858 31166
rect 44494 31154 44546 31166
rect 44942 31218 44994 31230
rect 44942 31154 44994 31166
rect 45838 31218 45890 31230
rect 45838 31154 45890 31166
rect 8206 31106 8258 31118
rect 5618 31054 5630 31106
rect 5682 31054 5694 31106
rect 8206 31042 8258 31054
rect 8430 31106 8482 31118
rect 21086 31106 21138 31118
rect 45950 31106 46002 31118
rect 14690 31054 14702 31106
rect 14754 31054 14766 31106
rect 19506 31054 19518 31106
rect 19570 31054 19582 31106
rect 22530 31054 22542 31106
rect 22594 31054 22606 31106
rect 26674 31054 26686 31106
rect 26738 31054 26750 31106
rect 27906 31054 27918 31106
rect 27970 31054 27982 31106
rect 29586 31054 29598 31106
rect 29650 31054 29662 31106
rect 33282 31054 33294 31106
rect 33346 31054 33358 31106
rect 42354 31054 42366 31106
rect 42418 31054 42430 31106
rect 43922 31054 43934 31106
rect 43986 31054 43998 31106
rect 8430 31042 8482 31054
rect 21086 31042 21138 31054
rect 45950 31042 46002 31054
rect 8542 30994 8594 31006
rect 7634 30942 7646 30994
rect 7698 30942 7710 30994
rect 8542 30930 8594 30942
rect 9102 30994 9154 31006
rect 9102 30930 9154 30942
rect 9886 30994 9938 31006
rect 41582 30994 41634 31006
rect 43486 30994 43538 31006
rect 13346 30942 13358 30994
rect 13410 30942 13422 30994
rect 14018 30942 14030 30994
rect 14082 30942 14094 30994
rect 20290 30942 20302 30994
rect 20354 30942 20366 30994
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 25218 30942 25230 30994
rect 25282 30942 25294 30994
rect 28354 30942 28366 30994
rect 28418 30942 28430 30994
rect 28914 30942 28926 30994
rect 28978 30942 28990 30994
rect 32386 30942 32398 30994
rect 32450 30942 32462 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 39778 30942 39790 30994
rect 39842 30942 39854 30994
rect 41346 30942 41358 30994
rect 41410 30942 41422 30994
rect 42018 30942 42030 30994
rect 42082 30942 42094 30994
rect 43026 30942 43038 30994
rect 43090 30942 43102 30994
rect 9886 30930 9938 30942
rect 41582 30930 41634 30942
rect 43486 30930 43538 30942
rect 20862 30882 20914 30894
rect 32174 30882 32226 30894
rect 40238 30882 40290 30894
rect 10434 30830 10446 30882
rect 10498 30830 10510 30882
rect 12562 30830 12574 30882
rect 12626 30830 12638 30882
rect 16818 30830 16830 30882
rect 16882 30830 16894 30882
rect 17378 30830 17390 30882
rect 17442 30830 17454 30882
rect 24658 30830 24670 30882
rect 24722 30830 24734 30882
rect 26562 30830 26574 30882
rect 26626 30830 26638 30882
rect 31714 30830 31726 30882
rect 31778 30830 31790 30882
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 20862 30818 20914 30830
rect 32174 30818 32226 30830
rect 40238 30818 40290 30830
rect 40910 30882 40962 30894
rect 40910 30818 40962 30830
rect 41694 30882 41746 30894
rect 41694 30818 41746 30830
rect 45390 30882 45442 30894
rect 45390 30818 45442 30830
rect 32062 30770 32114 30782
rect 32062 30706 32114 30718
rect 40126 30770 40178 30782
rect 40126 30706 40178 30718
rect 1344 30602 46592 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 46592 30602
rect 1344 30516 46592 30550
rect 12014 30434 12066 30446
rect 30818 30382 30830 30434
rect 30882 30382 30894 30434
rect 12014 30370 12066 30382
rect 19406 30322 19458 30334
rect 1698 30270 1710 30322
rect 1762 30270 1774 30322
rect 7410 30270 7422 30322
rect 7474 30270 7486 30322
rect 14018 30270 14030 30322
rect 14082 30270 14094 30322
rect 19406 30258 19458 30270
rect 26798 30322 26850 30334
rect 35186 30270 35198 30322
rect 35250 30270 35262 30322
rect 40450 30270 40462 30322
rect 40514 30270 40526 30322
rect 41570 30270 41582 30322
rect 41634 30270 41646 30322
rect 43698 30270 43710 30322
rect 43762 30270 43774 30322
rect 26798 30258 26850 30270
rect 5854 30210 5906 30222
rect 4610 30158 4622 30210
rect 4674 30158 4686 30210
rect 5854 30146 5906 30158
rect 6190 30210 6242 30222
rect 6190 30146 6242 30158
rect 6414 30210 6466 30222
rect 6414 30146 6466 30158
rect 7086 30210 7138 30222
rect 11230 30210 11282 30222
rect 10322 30158 10334 30210
rect 10386 30158 10398 30210
rect 7086 30146 7138 30158
rect 11230 30146 11282 30158
rect 11902 30210 11954 30222
rect 19294 30210 19346 30222
rect 17266 30158 17278 30210
rect 17330 30158 17342 30210
rect 19058 30158 19070 30210
rect 19122 30158 19134 30210
rect 11902 30146 11954 30158
rect 19294 30146 19346 30158
rect 20414 30210 20466 30222
rect 20414 30146 20466 30158
rect 21310 30210 21362 30222
rect 21310 30146 21362 30158
rect 21982 30210 22034 30222
rect 21982 30146 22034 30158
rect 22766 30210 22818 30222
rect 22766 30146 22818 30158
rect 22990 30210 23042 30222
rect 22990 30146 23042 30158
rect 23326 30210 23378 30222
rect 23326 30146 23378 30158
rect 23886 30210 23938 30222
rect 23886 30146 23938 30158
rect 24558 30210 24610 30222
rect 24558 30146 24610 30158
rect 25902 30210 25954 30222
rect 25902 30146 25954 30158
rect 26686 30210 26738 30222
rect 26686 30146 26738 30158
rect 27246 30210 27298 30222
rect 27246 30146 27298 30158
rect 27582 30210 27634 30222
rect 27582 30146 27634 30158
rect 27806 30210 27858 30222
rect 30158 30210 30210 30222
rect 28466 30158 28478 30210
rect 28530 30158 28542 30210
rect 27806 30146 27858 30158
rect 30158 30146 30210 30158
rect 31838 30210 31890 30222
rect 31838 30146 31890 30158
rect 32398 30210 32450 30222
rect 32398 30146 32450 30158
rect 33742 30210 33794 30222
rect 33742 30146 33794 30158
rect 34302 30210 34354 30222
rect 44046 30210 44098 30222
rect 34850 30158 34862 30210
rect 34914 30158 34926 30210
rect 37538 30158 37550 30210
rect 37602 30158 37614 30210
rect 38322 30158 38334 30210
rect 38386 30158 38398 30210
rect 40786 30158 40798 30210
rect 40850 30158 40862 30210
rect 34302 30146 34354 30158
rect 44046 30146 44098 30158
rect 44942 30210 44994 30222
rect 44942 30146 44994 30158
rect 45390 30210 45442 30222
rect 45390 30146 45442 30158
rect 46174 30210 46226 30222
rect 46174 30146 46226 30158
rect 5630 30098 5682 30110
rect 3826 30046 3838 30098
rect 3890 30046 3902 30098
rect 5630 30034 5682 30046
rect 5742 30098 5794 30110
rect 5742 30034 5794 30046
rect 6862 30098 6914 30110
rect 25230 30098 25282 30110
rect 9538 30046 9550 30098
rect 9602 30046 9614 30098
rect 24882 30046 24894 30098
rect 24946 30046 24958 30098
rect 6862 30034 6914 30046
rect 25230 30034 25282 30046
rect 25454 30098 25506 30110
rect 25454 30034 25506 30046
rect 28142 30098 28194 30110
rect 28142 30034 28194 30046
rect 29598 30098 29650 30110
rect 29598 30034 29650 30046
rect 30270 30098 30322 30110
rect 30270 30034 30322 30046
rect 30382 30098 30434 30110
rect 30382 30034 30434 30046
rect 35758 30098 35810 30110
rect 35758 30034 35810 30046
rect 36094 30098 36146 30110
rect 36094 30034 36146 30046
rect 44158 30098 44210 30110
rect 44158 30034 44210 30046
rect 45838 30098 45890 30110
rect 45838 30034 45890 30046
rect 6638 29986 6690 29998
rect 6638 29922 6690 29934
rect 10670 29986 10722 29998
rect 10670 29922 10722 29934
rect 12462 29986 12514 29998
rect 12462 29922 12514 29934
rect 19518 29986 19570 29998
rect 19518 29922 19570 29934
rect 19630 29986 19682 29998
rect 21422 29986 21474 29998
rect 20066 29934 20078 29986
rect 20130 29934 20142 29986
rect 19630 29922 19682 29934
rect 21422 29922 21474 29934
rect 21534 29986 21586 29998
rect 25678 29986 25730 29998
rect 22418 29934 22430 29986
rect 22482 29934 22494 29986
rect 21534 29922 21586 29934
rect 25678 29922 25730 29934
rect 26462 29986 26514 29998
rect 26462 29922 26514 29934
rect 26910 29986 26962 29998
rect 26910 29922 26962 29934
rect 27694 29986 27746 29998
rect 27694 29922 27746 29934
rect 28254 29986 28306 29998
rect 28254 29922 28306 29934
rect 29486 29986 29538 29998
rect 29486 29922 29538 29934
rect 31278 29986 31330 29998
rect 31278 29922 31330 29934
rect 32958 29986 33010 29998
rect 32958 29922 33010 29934
rect 33406 29986 33458 29998
rect 33406 29922 33458 29934
rect 35646 29986 35698 29998
rect 37214 29986 37266 29998
rect 36418 29934 36430 29986
rect 36482 29934 36494 29986
rect 35646 29922 35698 29934
rect 37214 29922 37266 29934
rect 1344 29818 46592 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 46592 29818
rect 1344 29732 46592 29766
rect 3166 29650 3218 29662
rect 3166 29586 3218 29598
rect 8094 29650 8146 29662
rect 8094 29586 8146 29598
rect 8654 29650 8706 29662
rect 8654 29586 8706 29598
rect 16382 29650 16434 29662
rect 16382 29586 16434 29598
rect 17614 29650 17666 29662
rect 17614 29586 17666 29598
rect 17726 29650 17778 29662
rect 17726 29586 17778 29598
rect 17838 29650 17890 29662
rect 17838 29586 17890 29598
rect 17950 29650 18002 29662
rect 17950 29586 18002 29598
rect 18510 29650 18562 29662
rect 23662 29650 23714 29662
rect 23202 29598 23214 29650
rect 23266 29598 23278 29650
rect 18510 29586 18562 29598
rect 23662 29586 23714 29598
rect 24558 29650 24610 29662
rect 24558 29586 24610 29598
rect 24670 29650 24722 29662
rect 33182 29650 33234 29662
rect 31378 29598 31390 29650
rect 31442 29598 31454 29650
rect 24670 29586 24722 29598
rect 33182 29586 33234 29598
rect 33406 29650 33458 29662
rect 33406 29586 33458 29598
rect 33518 29650 33570 29662
rect 33518 29586 33570 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 2606 29538 2658 29550
rect 7422 29538 7474 29550
rect 4386 29486 4398 29538
rect 4450 29486 4462 29538
rect 2606 29474 2658 29486
rect 7422 29474 7474 29486
rect 7870 29538 7922 29550
rect 7870 29474 7922 29486
rect 8430 29538 8482 29550
rect 8430 29474 8482 29486
rect 8878 29538 8930 29550
rect 8878 29474 8930 29486
rect 14142 29538 14194 29550
rect 14142 29474 14194 29486
rect 17390 29538 17442 29550
rect 23774 29538 23826 29550
rect 20962 29486 20974 29538
rect 21026 29486 21038 29538
rect 36082 29486 36094 29538
rect 36146 29486 36158 29538
rect 43810 29486 43822 29538
rect 43874 29486 43886 29538
rect 17390 29474 17442 29486
rect 23774 29474 23826 29486
rect 2158 29426 2210 29438
rect 2158 29362 2210 29374
rect 2494 29426 2546 29438
rect 2494 29362 2546 29374
rect 2830 29426 2882 29438
rect 2830 29362 2882 29374
rect 3054 29426 3106 29438
rect 7310 29426 7362 29438
rect 3714 29374 3726 29426
rect 3778 29374 3790 29426
rect 3054 29362 3106 29374
rect 7310 29362 7362 29374
rect 7646 29426 7698 29438
rect 7646 29362 7698 29374
rect 8094 29426 8146 29438
rect 8094 29362 8146 29374
rect 8990 29426 9042 29438
rect 14478 29426 14530 29438
rect 10882 29374 10894 29426
rect 10946 29374 10958 29426
rect 8990 29362 9042 29374
rect 14478 29362 14530 29374
rect 14926 29426 14978 29438
rect 22430 29426 22482 29438
rect 15362 29374 15374 29426
rect 15426 29374 15438 29426
rect 21634 29374 21646 29426
rect 21698 29374 21710 29426
rect 14926 29362 14978 29374
rect 22430 29362 22482 29374
rect 22878 29426 22930 29438
rect 22878 29362 22930 29374
rect 23998 29426 24050 29438
rect 23998 29362 24050 29374
rect 24446 29426 24498 29438
rect 31054 29426 31106 29438
rect 30482 29374 30494 29426
rect 30546 29374 30558 29426
rect 24446 29362 24498 29374
rect 31054 29362 31106 29374
rect 32286 29426 32338 29438
rect 32286 29362 32338 29374
rect 33294 29426 33346 29438
rect 39790 29426 39842 29438
rect 33730 29374 33742 29426
rect 33794 29374 33806 29426
rect 34066 29374 34078 29426
rect 34130 29374 34142 29426
rect 33294 29362 33346 29374
rect 39790 29362 39842 29374
rect 39902 29426 39954 29438
rect 39902 29362 39954 29374
rect 40014 29426 40066 29438
rect 40014 29362 40066 29374
rect 40126 29426 40178 29438
rect 40338 29374 40350 29426
rect 40402 29374 40414 29426
rect 42242 29374 42254 29426
rect 42306 29374 42318 29426
rect 40126 29362 40178 29374
rect 15822 29314 15874 29326
rect 6514 29262 6526 29314
rect 6578 29262 6590 29314
rect 11554 29262 11566 29314
rect 11618 29262 11630 29314
rect 13682 29262 13694 29314
rect 13746 29262 13758 29314
rect 15822 29250 15874 29262
rect 16942 29314 16994 29326
rect 22654 29314 22706 29326
rect 30830 29314 30882 29326
rect 18834 29262 18846 29314
rect 18898 29262 18910 29314
rect 25554 29262 25566 29314
rect 25618 29262 25630 29314
rect 31826 29262 31838 29314
rect 31890 29262 31902 29314
rect 16942 29250 16994 29262
rect 22654 29250 22706 29262
rect 30830 29250 30882 29262
rect 2046 29202 2098 29214
rect 2046 29138 2098 29150
rect 3166 29202 3218 29214
rect 3166 29138 3218 29150
rect 23662 29202 23714 29214
rect 23662 29138 23714 29150
rect 1344 29034 46592 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 46592 29034
rect 1344 28948 46592 28982
rect 6862 28866 6914 28878
rect 6862 28802 6914 28814
rect 25454 28866 25506 28878
rect 25454 28802 25506 28814
rect 26910 28866 26962 28878
rect 26910 28802 26962 28814
rect 6638 28754 6690 28766
rect 11118 28754 11170 28766
rect 1698 28702 1710 28754
rect 1762 28702 1774 28754
rect 7410 28702 7422 28754
rect 7474 28702 7486 28754
rect 6638 28690 6690 28702
rect 11118 28690 11170 28702
rect 13022 28754 13074 28766
rect 21646 28754 21698 28766
rect 25342 28754 25394 28766
rect 44942 28754 44994 28766
rect 20178 28702 20190 28754
rect 20242 28702 20254 28754
rect 22754 28702 22766 28754
rect 22818 28702 22830 28754
rect 24882 28702 24894 28754
rect 24946 28702 24958 28754
rect 28466 28702 28478 28754
rect 28530 28702 28542 28754
rect 29922 28702 29934 28754
rect 29986 28702 29998 28754
rect 32050 28702 32062 28754
rect 32114 28702 32126 28754
rect 33170 28702 33182 28754
rect 33234 28702 33246 28754
rect 35298 28702 35310 28754
rect 35362 28702 35374 28754
rect 36978 28702 36990 28754
rect 37042 28702 37054 28754
rect 40898 28702 40910 28754
rect 40962 28702 40974 28754
rect 41346 28702 41358 28754
rect 41410 28702 41422 28754
rect 13022 28690 13074 28702
rect 21646 28690 21698 28702
rect 25342 28690 25394 28702
rect 44942 28690 44994 28702
rect 45390 28754 45442 28766
rect 45390 28690 45442 28702
rect 6414 28642 6466 28654
rect 4610 28590 4622 28642
rect 4674 28590 4686 28642
rect 6414 28578 6466 28590
rect 6974 28642 7026 28654
rect 10782 28642 10834 28654
rect 9538 28590 9550 28642
rect 9602 28590 9614 28642
rect 10322 28590 10334 28642
rect 10386 28590 10398 28642
rect 6974 28578 7026 28590
rect 10782 28578 10834 28590
rect 11006 28642 11058 28654
rect 11006 28578 11058 28590
rect 11342 28642 11394 28654
rect 11342 28578 11394 28590
rect 12238 28642 12290 28654
rect 26126 28642 26178 28654
rect 19618 28590 19630 28642
rect 19682 28590 19694 28642
rect 20626 28590 20638 28642
rect 20690 28590 20702 28642
rect 21970 28590 21982 28642
rect 22034 28590 22046 28642
rect 12238 28578 12290 28590
rect 26126 28578 26178 28590
rect 26462 28642 26514 28654
rect 26462 28578 26514 28590
rect 26686 28642 26738 28654
rect 26686 28578 26738 28590
rect 27806 28642 27858 28654
rect 27806 28578 27858 28590
rect 28142 28642 28194 28654
rect 44830 28642 44882 28654
rect 29138 28590 29150 28642
rect 29202 28590 29214 28642
rect 32722 28590 32734 28642
rect 32786 28590 32798 28642
rect 35970 28590 35982 28642
rect 36034 28590 36046 28642
rect 39106 28590 39118 28642
rect 39170 28590 39182 28642
rect 39890 28590 39902 28642
rect 39954 28590 39966 28642
rect 40338 28590 40350 28642
rect 40402 28590 40414 28642
rect 41010 28590 41022 28642
rect 41074 28590 41086 28642
rect 43474 28590 43486 28642
rect 43538 28590 43550 28642
rect 44146 28590 44158 28642
rect 44210 28590 44222 28642
rect 28142 28578 28194 28590
rect 44830 28578 44882 28590
rect 45838 28642 45890 28654
rect 45838 28578 45890 28590
rect 11678 28530 11730 28542
rect 25790 28530 25842 28542
rect 3826 28478 3838 28530
rect 3890 28478 3902 28530
rect 5618 28478 5630 28530
rect 5682 28478 5694 28530
rect 16370 28478 16382 28530
rect 16434 28478 16446 28530
rect 11678 28466 11730 28478
rect 25790 28466 25842 28478
rect 32398 28530 32450 28542
rect 32398 28466 32450 28478
rect 40798 28530 40850 28542
rect 40798 28466 40850 28478
rect 5966 28418 6018 28430
rect 5966 28354 6018 28366
rect 6526 28418 6578 28430
rect 6526 28354 6578 28366
rect 11566 28418 11618 28430
rect 11566 28354 11618 28366
rect 11790 28418 11842 28430
rect 13806 28418 13858 28430
rect 13458 28366 13470 28418
rect 13522 28366 13534 28418
rect 11790 28354 11842 28366
rect 13806 28354 13858 28366
rect 20078 28418 20130 28430
rect 20078 28354 20130 28366
rect 20190 28418 20242 28430
rect 20190 28354 20242 28366
rect 20414 28418 20466 28430
rect 20414 28354 20466 28366
rect 26238 28418 26290 28430
rect 32510 28418 32562 28430
rect 27234 28366 27246 28418
rect 27298 28366 27310 28418
rect 26238 28354 26290 28366
rect 32510 28354 32562 28366
rect 40574 28418 40626 28430
rect 40574 28354 40626 28366
rect 1344 28250 46592 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 46592 28250
rect 1344 28164 46592 28198
rect 3838 28082 3890 28094
rect 3838 28018 3890 28030
rect 5742 28082 5794 28094
rect 5742 28018 5794 28030
rect 6302 28082 6354 28094
rect 6302 28018 6354 28030
rect 7198 28082 7250 28094
rect 7198 28018 7250 28030
rect 7422 28082 7474 28094
rect 7422 28018 7474 28030
rect 7758 28082 7810 28094
rect 7758 28018 7810 28030
rect 8318 28082 8370 28094
rect 8318 28018 8370 28030
rect 9662 28082 9714 28094
rect 9662 28018 9714 28030
rect 10446 28082 10498 28094
rect 10446 28018 10498 28030
rect 11790 28082 11842 28094
rect 11790 28018 11842 28030
rect 18846 28082 18898 28094
rect 18846 28018 18898 28030
rect 23214 28082 23266 28094
rect 23214 28018 23266 28030
rect 24558 28082 24610 28094
rect 24558 28018 24610 28030
rect 24670 28082 24722 28094
rect 31614 28082 31666 28094
rect 26786 28030 26798 28082
rect 26850 28030 26862 28082
rect 27234 28030 27246 28082
rect 27298 28030 27310 28082
rect 24670 28018 24722 28030
rect 31614 28018 31666 28030
rect 31950 28082 32002 28094
rect 31950 28018 32002 28030
rect 32062 28082 32114 28094
rect 32062 28018 32114 28030
rect 32286 28082 32338 28094
rect 32286 28018 32338 28030
rect 39566 28082 39618 28094
rect 39566 28018 39618 28030
rect 3166 27970 3218 27982
rect 3166 27906 3218 27918
rect 5294 27970 5346 27982
rect 5294 27906 5346 27918
rect 6414 27970 6466 27982
rect 6414 27906 6466 27918
rect 8766 27970 8818 27982
rect 17838 27970 17890 27982
rect 12114 27918 12126 27970
rect 12178 27918 12190 27970
rect 14690 27918 14702 27970
rect 14754 27918 14766 27970
rect 8766 27906 8818 27918
rect 17838 27906 17890 27918
rect 17950 27970 18002 27982
rect 17950 27906 18002 27918
rect 19518 27970 19570 27982
rect 19518 27906 19570 27918
rect 28254 27970 28306 27982
rect 28254 27906 28306 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 38334 27970 38386 27982
rect 38334 27906 38386 27918
rect 38894 27970 38946 27982
rect 41234 27918 41246 27970
rect 41298 27918 41310 27970
rect 38894 27906 38946 27918
rect 3054 27858 3106 27870
rect 3054 27794 3106 27806
rect 3502 27858 3554 27870
rect 3502 27794 3554 27806
rect 3950 27858 4002 27870
rect 3950 27794 4002 27806
rect 4174 27858 4226 27870
rect 4174 27794 4226 27806
rect 4622 27858 4674 27870
rect 4622 27794 4674 27806
rect 4958 27858 5010 27870
rect 4958 27794 5010 27806
rect 5182 27858 5234 27870
rect 5182 27794 5234 27806
rect 5518 27858 5570 27870
rect 5518 27794 5570 27806
rect 5854 27858 5906 27870
rect 5854 27794 5906 27806
rect 7086 27858 7138 27870
rect 7086 27794 7138 27806
rect 7646 27858 7698 27870
rect 7646 27794 7698 27806
rect 7982 27858 8034 27870
rect 7982 27794 8034 27806
rect 8094 27858 8146 27870
rect 8094 27794 8146 27806
rect 8542 27858 8594 27870
rect 8542 27794 8594 27806
rect 12462 27858 12514 27870
rect 12462 27794 12514 27806
rect 13246 27858 13298 27870
rect 13246 27794 13298 27806
rect 13358 27858 13410 27870
rect 18622 27858 18674 27870
rect 22990 27858 23042 27870
rect 13570 27806 13582 27858
rect 13634 27806 13646 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 18386 27806 18398 27858
rect 18450 27806 18462 27858
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 22642 27806 22654 27858
rect 22706 27806 22718 27858
rect 13358 27794 13410 27806
rect 18622 27794 18674 27806
rect 22990 27794 23042 27806
rect 23326 27858 23378 27870
rect 23326 27794 23378 27806
rect 23662 27858 23714 27870
rect 23662 27794 23714 27806
rect 23998 27858 24050 27870
rect 23998 27794 24050 27806
rect 24446 27858 24498 27870
rect 26350 27858 26402 27870
rect 37662 27858 37714 27870
rect 26114 27806 26126 27858
rect 26178 27806 26190 27858
rect 28690 27806 28702 27858
rect 28754 27806 28766 27858
rect 30930 27806 30942 27858
rect 30994 27806 31006 27858
rect 32498 27806 32510 27858
rect 32562 27806 32574 27858
rect 33170 27806 33182 27858
rect 33234 27806 33246 27858
rect 37314 27806 37326 27858
rect 37378 27806 37390 27858
rect 24446 27794 24498 27806
rect 26350 27794 26402 27806
rect 37662 27794 37714 27806
rect 38782 27858 38834 27870
rect 38782 27794 38834 27806
rect 39454 27858 39506 27870
rect 39454 27794 39506 27806
rect 39790 27858 39842 27870
rect 39790 27794 39842 27806
rect 39902 27858 39954 27870
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 42130 27806 42142 27858
rect 42194 27806 42206 27858
rect 46050 27806 46062 27858
rect 46114 27806 46126 27858
rect 39902 27794 39954 27806
rect 10334 27746 10386 27758
rect 17502 27746 17554 27758
rect 16818 27694 16830 27746
rect 16882 27694 16894 27746
rect 10334 27682 10386 27694
rect 17502 27682 17554 27694
rect 18734 27746 18786 27758
rect 32174 27746 32226 27758
rect 36430 27746 36482 27758
rect 19842 27694 19854 27746
rect 19906 27694 19918 27746
rect 21970 27694 21982 27746
rect 22034 27694 22046 27746
rect 26002 27694 26014 27746
rect 26066 27694 26078 27746
rect 33842 27694 33854 27746
rect 33906 27694 33918 27746
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 18734 27682 18786 27694
rect 32174 27682 32226 27694
rect 36430 27682 36482 27694
rect 37774 27746 37826 27758
rect 37774 27682 37826 27694
rect 38110 27746 38162 27758
rect 39678 27746 39730 27758
rect 42702 27746 42754 27758
rect 38322 27694 38334 27746
rect 38386 27694 38398 27746
rect 41906 27694 41918 27746
rect 41970 27694 41982 27746
rect 43250 27694 43262 27746
rect 43314 27694 43326 27746
rect 45378 27694 45390 27746
rect 45442 27694 45454 27746
rect 38110 27682 38162 27694
rect 39678 27682 39730 27694
rect 42702 27682 42754 27694
rect 3166 27634 3218 27646
rect 3166 27570 3218 27582
rect 4734 27634 4786 27646
rect 4734 27570 4786 27582
rect 6302 27634 6354 27646
rect 6302 27570 6354 27582
rect 10222 27634 10274 27646
rect 17390 27634 17442 27646
rect 12786 27582 12798 27634
rect 12850 27582 12862 27634
rect 10222 27570 10274 27582
rect 17390 27570 17442 27582
rect 1344 27466 46592 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 46592 27466
rect 1344 27380 46592 27414
rect 27582 27298 27634 27310
rect 13794 27246 13806 27298
rect 13858 27295 13870 27298
rect 14130 27295 14142 27298
rect 13858 27249 14142 27295
rect 13858 27246 13870 27249
rect 14130 27246 14142 27249
rect 14194 27246 14206 27298
rect 27582 27234 27634 27246
rect 27918 27298 27970 27310
rect 27918 27234 27970 27246
rect 28254 27298 28306 27310
rect 28254 27234 28306 27246
rect 29486 27298 29538 27310
rect 30382 27298 30434 27310
rect 33294 27298 33346 27310
rect 29810 27246 29822 27298
rect 29874 27246 29886 27298
rect 30706 27246 30718 27298
rect 30770 27246 30782 27298
rect 29486 27234 29538 27246
rect 30382 27234 30434 27246
rect 33294 27234 33346 27246
rect 38894 27298 38946 27310
rect 38894 27234 38946 27246
rect 39902 27298 39954 27310
rect 39902 27234 39954 27246
rect 40462 27298 40514 27310
rect 40462 27234 40514 27246
rect 44718 27298 44770 27310
rect 44718 27234 44770 27246
rect 29262 27186 29314 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 12226 27134 12238 27186
rect 12290 27134 12302 27186
rect 13906 27134 13918 27186
rect 13970 27134 13982 27186
rect 16258 27134 16270 27186
rect 16322 27134 16334 27186
rect 18386 27134 18398 27186
rect 18450 27134 18462 27186
rect 19058 27134 19070 27186
rect 19122 27134 19134 27186
rect 19730 27134 19742 27186
rect 19794 27134 19806 27186
rect 24210 27134 24222 27186
rect 24274 27134 24286 27186
rect 29262 27122 29314 27134
rect 30158 27186 30210 27198
rect 30158 27122 30210 27134
rect 31614 27186 31666 27198
rect 31614 27122 31666 27134
rect 32510 27186 32562 27198
rect 32510 27122 32562 27134
rect 33182 27186 33234 27198
rect 33182 27122 33234 27134
rect 34190 27186 34242 27198
rect 35982 27186 36034 27198
rect 35298 27134 35310 27186
rect 35362 27134 35374 27186
rect 34190 27122 34242 27134
rect 35982 27122 36034 27134
rect 37886 27186 37938 27198
rect 37886 27122 37938 27134
rect 38446 27186 38498 27198
rect 38446 27122 38498 27134
rect 38782 27186 38834 27198
rect 43822 27186 43874 27198
rect 42578 27134 42590 27186
rect 42642 27134 42654 27186
rect 38782 27122 38834 27134
rect 43822 27122 43874 27134
rect 14142 27074 14194 27086
rect 24782 27074 24834 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 7074 27022 7086 27074
rect 7138 27022 7150 27074
rect 9426 27022 9438 27074
rect 9490 27022 9502 27074
rect 14242 27022 14254 27074
rect 14306 27022 14318 27074
rect 15474 27022 15486 27074
rect 15538 27022 15550 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 20066 27022 20078 27074
rect 20130 27022 20142 27074
rect 21410 27022 21422 27074
rect 21474 27022 21486 27074
rect 14142 27010 14194 27022
rect 24782 27010 24834 27022
rect 26462 27074 26514 27086
rect 26462 27010 26514 27022
rect 28366 27074 28418 27086
rect 28366 27010 28418 27022
rect 33742 27074 33794 27086
rect 33742 27010 33794 27022
rect 34862 27074 34914 27086
rect 34862 27010 34914 27022
rect 37102 27074 37154 27086
rect 37102 27010 37154 27022
rect 39230 27074 39282 27086
rect 39230 27010 39282 27022
rect 40014 27074 40066 27086
rect 41022 27074 41074 27086
rect 40786 27022 40798 27074
rect 40850 27022 40862 27074
rect 40014 27010 40066 27022
rect 41022 27010 41074 27022
rect 41246 27074 41298 27086
rect 41246 27010 41298 27022
rect 41358 27074 41410 27086
rect 42926 27074 42978 27086
rect 44046 27074 44098 27086
rect 45614 27074 45666 27086
rect 42466 27022 42478 27074
rect 42530 27022 42542 27074
rect 43138 27022 43150 27074
rect 43202 27022 43214 27074
rect 45042 27022 45054 27074
rect 45106 27022 45118 27074
rect 46050 27022 46062 27074
rect 46114 27022 46126 27074
rect 41358 27010 41410 27022
rect 42926 27010 42978 27022
rect 44046 27010 44098 27022
rect 45614 27010 45666 27022
rect 25678 26962 25730 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 10098 26910 10110 26962
rect 10162 26910 10174 26962
rect 19618 26910 19630 26962
rect 19682 26910 19694 26962
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 25678 26898 25730 26910
rect 27694 26962 27746 26974
rect 27694 26898 27746 26910
rect 31166 26962 31218 26974
rect 40350 26962 40402 26974
rect 37426 26910 37438 26962
rect 37490 26910 37502 26962
rect 41918 26962 41970 26974
rect 31166 26898 31218 26910
rect 40350 26898 40402 26910
rect 41806 26906 41858 26918
rect 26126 26850 26178 26862
rect 6850 26798 6862 26850
rect 6914 26798 6926 26850
rect 13682 26798 13694 26850
rect 13746 26798 13758 26850
rect 26126 26786 26178 26798
rect 31054 26850 31106 26862
rect 31054 26786 31106 26798
rect 36094 26850 36146 26862
rect 36094 26786 36146 26798
rect 39566 26850 39618 26862
rect 39566 26786 39618 26798
rect 41134 26850 41186 26862
rect 41918 26898 41970 26910
rect 42702 26962 42754 26974
rect 42702 26898 42754 26910
rect 44830 26962 44882 26974
rect 44830 26898 44882 26910
rect 45278 26962 45330 26974
rect 45278 26898 45330 26910
rect 41806 26842 41858 26854
rect 42142 26850 42194 26862
rect 41134 26786 41186 26798
rect 43474 26798 43486 26850
rect 43538 26798 43550 26850
rect 42142 26786 42194 26798
rect 1344 26682 46592 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 46592 26682
rect 1344 26596 46592 26630
rect 3166 26514 3218 26526
rect 3166 26450 3218 26462
rect 3950 26514 4002 26526
rect 3950 26450 4002 26462
rect 4622 26514 4674 26526
rect 4622 26450 4674 26462
rect 10334 26514 10386 26526
rect 10334 26450 10386 26462
rect 17614 26514 17666 26526
rect 17614 26450 17666 26462
rect 22990 26514 23042 26526
rect 22990 26450 23042 26462
rect 24110 26514 24162 26526
rect 24110 26450 24162 26462
rect 24782 26514 24834 26526
rect 37774 26514 37826 26526
rect 39902 26514 39954 26526
rect 28466 26462 28478 26514
rect 28530 26462 28542 26514
rect 38434 26462 38446 26514
rect 38498 26462 38510 26514
rect 24782 26450 24834 26462
rect 37774 26450 37826 26462
rect 39902 26450 39954 26462
rect 40350 26514 40402 26526
rect 40350 26450 40402 26462
rect 3054 26402 3106 26414
rect 3054 26338 3106 26350
rect 3838 26402 3890 26414
rect 3838 26338 3890 26350
rect 4398 26402 4450 26414
rect 23662 26402 23714 26414
rect 39454 26402 39506 26414
rect 9874 26350 9886 26402
rect 9938 26350 9950 26402
rect 17938 26350 17950 26402
rect 18002 26350 18014 26402
rect 21186 26350 21198 26402
rect 21250 26350 21262 26402
rect 26226 26350 26238 26402
rect 26290 26350 26302 26402
rect 30258 26350 30270 26402
rect 30322 26350 30334 26402
rect 42242 26350 42254 26402
rect 42306 26350 42318 26402
rect 4398 26338 4450 26350
rect 23662 26338 23714 26350
rect 39454 26338 39506 26350
rect 3726 26290 3778 26302
rect 3726 26226 3778 26238
rect 4286 26290 4338 26302
rect 4286 26226 4338 26238
rect 4734 26290 4786 26302
rect 22878 26290 22930 26302
rect 5730 26238 5742 26290
rect 5794 26238 5806 26290
rect 9650 26238 9662 26290
rect 9714 26238 9726 26290
rect 10770 26238 10782 26290
rect 10834 26238 10846 26290
rect 13906 26238 13918 26290
rect 13970 26238 13982 26290
rect 18274 26238 18286 26290
rect 18338 26238 18350 26290
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 21746 26238 21758 26290
rect 21810 26238 21822 26290
rect 4734 26226 4786 26238
rect 22878 26226 22930 26238
rect 23102 26290 23154 26302
rect 23102 26226 23154 26238
rect 23550 26290 23602 26302
rect 36878 26290 36930 26302
rect 37550 26290 37602 26302
rect 38782 26290 38834 26302
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 29586 26238 29598 26290
rect 29650 26238 29662 26290
rect 33394 26238 33406 26290
rect 33458 26238 33470 26290
rect 37314 26238 37326 26290
rect 37378 26238 37390 26290
rect 37986 26238 37998 26290
rect 38050 26238 38062 26290
rect 45490 26238 45502 26290
rect 45554 26238 45566 26290
rect 23550 26226 23602 26238
rect 36878 26226 36930 26238
rect 37550 26226 37602 26238
rect 38782 26226 38834 26238
rect 20526 26178 20578 26190
rect 6402 26126 6414 26178
rect 6466 26126 6478 26178
rect 8530 26126 8542 26178
rect 8594 26126 8606 26178
rect 11442 26126 11454 26178
rect 11506 26126 11518 26178
rect 13570 26126 13582 26178
rect 13634 26126 13646 26178
rect 14690 26126 14702 26178
rect 14754 26126 14766 26178
rect 16818 26126 16830 26178
rect 16882 26126 16894 26178
rect 20526 26114 20578 26126
rect 22654 26178 22706 26190
rect 36766 26178 36818 26190
rect 32386 26126 32398 26178
rect 32450 26126 32462 26178
rect 34178 26126 34190 26178
rect 34242 26126 34254 26178
rect 36306 26126 36318 26178
rect 36370 26126 36382 26178
rect 22654 26114 22706 26126
rect 36766 26114 36818 26126
rect 37662 26178 37714 26190
rect 37662 26114 37714 26126
rect 40238 26178 40290 26190
rect 40238 26114 40290 26126
rect 3166 26066 3218 26078
rect 3166 26002 3218 26014
rect 22430 26066 22482 26078
rect 22430 26002 22482 26014
rect 39342 26066 39394 26078
rect 39342 26002 39394 26014
rect 1344 25898 46592 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 46592 25898
rect 1344 25812 46592 25846
rect 6414 25730 6466 25742
rect 6414 25666 6466 25678
rect 21422 25730 21474 25742
rect 21422 25666 21474 25678
rect 29486 25730 29538 25742
rect 29486 25666 29538 25678
rect 35982 25730 36034 25742
rect 35982 25666 36034 25678
rect 36318 25730 36370 25742
rect 36318 25666 36370 25678
rect 37326 25730 37378 25742
rect 37326 25666 37378 25678
rect 44830 25730 44882 25742
rect 44830 25666 44882 25678
rect 45166 25730 45218 25742
rect 45166 25666 45218 25678
rect 12798 25618 12850 25630
rect 1698 25566 1710 25618
rect 1762 25566 1774 25618
rect 12798 25554 12850 25566
rect 17502 25618 17554 25630
rect 17502 25554 17554 25566
rect 19294 25618 19346 25630
rect 19294 25554 19346 25566
rect 20414 25618 20466 25630
rect 20414 25554 20466 25566
rect 21310 25618 21362 25630
rect 29710 25618 29762 25630
rect 24658 25566 24670 25618
rect 24722 25566 24734 25618
rect 21310 25554 21362 25566
rect 29710 25554 29762 25566
rect 30718 25618 30770 25630
rect 33182 25618 33234 25630
rect 31154 25566 31166 25618
rect 31218 25566 31230 25618
rect 32162 25566 32174 25618
rect 32226 25566 32238 25618
rect 30718 25554 30770 25566
rect 33182 25554 33234 25566
rect 35310 25618 35362 25630
rect 35310 25554 35362 25566
rect 37102 25618 37154 25630
rect 37102 25554 37154 25566
rect 40798 25618 40850 25630
rect 40798 25554 40850 25566
rect 45614 25618 45666 25630
rect 45614 25554 45666 25566
rect 46174 25618 46226 25630
rect 46174 25554 46226 25566
rect 18062 25506 18114 25518
rect 4498 25454 4510 25506
rect 4562 25454 4574 25506
rect 5842 25454 5854 25506
rect 5906 25454 5918 25506
rect 8306 25454 8318 25506
rect 8370 25454 8382 25506
rect 13570 25454 13582 25506
rect 13634 25454 13646 25506
rect 18062 25442 18114 25454
rect 18398 25506 18450 25518
rect 18398 25442 18450 25454
rect 18510 25506 18562 25518
rect 18510 25442 18562 25454
rect 18734 25506 18786 25518
rect 19406 25506 19458 25518
rect 18946 25454 18958 25506
rect 19010 25454 19022 25506
rect 18734 25442 18786 25454
rect 19406 25442 19458 25454
rect 19854 25506 19906 25518
rect 19854 25442 19906 25454
rect 20078 25506 20130 25518
rect 20078 25442 20130 25454
rect 20302 25506 20354 25518
rect 25118 25506 25170 25518
rect 21858 25454 21870 25506
rect 21922 25454 21934 25506
rect 20302 25442 20354 25454
rect 25118 25442 25170 25454
rect 25230 25506 25282 25518
rect 31278 25506 31330 25518
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 25230 25442 25282 25454
rect 31278 25442 31330 25454
rect 31502 25506 31554 25518
rect 32510 25506 32562 25518
rect 36206 25506 36258 25518
rect 32050 25454 32062 25506
rect 32114 25454 32126 25506
rect 32722 25454 32734 25506
rect 32786 25454 32798 25506
rect 35746 25454 35758 25506
rect 35810 25454 35822 25506
rect 31502 25442 31554 25454
rect 32510 25442 32562 25454
rect 36206 25442 36258 25454
rect 38558 25506 38610 25518
rect 38558 25442 38610 25454
rect 38894 25506 38946 25518
rect 38894 25442 38946 25454
rect 39230 25506 39282 25518
rect 39230 25442 39282 25454
rect 39678 25506 39730 25518
rect 39678 25442 39730 25454
rect 41470 25506 41522 25518
rect 41470 25442 41522 25454
rect 41582 25506 41634 25518
rect 41582 25442 41634 25454
rect 41694 25506 41746 25518
rect 46062 25506 46114 25518
rect 42018 25454 42030 25506
rect 42082 25454 42094 25506
rect 43250 25454 43262 25506
rect 43314 25454 43326 25506
rect 44258 25454 44270 25506
rect 44322 25454 44334 25506
rect 41694 25442 41746 25454
rect 46062 25442 46114 25454
rect 6750 25394 6802 25406
rect 25454 25394 25506 25406
rect 3826 25342 3838 25394
rect 3890 25342 3902 25394
rect 5618 25342 5630 25394
rect 5682 25342 5694 25394
rect 10994 25342 11006 25394
rect 11058 25342 11070 25394
rect 14242 25342 14254 25394
rect 14306 25342 14318 25394
rect 22530 25342 22542 25394
rect 22594 25342 22606 25394
rect 6750 25330 6802 25342
rect 25454 25330 25506 25342
rect 25566 25394 25618 25406
rect 26798 25394 26850 25406
rect 26002 25342 26014 25394
rect 26066 25342 26078 25394
rect 25566 25330 25618 25342
rect 26798 25330 26850 25342
rect 27134 25394 27186 25406
rect 27134 25330 27186 25342
rect 30606 25394 30658 25406
rect 30606 25330 30658 25342
rect 31166 25394 31218 25406
rect 31166 25330 31218 25342
rect 31726 25394 31778 25406
rect 31726 25330 31778 25342
rect 35422 25394 35474 25406
rect 35422 25330 35474 25342
rect 40126 25394 40178 25406
rect 40126 25330 40178 25342
rect 40350 25394 40402 25406
rect 42802 25342 42814 25394
rect 42866 25342 42878 25394
rect 40350 25330 40402 25342
rect 6526 25282 6578 25294
rect 18622 25282 18674 25294
rect 16482 25230 16494 25282
rect 16546 25230 16558 25282
rect 6526 25218 6578 25230
rect 18622 25218 18674 25230
rect 20526 25282 20578 25294
rect 20526 25218 20578 25230
rect 25342 25282 25394 25294
rect 25342 25218 25394 25230
rect 27246 25282 27298 25294
rect 32286 25282 32338 25294
rect 29138 25230 29150 25282
rect 29202 25230 29214 25282
rect 27246 25218 27298 25230
rect 32286 25218 32338 25230
rect 33630 25282 33682 25294
rect 33630 25218 33682 25230
rect 35198 25282 35250 25294
rect 38334 25282 38386 25294
rect 37650 25230 37662 25282
rect 37714 25230 37726 25282
rect 35198 25218 35250 25230
rect 38334 25218 38386 25230
rect 38894 25282 38946 25294
rect 38894 25218 38946 25230
rect 39902 25282 39954 25294
rect 39902 25218 39954 25230
rect 40686 25282 40738 25294
rect 40686 25218 40738 25230
rect 42366 25282 42418 25294
rect 45054 25282 45106 25294
rect 43138 25230 43150 25282
rect 43202 25230 43214 25282
rect 44146 25230 44158 25282
rect 44210 25230 44222 25282
rect 42366 25218 42418 25230
rect 45054 25218 45106 25230
rect 1344 25114 46592 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 46592 25114
rect 1344 25028 46592 25062
rect 3278 24946 3330 24958
rect 3278 24882 3330 24894
rect 3838 24946 3890 24958
rect 3838 24882 3890 24894
rect 5406 24946 5458 24958
rect 5406 24882 5458 24894
rect 7198 24946 7250 24958
rect 7198 24882 7250 24894
rect 7310 24946 7362 24958
rect 7310 24882 7362 24894
rect 7422 24946 7474 24958
rect 7422 24882 7474 24894
rect 9774 24946 9826 24958
rect 9774 24882 9826 24894
rect 23998 24946 24050 24958
rect 37550 24946 37602 24958
rect 25218 24894 25230 24946
rect 25282 24894 25294 24946
rect 23998 24882 24050 24894
rect 37550 24882 37602 24894
rect 38222 24946 38274 24958
rect 38222 24882 38274 24894
rect 5518 24834 5570 24846
rect 7982 24834 8034 24846
rect 4610 24782 4622 24834
rect 4674 24782 4686 24834
rect 6514 24782 6526 24834
rect 6578 24782 6590 24834
rect 5518 24770 5570 24782
rect 7982 24770 8034 24782
rect 8094 24834 8146 24846
rect 8094 24770 8146 24782
rect 8542 24834 8594 24846
rect 8542 24770 8594 24782
rect 8654 24834 8706 24846
rect 8654 24770 8706 24782
rect 16830 24834 16882 24846
rect 24110 24834 24162 24846
rect 34862 24834 34914 24846
rect 23314 24782 23326 24834
rect 23378 24782 23390 24834
rect 28354 24782 28366 24834
rect 28418 24782 28430 24834
rect 30370 24782 30382 24834
rect 30434 24782 30446 24834
rect 16830 24770 16882 24782
rect 24110 24770 24162 24782
rect 34862 24770 34914 24782
rect 36766 24834 36818 24846
rect 39902 24834 39954 24846
rect 36978 24782 36990 24834
rect 37042 24782 37054 24834
rect 36766 24770 36818 24782
rect 39902 24770 39954 24782
rect 40014 24834 40066 24846
rect 40014 24770 40066 24782
rect 41022 24834 41074 24846
rect 41022 24770 41074 24782
rect 41134 24834 41186 24846
rect 41134 24770 41186 24782
rect 41470 24834 41522 24846
rect 41470 24770 41522 24782
rect 3166 24722 3218 24734
rect 3166 24658 3218 24670
rect 3502 24722 3554 24734
rect 3502 24658 3554 24670
rect 3726 24722 3778 24734
rect 3726 24658 3778 24670
rect 3950 24722 4002 24734
rect 3950 24658 4002 24670
rect 4174 24722 4226 24734
rect 4174 24658 4226 24670
rect 4958 24722 5010 24734
rect 4958 24658 5010 24670
rect 6190 24722 6242 24734
rect 6190 24658 6242 24670
rect 6750 24722 6802 24734
rect 6750 24658 6802 24670
rect 8318 24722 8370 24734
rect 8318 24658 8370 24670
rect 8878 24722 8930 24734
rect 8878 24658 8930 24670
rect 9438 24722 9490 24734
rect 9438 24658 9490 24670
rect 9774 24722 9826 24734
rect 9774 24658 9826 24670
rect 10110 24722 10162 24734
rect 14478 24722 14530 24734
rect 10994 24670 11006 24722
rect 11058 24670 11070 24722
rect 10110 24658 10162 24670
rect 14478 24658 14530 24670
rect 14814 24722 14866 24734
rect 14814 24658 14866 24670
rect 15038 24722 15090 24734
rect 15038 24658 15090 24670
rect 16382 24722 16434 24734
rect 23662 24722 23714 24734
rect 17714 24670 17726 24722
rect 17778 24670 17790 24722
rect 16382 24658 16434 24670
rect 23662 24658 23714 24670
rect 25566 24722 25618 24734
rect 35422 24722 35474 24734
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 29698 24670 29710 24722
rect 29762 24670 29774 24722
rect 25566 24658 25618 24670
rect 35422 24658 35474 24670
rect 36654 24722 36706 24734
rect 37662 24722 37714 24734
rect 37090 24670 37102 24722
rect 37154 24670 37166 24722
rect 36654 24658 36706 24670
rect 37662 24658 37714 24670
rect 38110 24722 38162 24734
rect 38110 24658 38162 24670
rect 38334 24722 38386 24734
rect 38334 24658 38386 24670
rect 39454 24722 39506 24734
rect 39454 24658 39506 24670
rect 40238 24722 40290 24734
rect 40238 24658 40290 24670
rect 41582 24722 41634 24734
rect 42242 24670 42254 24722
rect 42306 24670 42318 24722
rect 43362 24670 43374 24722
rect 43426 24670 43438 24722
rect 41582 24658 41634 24670
rect 14702 24610 14754 24622
rect 24558 24610 24610 24622
rect 34190 24610 34242 24622
rect 39006 24610 39058 24622
rect 42926 24610 42978 24622
rect 11778 24558 11790 24610
rect 11842 24558 11854 24610
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 22306 24558 22318 24610
rect 22370 24558 22382 24610
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 32498 24558 32510 24610
rect 32562 24558 32574 24610
rect 34962 24558 34974 24610
rect 35026 24558 35038 24610
rect 42466 24558 42478 24610
rect 42530 24558 42542 24610
rect 44034 24558 44046 24610
rect 44098 24558 44110 24610
rect 46162 24558 46174 24610
rect 46226 24558 46238 24610
rect 14702 24546 14754 24558
rect 24558 24546 24610 24558
rect 34190 24546 34242 24558
rect 39006 24546 39058 24558
rect 42926 24546 42978 24558
rect 5406 24498 5458 24510
rect 5406 24434 5458 24446
rect 16718 24498 16770 24510
rect 16718 24434 16770 24446
rect 24446 24498 24498 24510
rect 24446 24434 24498 24446
rect 34302 24498 34354 24510
rect 34302 24434 34354 24446
rect 34638 24498 34690 24510
rect 34638 24434 34690 24446
rect 35534 24498 35586 24510
rect 35534 24434 35586 24446
rect 35758 24498 35810 24510
rect 35758 24434 35810 24446
rect 35870 24498 35922 24510
rect 35870 24434 35922 24446
rect 39230 24498 39282 24510
rect 39230 24434 39282 24446
rect 41022 24498 41074 24510
rect 41022 24434 41074 24446
rect 1344 24330 46592 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 46592 24330
rect 1344 24244 46592 24278
rect 12350 24162 12402 24174
rect 12350 24098 12402 24110
rect 12686 24162 12738 24174
rect 12686 24098 12738 24110
rect 29486 24162 29538 24174
rect 29486 24098 29538 24110
rect 30270 24162 30322 24174
rect 30270 24098 30322 24110
rect 40350 24162 40402 24174
rect 40350 24098 40402 24110
rect 43374 24162 43426 24174
rect 43374 24098 43426 24110
rect 43710 24162 43762 24174
rect 43710 24098 43762 24110
rect 44830 24162 44882 24174
rect 44830 24098 44882 24110
rect 46062 24162 46114 24174
rect 46062 24098 46114 24110
rect 7198 24050 7250 24062
rect 7198 23986 7250 23998
rect 7646 24050 7698 24062
rect 7646 23986 7698 23998
rect 7758 24050 7810 24062
rect 13918 24050 13970 24062
rect 8642 23998 8654 24050
rect 8706 23998 8718 24050
rect 7758 23986 7810 23998
rect 13918 23986 13970 23998
rect 14702 24050 14754 24062
rect 14702 23986 14754 23998
rect 14814 24050 14866 24062
rect 30046 24050 30098 24062
rect 39566 24050 39618 24062
rect 16370 23998 16382 24050
rect 16434 23998 16446 24050
rect 18498 23998 18510 24050
rect 18562 23998 18574 24050
rect 31826 23998 31838 24050
rect 31890 23998 31902 24050
rect 33954 23998 33966 24050
rect 34018 23998 34030 24050
rect 34402 23998 34414 24050
rect 34466 23998 34478 24050
rect 14814 23986 14866 23998
rect 30046 23986 30098 23998
rect 39566 23986 39618 23998
rect 40462 24050 40514 24062
rect 40462 23986 40514 23998
rect 40910 24050 40962 24062
rect 40910 23986 40962 23998
rect 41470 24050 41522 24062
rect 41470 23986 41522 23998
rect 42478 24050 42530 24062
rect 45838 24050 45890 24062
rect 45154 23998 45166 24050
rect 45218 23998 45230 24050
rect 42478 23986 42530 23998
rect 45838 23986 45890 23998
rect 46174 24050 46226 24062
rect 46174 23986 46226 23998
rect 3838 23938 3890 23950
rect 3838 23874 3890 23886
rect 4062 23938 4114 23950
rect 4062 23874 4114 23886
rect 6862 23938 6914 23950
rect 6862 23874 6914 23886
rect 7086 23938 7138 23950
rect 12462 23938 12514 23950
rect 13806 23938 13858 23950
rect 19182 23938 19234 23950
rect 19854 23938 19906 23950
rect 7970 23886 7982 23938
rect 8034 23886 8046 23938
rect 11442 23886 11454 23938
rect 11506 23886 11518 23938
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 15698 23886 15710 23938
rect 15762 23886 15774 23938
rect 19394 23886 19406 23938
rect 19458 23935 19470 23938
rect 19618 23935 19630 23938
rect 19458 23889 19630 23935
rect 19458 23886 19470 23889
rect 19618 23886 19630 23889
rect 19682 23886 19694 23938
rect 7086 23874 7138 23886
rect 12462 23874 12514 23886
rect 13806 23874 13858 23886
rect 19182 23874 19234 23886
rect 19854 23874 19906 23886
rect 20078 23938 20130 23950
rect 20078 23874 20130 23886
rect 20302 23938 20354 23950
rect 20302 23874 20354 23886
rect 21198 23938 21250 23950
rect 21198 23874 21250 23886
rect 21534 23938 21586 23950
rect 21534 23874 21586 23886
rect 22206 23938 22258 23950
rect 29710 23938 29762 23950
rect 35310 23938 35362 23950
rect 36206 23938 36258 23950
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 31154 23886 31166 23938
rect 31218 23886 31230 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 35634 23886 35646 23938
rect 35698 23886 35710 23938
rect 22206 23874 22258 23886
rect 29710 23874 29762 23886
rect 35310 23874 35362 23886
rect 36206 23874 36258 23886
rect 37214 23938 37266 23950
rect 37214 23874 37266 23886
rect 37550 23938 37602 23950
rect 37550 23874 37602 23886
rect 37886 23938 37938 23950
rect 37886 23874 37938 23886
rect 39454 23938 39506 23950
rect 39454 23874 39506 23886
rect 39678 23938 39730 23950
rect 39678 23874 39730 23886
rect 40126 23938 40178 23950
rect 40126 23874 40178 23886
rect 42254 23938 42306 23950
rect 42254 23874 42306 23886
rect 42366 23938 42418 23950
rect 43598 23938 43650 23950
rect 42802 23886 42814 23938
rect 42866 23886 42878 23938
rect 43138 23886 43150 23938
rect 43202 23886 43214 23938
rect 42366 23874 42418 23886
rect 43598 23874 43650 23886
rect 3502 23826 3554 23838
rect 3502 23762 3554 23774
rect 6078 23826 6130 23838
rect 6078 23762 6130 23774
rect 6414 23826 6466 23838
rect 6414 23762 6466 23774
rect 7310 23826 7362 23838
rect 12014 23826 12066 23838
rect 10770 23774 10782 23826
rect 10834 23774 10846 23826
rect 7310 23762 7362 23774
rect 12014 23762 12066 23774
rect 19070 23826 19122 23838
rect 19070 23762 19122 23774
rect 22430 23826 22482 23838
rect 22430 23762 22482 23774
rect 22542 23826 22594 23838
rect 36094 23826 36146 23838
rect 25330 23774 25342 23826
rect 25394 23774 25406 23826
rect 22542 23762 22594 23774
rect 36094 23762 36146 23774
rect 36318 23826 36370 23838
rect 36318 23762 36370 23774
rect 36990 23826 37042 23838
rect 36990 23762 37042 23774
rect 38334 23826 38386 23838
rect 38334 23762 38386 23774
rect 44158 23826 44210 23838
rect 44158 23762 44210 23774
rect 45054 23826 45106 23838
rect 45054 23762 45106 23774
rect 3614 23714 3666 23726
rect 4734 23714 4786 23726
rect 4386 23662 4398 23714
rect 4450 23662 4462 23714
rect 3614 23650 3666 23662
rect 4734 23650 4786 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 14030 23714 14082 23726
rect 14030 23650 14082 23662
rect 14254 23714 14306 23726
rect 14254 23650 14306 23662
rect 14926 23714 14978 23726
rect 14926 23650 14978 23662
rect 20414 23714 20466 23726
rect 20414 23650 20466 23662
rect 20526 23714 20578 23726
rect 20526 23650 20578 23662
rect 21422 23714 21474 23726
rect 21422 23650 21474 23662
rect 22094 23714 22146 23726
rect 22094 23650 22146 23662
rect 22990 23714 23042 23726
rect 37438 23714 37490 23726
rect 29138 23662 29150 23714
rect 29202 23662 29214 23714
rect 30594 23662 30606 23714
rect 30658 23662 30670 23714
rect 22990 23650 23042 23662
rect 37438 23650 37490 23662
rect 37998 23714 38050 23726
rect 37998 23650 38050 23662
rect 38110 23714 38162 23726
rect 38110 23650 38162 23662
rect 41806 23714 41858 23726
rect 41806 23650 41858 23662
rect 42590 23714 42642 23726
rect 42590 23650 42642 23662
rect 44046 23714 44098 23726
rect 44046 23650 44098 23662
rect 1344 23546 46592 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 46592 23546
rect 1344 23460 46592 23494
rect 4958 23378 5010 23390
rect 4958 23314 5010 23326
rect 5518 23378 5570 23390
rect 5518 23314 5570 23326
rect 8990 23378 9042 23390
rect 8990 23314 9042 23326
rect 9774 23378 9826 23390
rect 22542 23378 22594 23390
rect 13570 23326 13582 23378
rect 13634 23326 13646 23378
rect 9774 23314 9826 23326
rect 22542 23314 22594 23326
rect 25790 23378 25842 23390
rect 25790 23314 25842 23326
rect 25902 23378 25954 23390
rect 25902 23314 25954 23326
rect 26126 23378 26178 23390
rect 26126 23314 26178 23326
rect 27358 23378 27410 23390
rect 27358 23314 27410 23326
rect 27470 23378 27522 23390
rect 27470 23314 27522 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 28142 23378 28194 23390
rect 28142 23314 28194 23326
rect 28702 23378 28754 23390
rect 28702 23314 28754 23326
rect 35646 23378 35698 23390
rect 35646 23314 35698 23326
rect 36878 23378 36930 23390
rect 36878 23314 36930 23326
rect 40350 23378 40402 23390
rect 40350 23314 40402 23326
rect 41358 23378 41410 23390
rect 41358 23314 41410 23326
rect 5742 23266 5794 23278
rect 2482 23214 2494 23266
rect 2546 23214 2558 23266
rect 5742 23202 5794 23214
rect 7646 23266 7698 23278
rect 7646 23202 7698 23214
rect 8654 23266 8706 23278
rect 8654 23202 8706 23214
rect 8766 23266 8818 23278
rect 8766 23202 8818 23214
rect 10558 23266 10610 23278
rect 22990 23266 23042 23278
rect 14690 23214 14702 23266
rect 14754 23214 14766 23266
rect 17938 23214 17950 23266
rect 18002 23214 18014 23266
rect 20178 23214 20190 23266
rect 20242 23214 20254 23266
rect 10558 23202 10610 23214
rect 22990 23202 23042 23214
rect 23102 23266 23154 23278
rect 23102 23202 23154 23214
rect 24222 23266 24274 23278
rect 24222 23202 24274 23214
rect 26014 23266 26066 23278
rect 26014 23202 26066 23214
rect 26686 23266 26738 23278
rect 26686 23202 26738 23214
rect 33742 23266 33794 23278
rect 33742 23202 33794 23214
rect 39118 23266 39170 23278
rect 39118 23202 39170 23214
rect 40238 23266 40290 23278
rect 40238 23202 40290 23214
rect 41582 23266 41634 23278
rect 41582 23202 41634 23214
rect 42254 23266 42306 23278
rect 42254 23202 42306 23214
rect 42366 23266 42418 23278
rect 42366 23202 42418 23214
rect 42478 23266 42530 23278
rect 45378 23214 45390 23266
rect 45442 23214 45454 23266
rect 42478 23202 42530 23214
rect 5294 23154 5346 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 5294 23090 5346 23102
rect 5854 23154 5906 23166
rect 6638 23154 6690 23166
rect 6402 23102 6414 23154
rect 6466 23102 6478 23154
rect 5854 23090 5906 23102
rect 6638 23090 6690 23102
rect 6862 23154 6914 23166
rect 6862 23090 6914 23102
rect 7198 23154 7250 23166
rect 7198 23090 7250 23102
rect 7534 23154 7586 23166
rect 9438 23154 9490 23166
rect 7746 23102 7758 23154
rect 7810 23102 7822 23154
rect 8194 23102 8206 23154
rect 8258 23102 8270 23154
rect 7534 23090 7586 23102
rect 9438 23090 9490 23102
rect 9886 23154 9938 23166
rect 9886 23090 9938 23102
rect 10110 23154 10162 23166
rect 10110 23090 10162 23102
rect 10334 23154 10386 23166
rect 10334 23090 10386 23102
rect 10670 23154 10722 23166
rect 10670 23090 10722 23102
rect 13022 23154 13074 23166
rect 13022 23090 13074 23102
rect 13246 23154 13298 23166
rect 20638 23154 20690 23166
rect 22654 23154 22706 23166
rect 14018 23102 14030 23154
rect 14082 23102 14094 23154
rect 18274 23102 18286 23154
rect 18338 23102 18350 23154
rect 19618 23102 19630 23154
rect 19682 23102 19694 23154
rect 21746 23102 21758 23154
rect 21810 23102 21822 23154
rect 13246 23090 13298 23102
rect 20638 23090 20690 23102
rect 22654 23090 22706 23102
rect 23662 23154 23714 23166
rect 23662 23090 23714 23102
rect 23998 23154 24050 23166
rect 23998 23090 24050 23102
rect 24334 23154 24386 23166
rect 27246 23154 27298 23166
rect 25554 23102 25566 23154
rect 25618 23102 25630 23154
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 24334 23090 24386 23102
rect 27246 23090 27298 23102
rect 29486 23154 29538 23166
rect 29486 23090 29538 23102
rect 29710 23154 29762 23166
rect 31166 23154 31218 23166
rect 30482 23102 30494 23154
rect 30546 23102 30558 23154
rect 29710 23090 29762 23102
rect 31166 23090 31218 23102
rect 31614 23154 31666 23166
rect 31614 23090 31666 23102
rect 31838 23154 31890 23166
rect 31838 23090 31890 23102
rect 32398 23154 32450 23166
rect 34190 23154 34242 23166
rect 35422 23154 35474 23166
rect 33506 23102 33518 23154
rect 33570 23102 33582 23154
rect 34626 23102 34638 23154
rect 34690 23102 34702 23154
rect 32398 23090 32450 23102
rect 34190 23090 34242 23102
rect 35422 23090 35474 23102
rect 35758 23154 35810 23166
rect 35758 23090 35810 23102
rect 35870 23154 35922 23166
rect 35870 23090 35922 23102
rect 38222 23154 38274 23166
rect 38222 23090 38274 23102
rect 38558 23154 38610 23166
rect 38558 23090 38610 23102
rect 39006 23154 39058 23166
rect 39006 23090 39058 23102
rect 39230 23154 39282 23166
rect 41022 23154 41074 23166
rect 39442 23102 39454 23154
rect 39506 23102 39518 23154
rect 39230 23090 39282 23102
rect 41022 23090 41074 23102
rect 41134 23154 41186 23166
rect 41134 23090 41186 23102
rect 41246 23154 41298 23166
rect 46050 23102 46062 23154
rect 46114 23102 46126 23154
rect 41246 23090 41298 23102
rect 17726 23042 17778 23054
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 16818 22990 16830 23042
rect 16882 22990 16894 23042
rect 17726 22978 17778 22990
rect 26574 23042 26626 23054
rect 26574 22978 26626 22990
rect 29150 23042 29202 23054
rect 31726 23042 31778 23054
rect 30818 22990 30830 23042
rect 30882 22990 30894 23042
rect 29150 22978 29202 22990
rect 31726 22978 31778 22990
rect 35086 23042 35138 23054
rect 36430 23042 36482 23054
rect 36082 22990 36094 23042
rect 36146 22990 36158 23042
rect 43250 22990 43262 23042
rect 43314 22990 43326 23042
rect 35086 22978 35138 22990
rect 7086 22930 7138 22942
rect 22542 22930 22594 22942
rect 8082 22878 8094 22930
rect 8146 22878 8158 22930
rect 7086 22866 7138 22878
rect 22542 22866 22594 22878
rect 23102 22930 23154 22942
rect 23102 22866 23154 22878
rect 23774 22930 23826 22942
rect 30034 22878 30046 22930
rect 30098 22878 30110 22930
rect 36097 22927 36143 22990
rect 36430 22978 36482 22990
rect 38110 22930 38162 22942
rect 36418 22927 36430 22930
rect 36097 22881 36430 22927
rect 36418 22878 36430 22881
rect 36482 22878 36494 22930
rect 23774 22866 23826 22878
rect 38110 22866 38162 22878
rect 38446 22930 38498 22942
rect 38446 22866 38498 22878
rect 39902 22930 39954 22942
rect 42914 22878 42926 22930
rect 42978 22878 42990 22930
rect 39902 22866 39954 22878
rect 1344 22762 46592 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 46592 22762
rect 1344 22676 46592 22710
rect 27246 22594 27298 22606
rect 19618 22542 19630 22594
rect 19682 22542 19694 22594
rect 21298 22542 21310 22594
rect 21362 22591 21374 22594
rect 21522 22591 21534 22594
rect 21362 22545 21534 22591
rect 21362 22542 21374 22545
rect 21522 22542 21534 22545
rect 21586 22542 21598 22594
rect 27246 22530 27298 22542
rect 27582 22594 27634 22606
rect 27582 22530 27634 22542
rect 41022 22594 41074 22606
rect 41022 22530 41074 22542
rect 42366 22594 42418 22606
rect 42366 22530 42418 22542
rect 43822 22594 43874 22606
rect 43822 22530 43874 22542
rect 17950 22482 18002 22494
rect 43150 22482 43202 22494
rect 4722 22430 4734 22482
rect 4786 22430 4798 22482
rect 6738 22430 6750 22482
rect 6802 22430 6814 22482
rect 12898 22430 12910 22482
rect 12962 22430 12974 22482
rect 18498 22430 18510 22482
rect 18562 22430 18574 22482
rect 19282 22430 19294 22482
rect 19346 22430 19358 22482
rect 23090 22430 23102 22482
rect 23154 22430 23166 22482
rect 25218 22430 25230 22482
rect 25282 22430 25294 22482
rect 26786 22430 26798 22482
rect 26850 22430 26862 22482
rect 39218 22430 39230 22482
rect 39282 22430 39294 22482
rect 17950 22418 18002 22430
rect 43150 22418 43202 22430
rect 43710 22482 43762 22494
rect 43710 22418 43762 22430
rect 45054 22482 45106 22494
rect 45054 22418 45106 22430
rect 45614 22482 45666 22494
rect 45614 22418 45666 22430
rect 21870 22370 21922 22382
rect 25790 22370 25842 22382
rect 4050 22318 4062 22370
rect 4114 22318 4126 22370
rect 4386 22318 4398 22370
rect 4450 22318 4462 22370
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 9986 22318 9998 22370
rect 10050 22318 10062 22370
rect 13682 22318 13694 22370
rect 13746 22318 13758 22370
rect 15698 22318 15710 22370
rect 15762 22318 15774 22370
rect 18610 22318 18622 22370
rect 18674 22318 18686 22370
rect 19730 22318 19742 22370
rect 19794 22318 19806 22370
rect 22306 22318 22318 22370
rect 22370 22318 22382 22370
rect 21870 22306 21922 22318
rect 25790 22306 25842 22318
rect 28030 22370 28082 22382
rect 30046 22370 30098 22382
rect 37662 22370 37714 22382
rect 42702 22370 42754 22382
rect 29362 22318 29374 22370
rect 29426 22318 29438 22370
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 39330 22318 39342 22370
rect 39394 22318 39406 22370
rect 40002 22318 40014 22370
rect 40066 22318 40078 22370
rect 28030 22306 28082 22318
rect 30046 22306 30098 22318
rect 37662 22306 37714 22318
rect 42702 22306 42754 22318
rect 43038 22370 43090 22382
rect 43038 22306 43090 22318
rect 44046 22370 44098 22382
rect 44046 22306 44098 22318
rect 5742 22258 5794 22270
rect 3378 22206 3390 22258
rect 3442 22206 3454 22258
rect 4946 22206 4958 22258
rect 5010 22206 5022 22258
rect 5742 22194 5794 22206
rect 5854 22258 5906 22270
rect 14814 22258 14866 22270
rect 8866 22206 8878 22258
rect 8930 22206 8942 22258
rect 10770 22206 10782 22258
rect 10834 22206 10846 22258
rect 5854 22194 5906 22206
rect 14814 22194 14866 22206
rect 16270 22258 16322 22270
rect 16270 22194 16322 22206
rect 20414 22258 20466 22270
rect 20414 22194 20466 22206
rect 25678 22258 25730 22270
rect 25678 22194 25730 22206
rect 27358 22258 27410 22270
rect 27358 22194 27410 22206
rect 29150 22258 29202 22270
rect 29150 22194 29202 22206
rect 29598 22258 29650 22270
rect 37326 22258 37378 22270
rect 40910 22258 40962 22270
rect 33842 22206 33854 22258
rect 33906 22206 33918 22258
rect 37986 22206 37998 22258
rect 38050 22206 38062 22258
rect 39554 22206 39566 22258
rect 39618 22206 39630 22258
rect 29598 22194 29650 22206
rect 37326 22194 37378 22206
rect 40910 22194 40962 22206
rect 41806 22258 41858 22270
rect 41806 22194 41858 22206
rect 43262 22258 43314 22270
rect 43262 22194 43314 22206
rect 44158 22258 44210 22270
rect 44158 22194 44210 22206
rect 45838 22258 45890 22270
rect 45838 22194 45890 22206
rect 46174 22258 46226 22270
rect 46174 22194 46226 22206
rect 5518 22146 5570 22158
rect 5518 22082 5570 22094
rect 6302 22146 6354 22158
rect 20526 22146 20578 22158
rect 13794 22094 13806 22146
rect 13858 22094 13870 22146
rect 6302 22082 6354 22094
rect 20526 22082 20578 22094
rect 21534 22146 21586 22158
rect 21534 22082 21586 22094
rect 21982 22146 22034 22158
rect 21982 22082 22034 22094
rect 25454 22146 25506 22158
rect 25454 22082 25506 22094
rect 26350 22146 26402 22158
rect 26350 22082 26402 22094
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 29038 22146 29090 22158
rect 36430 22146 36482 22158
rect 35970 22094 35982 22146
rect 36034 22143 36046 22146
rect 36194 22143 36206 22146
rect 36034 22097 36206 22143
rect 36034 22094 36046 22097
rect 36194 22094 36206 22097
rect 36258 22094 36270 22146
rect 29038 22082 29090 22094
rect 36430 22082 36482 22094
rect 36990 22146 37042 22158
rect 36990 22082 37042 22094
rect 38894 22146 38946 22158
rect 38894 22082 38946 22094
rect 42142 22146 42194 22158
rect 42142 22082 42194 22094
rect 42254 22146 42306 22158
rect 42254 22082 42306 22094
rect 1344 21978 46592 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 46592 21978
rect 1344 21892 46592 21926
rect 5966 21810 6018 21822
rect 5966 21746 6018 21758
rect 6974 21810 7026 21822
rect 6974 21746 7026 21758
rect 7870 21810 7922 21822
rect 7870 21746 7922 21758
rect 8430 21810 8482 21822
rect 8430 21746 8482 21758
rect 9662 21810 9714 21822
rect 9662 21746 9714 21758
rect 14142 21810 14194 21822
rect 14142 21746 14194 21758
rect 15934 21810 15986 21822
rect 15934 21746 15986 21758
rect 17726 21810 17778 21822
rect 17726 21746 17778 21758
rect 23214 21810 23266 21822
rect 23214 21746 23266 21758
rect 24334 21810 24386 21822
rect 24334 21746 24386 21758
rect 26126 21810 26178 21822
rect 26126 21746 26178 21758
rect 29710 21810 29762 21822
rect 29710 21746 29762 21758
rect 32062 21810 32114 21822
rect 32062 21746 32114 21758
rect 33742 21810 33794 21822
rect 33742 21746 33794 21758
rect 37774 21810 37826 21822
rect 37774 21746 37826 21758
rect 38894 21810 38946 21822
rect 38894 21746 38946 21758
rect 39678 21810 39730 21822
rect 39678 21746 39730 21758
rect 39790 21810 39842 21822
rect 39790 21746 39842 21758
rect 39902 21810 39954 21822
rect 39902 21746 39954 21758
rect 40238 21810 40290 21822
rect 40238 21746 40290 21758
rect 5854 21698 5906 21710
rect 4946 21646 4958 21698
rect 5010 21646 5022 21698
rect 5854 21634 5906 21646
rect 7086 21698 7138 21710
rect 7086 21634 7138 21646
rect 7758 21698 7810 21710
rect 7758 21634 7810 21646
rect 8318 21698 8370 21710
rect 8318 21634 8370 21646
rect 10110 21698 10162 21710
rect 10110 21634 10162 21646
rect 13358 21698 13410 21710
rect 13358 21634 13410 21646
rect 13918 21698 13970 21710
rect 22990 21698 23042 21710
rect 17378 21646 17390 21698
rect 17442 21646 17454 21698
rect 18834 21646 18846 21698
rect 18898 21646 18910 21698
rect 13918 21634 13970 21646
rect 22990 21634 23042 21646
rect 24110 21698 24162 21710
rect 24110 21634 24162 21646
rect 25230 21698 25282 21710
rect 28690 21646 28702 21698
rect 28754 21646 28766 21698
rect 32386 21646 32398 21698
rect 32450 21646 32462 21698
rect 35298 21646 35310 21698
rect 35362 21646 35374 21698
rect 38098 21646 38110 21698
rect 38162 21646 38174 21698
rect 45378 21646 45390 21698
rect 45442 21646 45454 21698
rect 25230 21634 25282 21646
rect 5294 21586 5346 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 5294 21522 5346 21534
rect 6190 21586 6242 21598
rect 6190 21522 6242 21534
rect 6750 21586 6802 21598
rect 6750 21522 6802 21534
rect 8094 21586 8146 21598
rect 8094 21522 8146 21534
rect 8654 21586 8706 21598
rect 8654 21522 8706 21534
rect 9438 21586 9490 21598
rect 9438 21522 9490 21534
rect 9774 21586 9826 21598
rect 14814 21586 14866 21598
rect 14466 21534 14478 21586
rect 14530 21534 14542 21586
rect 9774 21522 9826 21534
rect 14814 21522 14866 21534
rect 15038 21586 15090 21598
rect 22542 21586 22594 21598
rect 30158 21586 30210 21598
rect 31502 21586 31554 21598
rect 38558 21586 38610 21598
rect 16706 21534 16718 21586
rect 16770 21534 16782 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 22082 21534 22094 21586
rect 22146 21534 22158 21586
rect 22866 21534 22878 21586
rect 22930 21534 22942 21586
rect 23986 21534 23998 21586
rect 24050 21534 24062 21586
rect 25554 21534 25566 21586
rect 25618 21534 25630 21586
rect 29474 21534 29486 21586
rect 29538 21534 29550 21586
rect 31154 21534 31166 21586
rect 31218 21534 31230 21586
rect 34514 21534 34526 21586
rect 34578 21534 34590 21586
rect 15038 21522 15090 21534
rect 22542 21522 22594 21534
rect 30158 21522 30210 21534
rect 31502 21522 31554 21534
rect 38558 21522 38610 21534
rect 39230 21586 39282 21598
rect 39230 21522 39282 21534
rect 42366 21586 42418 21598
rect 46050 21534 46062 21586
rect 46114 21534 46126 21586
rect 42366 21522 42418 21534
rect 14030 21474 14082 21486
rect 23102 21474 23154 21486
rect 2482 21422 2494 21474
rect 2546 21422 2558 21474
rect 4610 21422 4622 21474
rect 4674 21422 4686 21474
rect 13234 21422 13246 21474
rect 13298 21422 13310 21474
rect 16370 21422 16382 21474
rect 16434 21422 16446 21474
rect 19170 21422 19182 21474
rect 19234 21422 19246 21474
rect 21298 21422 21310 21474
rect 21362 21422 21374 21474
rect 14030 21410 14082 21422
rect 23102 21410 23154 21422
rect 24222 21474 24274 21486
rect 24222 21410 24274 21422
rect 25342 21474 25394 21486
rect 25342 21410 25394 21422
rect 26238 21474 26290 21486
rect 30606 21474 30658 21486
rect 26562 21422 26574 21474
rect 26626 21422 26638 21474
rect 26238 21410 26290 21422
rect 30606 21410 30658 21422
rect 31726 21474 31778 21486
rect 31726 21410 31778 21422
rect 33182 21474 33234 21486
rect 39006 21474 39058 21486
rect 37426 21422 37438 21474
rect 37490 21422 37502 21474
rect 33182 21410 33234 21422
rect 39006 21410 39058 21422
rect 40350 21474 40402 21486
rect 40350 21410 40402 21422
rect 41806 21474 41858 21486
rect 41806 21410 41858 21422
rect 42142 21474 42194 21486
rect 43250 21422 43262 21474
rect 43314 21422 43326 21474
rect 42142 21410 42194 21422
rect 13582 21362 13634 21374
rect 18734 21362 18786 21374
rect 15362 21310 15374 21362
rect 15426 21310 15438 21362
rect 13582 21298 13634 21310
rect 18734 21298 18786 21310
rect 23662 21362 23714 21374
rect 23662 21298 23714 21310
rect 30382 21362 30434 21374
rect 30382 21298 30434 21310
rect 33070 21362 33122 21374
rect 41582 21362 41634 21374
rect 41234 21310 41246 21362
rect 41298 21310 41310 21362
rect 42690 21310 42702 21362
rect 42754 21310 42766 21362
rect 33070 21298 33122 21310
rect 41582 21298 41634 21310
rect 1344 21194 46592 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 46592 21194
rect 1344 21108 46592 21142
rect 21310 21026 21362 21038
rect 20514 20974 20526 21026
rect 20578 21023 20590 21026
rect 20850 21023 20862 21026
rect 20578 20977 20862 21023
rect 20578 20974 20590 20977
rect 20850 20974 20862 20977
rect 20914 20974 20926 21026
rect 21310 20962 21362 20974
rect 35310 21026 35362 21038
rect 35310 20962 35362 20974
rect 35646 21026 35698 21038
rect 44942 21026 44994 21038
rect 35858 20974 35870 21026
rect 35922 21023 35934 21026
rect 36418 21023 36430 21026
rect 35922 20977 36430 21023
rect 35922 20974 35934 20977
rect 36418 20974 36430 20977
rect 36482 20974 36494 21026
rect 35646 20962 35698 20974
rect 44942 20962 44994 20974
rect 45166 21026 45218 21038
rect 45166 20962 45218 20974
rect 45278 21026 45330 21038
rect 45278 20962 45330 20974
rect 12910 20914 12962 20926
rect 21534 20914 21586 20926
rect 8754 20862 8766 20914
rect 8818 20862 8830 20914
rect 10882 20862 10894 20914
rect 10946 20862 10958 20914
rect 18162 20862 18174 20914
rect 18226 20862 18238 20914
rect 12910 20850 12962 20862
rect 21534 20850 21586 20862
rect 21870 20914 21922 20926
rect 21870 20850 21922 20862
rect 29598 20914 29650 20926
rect 35086 20914 35138 20926
rect 34178 20862 34190 20914
rect 34242 20862 34254 20914
rect 29598 20850 29650 20862
rect 35086 20850 35138 20862
rect 36206 20914 36258 20926
rect 36206 20850 36258 20862
rect 39566 20914 39618 20926
rect 39566 20850 39618 20862
rect 40350 20914 40402 20926
rect 45950 20914 46002 20926
rect 41010 20862 41022 20914
rect 41074 20862 41086 20914
rect 41346 20862 41358 20914
rect 41410 20862 41422 20914
rect 40350 20850 40402 20862
rect 45950 20850 46002 20862
rect 2382 20802 2434 20814
rect 2382 20738 2434 20750
rect 2718 20802 2770 20814
rect 2718 20738 2770 20750
rect 3950 20802 4002 20814
rect 3950 20738 4002 20750
rect 4622 20802 4674 20814
rect 12686 20802 12738 20814
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 4622 20738 4674 20750
rect 12686 20738 12738 20750
rect 14030 20802 14082 20814
rect 14030 20738 14082 20750
rect 14254 20802 14306 20814
rect 19070 20802 19122 20814
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 14254 20738 14306 20750
rect 19070 20738 19122 20750
rect 19182 20802 19234 20814
rect 19182 20738 19234 20750
rect 19854 20802 19906 20814
rect 19854 20738 19906 20750
rect 21758 20802 21810 20814
rect 21758 20738 21810 20750
rect 21982 20802 22034 20814
rect 23998 20802 24050 20814
rect 29038 20802 29090 20814
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 24994 20750 25006 20802
rect 25058 20750 25070 20802
rect 26338 20750 26350 20802
rect 26402 20750 26414 20802
rect 27010 20750 27022 20802
rect 27074 20750 27086 20802
rect 21982 20738 22034 20750
rect 23998 20738 24050 20750
rect 29038 20738 29090 20750
rect 29710 20802 29762 20814
rect 37326 20802 37378 20814
rect 39678 20802 39730 20814
rect 31378 20750 31390 20802
rect 31442 20750 31454 20802
rect 32050 20750 32062 20802
rect 32114 20750 32126 20802
rect 37762 20750 37774 20802
rect 37826 20750 37838 20802
rect 44258 20750 44270 20802
rect 44322 20750 44334 20802
rect 29710 20738 29762 20750
rect 37326 20738 37378 20750
rect 39678 20738 39730 20750
rect 2830 20690 2882 20702
rect 2830 20626 2882 20638
rect 3054 20690 3106 20702
rect 3054 20626 3106 20638
rect 3278 20690 3330 20702
rect 3278 20626 3330 20638
rect 3502 20690 3554 20702
rect 3502 20626 3554 20638
rect 4174 20690 4226 20702
rect 4174 20626 4226 20638
rect 4510 20690 4562 20702
rect 11230 20690 11282 20702
rect 18958 20690 19010 20702
rect 27246 20690 27298 20702
rect 6626 20638 6638 20690
rect 6690 20638 6702 20690
rect 9426 20638 9438 20690
rect 9490 20638 9502 20690
rect 16034 20638 16046 20690
rect 16098 20638 16110 20690
rect 25778 20638 25790 20690
rect 25842 20638 25854 20690
rect 4510 20626 4562 20638
rect 11230 20626 11282 20638
rect 18958 20626 19010 20638
rect 27246 20626 27298 20638
rect 27358 20690 27410 20702
rect 27358 20626 27410 20638
rect 30718 20690 30770 20702
rect 38782 20690 38834 20702
rect 36978 20638 36990 20690
rect 37042 20638 37054 20690
rect 37986 20638 37998 20690
rect 38050 20638 38062 20690
rect 30718 20626 30770 20638
rect 38782 20626 38834 20638
rect 39902 20690 39954 20702
rect 39902 20626 39954 20638
rect 40686 20690 40738 20702
rect 40686 20626 40738 20638
rect 40910 20690 40962 20702
rect 44830 20690 44882 20702
rect 43474 20638 43486 20690
rect 43538 20638 43550 20690
rect 40910 20626 40962 20638
rect 44830 20626 44882 20638
rect 2046 20578 2098 20590
rect 2046 20514 2098 20526
rect 2270 20578 2322 20590
rect 2270 20514 2322 20526
rect 3614 20578 3666 20590
rect 3614 20514 3666 20526
rect 4286 20578 4338 20590
rect 4286 20514 4338 20526
rect 9102 20578 9154 20590
rect 9102 20514 9154 20526
rect 11006 20578 11058 20590
rect 11006 20514 11058 20526
rect 11790 20578 11842 20590
rect 14142 20578 14194 20590
rect 12338 20526 12350 20578
rect 12402 20526 12414 20578
rect 11790 20514 11842 20526
rect 14142 20514 14194 20526
rect 14478 20578 14530 20590
rect 20302 20578 20354 20590
rect 18498 20526 18510 20578
rect 18562 20526 18574 20578
rect 14478 20514 14530 20526
rect 20302 20514 20354 20526
rect 20750 20578 20802 20590
rect 28142 20578 28194 20590
rect 29486 20578 29538 20590
rect 22754 20526 22766 20578
rect 22818 20526 22830 20578
rect 27794 20526 27806 20578
rect 27858 20526 27870 20578
rect 28466 20526 28478 20578
rect 28530 20526 28542 20578
rect 20750 20514 20802 20526
rect 28142 20514 28194 20526
rect 29486 20514 29538 20526
rect 30046 20578 30098 20590
rect 30830 20578 30882 20590
rect 30370 20526 30382 20578
rect 30434 20526 30446 20578
rect 30046 20514 30098 20526
rect 30830 20514 30882 20526
rect 34750 20578 34802 20590
rect 34750 20514 34802 20526
rect 38558 20578 38610 20590
rect 38558 20514 38610 20526
rect 38894 20578 38946 20590
rect 38894 20514 38946 20526
rect 39342 20578 39394 20590
rect 39342 20514 39394 20526
rect 39454 20578 39506 20590
rect 39454 20514 39506 20526
rect 40238 20578 40290 20590
rect 40238 20514 40290 20526
rect 1344 20410 46592 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 46592 20410
rect 1344 20324 46592 20358
rect 17614 20242 17666 20254
rect 17614 20178 17666 20190
rect 23662 20242 23714 20254
rect 23662 20178 23714 20190
rect 27806 20242 27858 20254
rect 27806 20178 27858 20190
rect 30046 20242 30098 20254
rect 30046 20178 30098 20190
rect 30718 20242 30770 20254
rect 30718 20178 30770 20190
rect 31726 20242 31778 20254
rect 31726 20178 31778 20190
rect 33406 20242 33458 20254
rect 33406 20178 33458 20190
rect 38894 20242 38946 20254
rect 38894 20178 38946 20190
rect 2046 20130 2098 20142
rect 2046 20066 2098 20078
rect 2270 20130 2322 20142
rect 2270 20066 2322 20078
rect 8542 20130 8594 20142
rect 8542 20066 8594 20078
rect 8878 20130 8930 20142
rect 17838 20130 17890 20142
rect 15250 20078 15262 20130
rect 15314 20078 15326 20130
rect 8878 20066 8930 20078
rect 17838 20066 17890 20078
rect 18174 20130 18226 20142
rect 18174 20066 18226 20078
rect 19294 20130 19346 20142
rect 19294 20066 19346 20078
rect 20078 20130 20130 20142
rect 24334 20130 24386 20142
rect 21186 20078 21198 20130
rect 21250 20078 21262 20130
rect 20078 20066 20130 20078
rect 24334 20066 24386 20078
rect 27358 20130 27410 20142
rect 27358 20066 27410 20078
rect 34190 20130 34242 20142
rect 34190 20066 34242 20078
rect 36094 20130 36146 20142
rect 36094 20066 36146 20078
rect 38446 20130 38498 20142
rect 38446 20066 38498 20078
rect 39006 20130 39058 20142
rect 39006 20066 39058 20078
rect 39118 20130 39170 20142
rect 39118 20066 39170 20078
rect 2606 20018 2658 20030
rect 18286 20018 18338 20030
rect 23774 20018 23826 20030
rect 8194 19966 8206 20018
rect 8258 19966 8270 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 20514 19966 20526 20018
rect 20578 19966 20590 20018
rect 2606 19954 2658 19966
rect 18286 19954 18338 19966
rect 23774 19954 23826 19966
rect 26462 20018 26514 20030
rect 26462 19954 26514 19966
rect 26686 20018 26738 20030
rect 26686 19954 26738 19966
rect 26798 20018 26850 20030
rect 26798 19954 26850 19966
rect 27022 20018 27074 20030
rect 27022 19954 27074 19966
rect 27582 20018 27634 20030
rect 33294 20018 33346 20030
rect 33058 19966 33070 20018
rect 33122 19966 33134 20018
rect 27582 19954 27634 19966
rect 33294 19954 33346 19966
rect 33518 20018 33570 20030
rect 33518 19954 33570 19966
rect 33630 20018 33682 20030
rect 33630 19954 33682 19966
rect 34302 20018 34354 20030
rect 34302 19954 34354 19966
rect 34526 20018 34578 20030
rect 38782 20018 38834 20030
rect 40014 20018 40066 20030
rect 34738 19966 34750 20018
rect 34802 19966 34814 20018
rect 39554 19966 39566 20018
rect 39618 19966 39630 20018
rect 40226 19966 40238 20018
rect 40290 19966 40302 20018
rect 40898 19966 40910 20018
rect 40962 19966 40974 20018
rect 34526 19954 34578 19966
rect 38782 19954 38834 19966
rect 40014 19954 40066 19966
rect 2494 19906 2546 19918
rect 9774 19906 9826 19918
rect 3378 19854 3390 19906
rect 3442 19854 3454 19906
rect 2494 19842 2546 19854
rect 9774 19842 9826 19854
rect 17950 19906 18002 19918
rect 24670 19906 24722 19918
rect 18834 19854 18846 19906
rect 18898 19854 18910 19906
rect 23314 19854 23326 19906
rect 23378 19854 23390 19906
rect 17950 19842 18002 19854
rect 24670 19842 24722 19854
rect 26014 19906 26066 19918
rect 26014 19842 26066 19854
rect 27694 19906 27746 19918
rect 27694 19842 27746 19854
rect 28254 19906 28306 19918
rect 28254 19842 28306 19854
rect 28702 19906 28754 19918
rect 28702 19842 28754 19854
rect 29150 19906 29202 19918
rect 29150 19842 29202 19854
rect 29598 19906 29650 19918
rect 29598 19842 29650 19854
rect 31278 19906 31330 19918
rect 31278 19842 31330 19854
rect 34414 19906 34466 19918
rect 34414 19842 34466 19854
rect 35086 19906 35138 19918
rect 35086 19842 35138 19854
rect 35646 19906 35698 19918
rect 35646 19842 35698 19854
rect 36654 19906 36706 19918
rect 36654 19842 36706 19854
rect 37102 19906 37154 19918
rect 37102 19842 37154 19854
rect 37550 19906 37602 19918
rect 37550 19842 37602 19854
rect 37886 19906 37938 19918
rect 44706 19854 44718 19906
rect 44770 19854 44782 19906
rect 37886 19842 37938 19854
rect 31166 19794 31218 19806
rect 31166 19730 31218 19742
rect 35198 19794 35250 19806
rect 35198 19730 35250 19742
rect 35534 19794 35586 19806
rect 35534 19730 35586 19742
rect 38222 19794 38274 19806
rect 38222 19730 38274 19742
rect 39902 19794 39954 19806
rect 39902 19730 39954 19742
rect 1344 19626 46592 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 46592 19626
rect 1344 19540 46592 19574
rect 8542 19458 8594 19470
rect 8082 19406 8094 19458
rect 8146 19406 8158 19458
rect 8542 19394 8594 19406
rect 16158 19458 16210 19470
rect 16158 19394 16210 19406
rect 16270 19458 16322 19470
rect 16270 19394 16322 19406
rect 16494 19458 16546 19470
rect 45278 19458 45330 19470
rect 29586 19455 29598 19458
rect 16494 19394 16546 19406
rect 29041 19409 29598 19455
rect 6638 19346 6690 19358
rect 21534 19346 21586 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 12898 19294 12910 19346
rect 12962 19294 12974 19346
rect 13794 19294 13806 19346
rect 13858 19294 13870 19346
rect 18162 19294 18174 19346
rect 18226 19294 18238 19346
rect 6638 19282 6690 19294
rect 21534 19282 21586 19294
rect 22430 19346 22482 19358
rect 22430 19282 22482 19294
rect 23102 19346 23154 19358
rect 29041 19346 29087 19409
rect 29586 19406 29598 19409
rect 29650 19406 29662 19458
rect 45278 19394 45330 19406
rect 45726 19458 45778 19470
rect 45726 19394 45778 19406
rect 39678 19346 39730 19358
rect 25330 19294 25342 19346
rect 25394 19294 25406 19346
rect 29026 19294 29038 19346
rect 29090 19294 29102 19346
rect 30706 19294 30718 19346
rect 30770 19294 30782 19346
rect 32834 19294 32846 19346
rect 32898 19294 32910 19346
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 35634 19294 35646 19346
rect 35698 19294 35710 19346
rect 38658 19294 38670 19346
rect 38722 19294 38734 19346
rect 23102 19282 23154 19294
rect 39678 19282 39730 19294
rect 41022 19346 41074 19358
rect 41346 19294 41358 19346
rect 41410 19294 41422 19346
rect 41022 19282 41074 19294
rect 5518 19234 5570 19246
rect 1810 19182 1822 19234
rect 1874 19182 1886 19234
rect 5518 19170 5570 19182
rect 6190 19234 6242 19246
rect 6190 19170 6242 19182
rect 6414 19234 6466 19246
rect 6414 19170 6466 19182
rect 6750 19234 6802 19246
rect 6750 19170 6802 19182
rect 7534 19234 7586 19246
rect 7534 19170 7586 19182
rect 7758 19234 7810 19246
rect 7758 19170 7810 19182
rect 8654 19234 8706 19246
rect 13582 19234 13634 19246
rect 15038 19234 15090 19246
rect 10098 19182 10110 19234
rect 10162 19182 10174 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 8654 19170 8706 19182
rect 13582 19170 13634 19182
rect 15038 19170 15090 19182
rect 15262 19234 15314 19246
rect 17054 19234 17106 19246
rect 16706 19182 16718 19234
rect 16770 19182 16782 19234
rect 15262 19170 15314 19182
rect 17054 19170 17106 19182
rect 17390 19234 17442 19246
rect 39006 19234 39058 19246
rect 44942 19234 44994 19246
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 19506 19182 19518 19234
rect 19570 19182 19582 19234
rect 21970 19182 21982 19234
rect 22034 19182 22046 19234
rect 24658 19182 24670 19234
rect 24722 19182 24734 19234
rect 29922 19182 29934 19234
rect 29986 19182 29998 19234
rect 36418 19182 36430 19234
rect 36482 19182 36494 19234
rect 40450 19182 40462 19234
rect 40514 19182 40526 19234
rect 40786 19182 40798 19234
rect 40850 19182 40862 19234
rect 44258 19182 44270 19234
rect 44322 19182 44334 19234
rect 17390 19170 17442 19182
rect 39006 19170 39058 19182
rect 44942 19170 44994 19182
rect 45166 19234 45218 19246
rect 45166 19170 45218 19182
rect 45838 19234 45890 19246
rect 45838 19170 45890 19182
rect 5742 19122 5794 19134
rect 5742 19058 5794 19070
rect 5854 19122 5906 19134
rect 17166 19122 17218 19134
rect 10770 19070 10782 19122
rect 10834 19070 10846 19122
rect 5854 19058 5906 19070
rect 17166 19058 17218 19070
rect 19966 19122 20018 19134
rect 37214 19122 37266 19134
rect 20402 19070 20414 19122
rect 20466 19070 20478 19122
rect 19966 19058 20018 19070
rect 37214 19058 37266 19070
rect 39230 19122 39282 19134
rect 44830 19122 44882 19134
rect 43474 19070 43486 19122
rect 43538 19070 43550 19122
rect 39230 19058 39282 19070
rect 44830 19058 44882 19070
rect 45950 19122 46002 19134
rect 45950 19058 46002 19070
rect 7198 19010 7250 19022
rect 7198 18946 7250 18958
rect 8542 19010 8594 19022
rect 8542 18946 8594 18958
rect 9102 19010 9154 19022
rect 20750 19010 20802 19022
rect 15586 18958 15598 19010
rect 15650 18958 15662 19010
rect 9102 18946 9154 18958
rect 20750 18946 20802 18958
rect 21422 19010 21474 19022
rect 21422 18946 21474 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 36878 19010 36930 19022
rect 36878 18946 36930 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 37886 19010 37938 19022
rect 38670 19010 38722 19022
rect 38210 18958 38222 19010
rect 38274 18958 38286 19010
rect 37886 18946 37938 18958
rect 38670 18946 38722 18958
rect 38782 19010 38834 19022
rect 38782 18946 38834 18958
rect 1344 18842 46592 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 46592 18842
rect 1344 18756 46592 18790
rect 8654 18674 8706 18686
rect 8654 18610 8706 18622
rect 11006 18674 11058 18686
rect 11006 18610 11058 18622
rect 12014 18674 12066 18686
rect 12014 18610 12066 18622
rect 17726 18674 17778 18686
rect 17726 18610 17778 18622
rect 31726 18674 31778 18686
rect 31726 18610 31778 18622
rect 31838 18674 31890 18686
rect 31838 18610 31890 18622
rect 39790 18674 39842 18686
rect 39790 18610 39842 18622
rect 19406 18562 19458 18574
rect 17378 18510 17390 18562
rect 17442 18510 17454 18562
rect 18274 18510 18286 18562
rect 18338 18510 18350 18562
rect 19406 18498 19458 18510
rect 20190 18562 20242 18574
rect 20190 18498 20242 18510
rect 25230 18562 25282 18574
rect 25230 18498 25282 18510
rect 30046 18562 30098 18574
rect 30046 18498 30098 18510
rect 32062 18562 32114 18574
rect 39566 18562 39618 18574
rect 38882 18510 38894 18562
rect 38946 18510 38958 18562
rect 32062 18498 32114 18510
rect 39566 18498 39618 18510
rect 44158 18562 44210 18574
rect 44158 18498 44210 18510
rect 44942 18562 44994 18574
rect 44942 18498 44994 18510
rect 45166 18562 45218 18574
rect 45166 18498 45218 18510
rect 45278 18562 45330 18574
rect 45278 18498 45330 18510
rect 12238 18450 12290 18462
rect 16606 18450 16658 18462
rect 20414 18450 20466 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 2482 18398 2494 18450
rect 2546 18398 2558 18450
rect 5282 18398 5294 18450
rect 5346 18398 5358 18450
rect 6066 18398 6078 18450
rect 6130 18398 6142 18450
rect 15362 18398 15374 18450
rect 15426 18398 15438 18450
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 19058 18398 19070 18450
rect 19122 18398 19134 18450
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 12238 18386 12290 18398
rect 16606 18386 16658 18398
rect 20414 18386 20466 18398
rect 20526 18450 20578 18462
rect 20526 18386 20578 18398
rect 21310 18450 21362 18462
rect 21310 18386 21362 18398
rect 21534 18450 21586 18462
rect 21534 18386 21586 18398
rect 21758 18450 21810 18462
rect 21758 18386 21810 18398
rect 22094 18450 22146 18462
rect 22094 18386 22146 18398
rect 22430 18450 22482 18462
rect 22430 18386 22482 18398
rect 23326 18450 23378 18462
rect 23326 18386 23378 18398
rect 24334 18450 24386 18462
rect 29822 18450 29874 18462
rect 25442 18398 25454 18450
rect 25506 18398 25518 18450
rect 26338 18398 26350 18450
rect 26402 18398 26414 18450
rect 29586 18398 29598 18450
rect 29650 18398 29662 18450
rect 24334 18386 24386 18398
rect 29822 18386 29874 18398
rect 30158 18450 30210 18462
rect 30158 18386 30210 18398
rect 31502 18450 31554 18462
rect 31502 18386 31554 18398
rect 31614 18450 31666 18462
rect 31614 18386 31666 18398
rect 32510 18450 32562 18462
rect 32510 18386 32562 18398
rect 33518 18450 33570 18462
rect 44382 18450 44434 18462
rect 33842 18398 33854 18450
rect 33906 18398 33918 18450
rect 40898 18398 40910 18450
rect 40962 18398 40974 18450
rect 41682 18398 41694 18450
rect 41746 18398 41758 18450
rect 33518 18386 33570 18398
rect 44382 18386 44434 18398
rect 44830 18450 44882 18462
rect 44830 18386 44882 18398
rect 8542 18338 8594 18350
rect 4610 18286 4622 18338
rect 4674 18286 4686 18338
rect 8194 18286 8206 18338
rect 8258 18286 8270 18338
rect 8542 18274 8594 18286
rect 11118 18338 11170 18350
rect 15934 18338 15986 18350
rect 11890 18286 11902 18338
rect 11954 18286 11966 18338
rect 12562 18286 12574 18338
rect 12626 18286 12638 18338
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 11118 18274 11170 18286
rect 15934 18274 15986 18286
rect 16830 18338 16882 18350
rect 20302 18338 20354 18350
rect 18722 18286 18734 18338
rect 18786 18286 18798 18338
rect 16830 18274 16882 18286
rect 20302 18274 20354 18286
rect 21646 18338 21698 18350
rect 21646 18274 21698 18286
rect 22990 18338 23042 18350
rect 22990 18274 23042 18286
rect 23886 18338 23938 18350
rect 29934 18338 29986 18350
rect 27122 18286 27134 18338
rect 27186 18286 27198 18338
rect 29250 18286 29262 18338
rect 29314 18286 29326 18338
rect 23886 18274 23938 18286
rect 29934 18274 29986 18286
rect 30718 18338 30770 18350
rect 40238 18338 40290 18350
rect 44606 18338 44658 18350
rect 39890 18286 39902 18338
rect 39954 18286 39966 18338
rect 43810 18286 43822 18338
rect 43874 18286 43886 18338
rect 30718 18274 30770 18286
rect 40238 18274 40290 18286
rect 44606 18274 44658 18286
rect 45726 18338 45778 18350
rect 45726 18274 45778 18286
rect 46174 18338 46226 18350
rect 46174 18274 46226 18286
rect 11230 18226 11282 18238
rect 40350 18226 40402 18238
rect 16258 18174 16270 18226
rect 16322 18174 16334 18226
rect 11230 18162 11282 18174
rect 40350 18162 40402 18174
rect 45614 18226 45666 18238
rect 45614 18162 45666 18174
rect 1344 18058 46592 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 46592 18058
rect 1344 17972 46592 18006
rect 27806 17890 27858 17902
rect 20402 17838 20414 17890
rect 20466 17887 20478 17890
rect 20466 17841 20799 17887
rect 20466 17838 20478 17841
rect 6526 17778 6578 17790
rect 20753 17778 20799 17841
rect 27806 17826 27858 17838
rect 29150 17890 29202 17902
rect 29150 17826 29202 17838
rect 31726 17890 31778 17902
rect 31726 17826 31778 17838
rect 42590 17890 42642 17902
rect 42590 17826 42642 17838
rect 22206 17778 22258 17790
rect 27918 17778 27970 17790
rect 31390 17778 31442 17790
rect 42702 17778 42754 17790
rect 10770 17726 10782 17778
rect 10834 17726 10846 17778
rect 12898 17726 12910 17778
rect 12962 17726 12974 17778
rect 19842 17726 19854 17778
rect 19906 17726 19918 17778
rect 20738 17726 20750 17778
rect 20802 17726 20814 17778
rect 24546 17726 24558 17778
rect 24610 17726 24622 17778
rect 26674 17726 26686 17778
rect 26738 17726 26750 17778
rect 29474 17726 29486 17778
rect 29538 17726 29550 17778
rect 32050 17726 32062 17778
rect 32114 17726 32126 17778
rect 33394 17726 33406 17778
rect 33458 17726 33470 17778
rect 6526 17714 6578 17726
rect 22206 17714 22258 17726
rect 27918 17714 27970 17726
rect 31390 17714 31442 17726
rect 42702 17714 42754 17726
rect 43374 17778 43426 17790
rect 43374 17714 43426 17726
rect 44942 17778 44994 17790
rect 44942 17714 44994 17726
rect 45390 17778 45442 17790
rect 45390 17714 45442 17726
rect 2718 17666 2770 17678
rect 2718 17602 2770 17614
rect 3054 17666 3106 17678
rect 3054 17602 3106 17614
rect 3838 17666 3890 17678
rect 3838 17602 3890 17614
rect 4174 17666 4226 17678
rect 4174 17602 4226 17614
rect 6078 17666 6130 17678
rect 14254 17666 14306 17678
rect 10098 17614 10110 17666
rect 10162 17614 10174 17666
rect 13906 17614 13918 17666
rect 13970 17614 13982 17666
rect 6078 17602 6130 17614
rect 14254 17602 14306 17614
rect 14478 17666 14530 17678
rect 22318 17666 22370 17678
rect 16034 17614 16046 17666
rect 16098 17614 16110 17666
rect 14478 17602 14530 17614
rect 22318 17602 22370 17614
rect 22766 17666 22818 17678
rect 29822 17666 29874 17678
rect 23090 17614 23102 17666
rect 23154 17614 23166 17666
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 22766 17602 22818 17614
rect 29822 17602 29874 17614
rect 30830 17666 30882 17678
rect 30830 17602 30882 17614
rect 32398 17666 32450 17678
rect 33742 17666 33794 17678
rect 34526 17666 34578 17678
rect 43262 17666 43314 17678
rect 32834 17614 32846 17666
rect 32898 17614 32910 17666
rect 33282 17614 33294 17666
rect 33346 17614 33358 17666
rect 33954 17614 33966 17666
rect 34018 17614 34030 17666
rect 36306 17614 36318 17666
rect 36370 17614 36382 17666
rect 40786 17614 40798 17666
rect 40850 17614 40862 17666
rect 43026 17614 43038 17666
rect 43090 17614 43102 17666
rect 32398 17602 32450 17614
rect 33742 17602 33794 17614
rect 34526 17602 34578 17614
rect 43262 17602 43314 17614
rect 2830 17554 2882 17566
rect 2830 17490 2882 17502
rect 5742 17554 5794 17566
rect 28590 17554 28642 17566
rect 23314 17502 23326 17554
rect 23378 17502 23390 17554
rect 5742 17490 5794 17502
rect 28590 17490 28642 17502
rect 31950 17554 32002 17566
rect 31950 17490 32002 17502
rect 34302 17554 34354 17566
rect 34302 17490 34354 17502
rect 34862 17554 34914 17566
rect 43710 17554 43762 17566
rect 35522 17502 35534 17554
rect 35586 17502 35598 17554
rect 36082 17502 36094 17554
rect 36146 17502 36158 17554
rect 37426 17502 37438 17554
rect 37490 17502 37502 17554
rect 34862 17490 34914 17502
rect 43710 17490 43762 17502
rect 46174 17554 46226 17566
rect 46174 17490 46226 17502
rect 3950 17442 4002 17454
rect 3950 17378 4002 17390
rect 14366 17442 14418 17454
rect 14366 17378 14418 17390
rect 20526 17442 20578 17454
rect 20526 17378 20578 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 22094 17442 22146 17454
rect 22094 17378 22146 17390
rect 29374 17442 29426 17454
rect 33518 17442 33570 17454
rect 30146 17390 30158 17442
rect 30210 17390 30222 17442
rect 30482 17390 30494 17442
rect 30546 17390 30558 17442
rect 29374 17378 29426 17390
rect 33518 17378 33570 17390
rect 34750 17442 34802 17454
rect 34750 17378 34802 17390
rect 35198 17442 35250 17454
rect 35198 17378 35250 17390
rect 43486 17442 43538 17454
rect 43486 17378 43538 17390
rect 44158 17442 44210 17454
rect 44158 17378 44210 17390
rect 45838 17442 45890 17454
rect 45838 17378 45890 17390
rect 1344 17274 46592 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 46592 17274
rect 1344 17188 46592 17222
rect 13246 17106 13298 17118
rect 13246 17042 13298 17054
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 20526 17106 20578 17118
rect 27694 17106 27746 17118
rect 24658 17054 24670 17106
rect 24722 17054 24734 17106
rect 20526 17042 20578 17054
rect 27694 17042 27746 17054
rect 38334 17106 38386 17118
rect 38334 17042 38386 17054
rect 38446 17106 38498 17118
rect 38446 17042 38498 17054
rect 38670 17106 38722 17118
rect 38670 17042 38722 17054
rect 39342 17106 39394 17118
rect 39342 17042 39394 17054
rect 39454 17106 39506 17118
rect 39454 17042 39506 17054
rect 41358 17106 41410 17118
rect 41358 17042 41410 17054
rect 41582 17106 41634 17118
rect 41582 17042 41634 17054
rect 42478 17106 42530 17118
rect 42478 17042 42530 17054
rect 42702 17106 42754 17118
rect 42702 17042 42754 17054
rect 12798 16994 12850 17006
rect 19742 16994 19794 17006
rect 27134 16994 27186 17006
rect 10322 16942 10334 16994
rect 10386 16942 10398 16994
rect 19506 16942 19518 16994
rect 19570 16942 19582 16994
rect 22866 16942 22878 16994
rect 22930 16942 22942 16994
rect 12798 16930 12850 16942
rect 19742 16930 19794 16942
rect 27134 16930 27186 16942
rect 28142 16994 28194 17006
rect 28142 16930 28194 16942
rect 31726 16994 31778 17006
rect 31726 16930 31778 16942
rect 33070 16994 33122 17006
rect 39230 16994 39282 17006
rect 34290 16942 34302 16994
rect 34354 16942 34366 16994
rect 35410 16942 35422 16994
rect 35474 16942 35486 16994
rect 33070 16930 33122 16942
rect 39230 16930 39282 16942
rect 39902 16994 39954 17006
rect 44034 16942 44046 16994
rect 44098 16942 44110 16994
rect 39902 16930 39954 16942
rect 13022 16882 13074 16894
rect 18286 16882 18338 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 6178 16830 6190 16882
rect 6242 16830 6254 16882
rect 9650 16830 9662 16882
rect 9714 16830 9726 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 13022 16818 13074 16830
rect 18286 16818 18338 16830
rect 19182 16882 19234 16894
rect 25454 16882 25506 16894
rect 26350 16882 26402 16894
rect 23650 16830 23662 16882
rect 23714 16830 23726 16882
rect 26114 16830 26126 16882
rect 26178 16830 26190 16882
rect 19182 16818 19234 16830
rect 25454 16818 25506 16830
rect 26350 16818 26402 16830
rect 27246 16882 27298 16894
rect 32286 16882 32338 16894
rect 38558 16882 38610 16894
rect 40014 16882 40066 16894
rect 31266 16830 31278 16882
rect 31330 16830 31342 16882
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 34066 16830 34078 16882
rect 34130 16830 34142 16882
rect 34626 16830 34638 16882
rect 34690 16830 34702 16882
rect 38882 16830 38894 16882
rect 38946 16830 38958 16882
rect 41122 16830 41134 16882
rect 41186 16830 41198 16882
rect 41794 16830 41806 16882
rect 41858 16830 41870 16882
rect 42242 16830 42254 16882
rect 42306 16830 42318 16882
rect 42914 16830 42926 16882
rect 42978 16830 42990 16882
rect 43362 16830 43374 16882
rect 43426 16830 43438 16882
rect 27246 16818 27298 16830
rect 32286 16818 32338 16830
rect 38558 16818 38610 16830
rect 40014 16818 40066 16830
rect 5518 16770 5570 16782
rect 12910 16770 12962 16782
rect 17950 16770 18002 16782
rect 2482 16718 2494 16770
rect 2546 16718 2558 16770
rect 4610 16718 4622 16770
rect 4674 16718 4686 16770
rect 6850 16718 6862 16770
rect 6914 16718 6926 16770
rect 8978 16718 8990 16770
rect 9042 16718 9054 16770
rect 12450 16718 12462 16770
rect 12514 16718 12526 16770
rect 14690 16718 14702 16770
rect 14754 16718 14766 16770
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 5518 16706 5570 16718
rect 12910 16706 12962 16718
rect 17950 16706 18002 16718
rect 18174 16770 18226 16782
rect 18174 16706 18226 16718
rect 19966 16770 20018 16782
rect 24110 16770 24162 16782
rect 20738 16718 20750 16770
rect 20802 16718 20814 16770
rect 19966 16706 20018 16718
rect 24110 16706 24162 16718
rect 24334 16770 24386 16782
rect 41470 16770 41522 16782
rect 28466 16718 28478 16770
rect 28530 16718 28542 16770
rect 30594 16718 30606 16770
rect 30658 16718 30670 16770
rect 37538 16718 37550 16770
rect 37602 16718 37614 16770
rect 24334 16706 24386 16718
rect 41470 16706 41522 16718
rect 42590 16770 42642 16782
rect 46162 16718 46174 16770
rect 46226 16718 46238 16770
rect 42590 16706 42642 16718
rect 5294 16658 5346 16670
rect 4946 16606 4958 16658
rect 5010 16606 5022 16658
rect 5294 16594 5346 16606
rect 18958 16658 19010 16670
rect 18958 16594 19010 16606
rect 27134 16658 27186 16670
rect 27134 16594 27186 16606
rect 1344 16490 46592 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 46592 16490
rect 1344 16404 46592 16438
rect 4734 16322 4786 16334
rect 11566 16322 11618 16334
rect 11218 16270 11230 16322
rect 11282 16270 11294 16322
rect 4734 16258 4786 16270
rect 11566 16258 11618 16270
rect 14926 16322 14978 16334
rect 14926 16258 14978 16270
rect 15598 16322 15650 16334
rect 15598 16258 15650 16270
rect 15934 16322 15986 16334
rect 15934 16258 15986 16270
rect 17726 16322 17778 16334
rect 17726 16258 17778 16270
rect 18398 16322 18450 16334
rect 30606 16322 30658 16334
rect 21186 16270 21198 16322
rect 21250 16319 21262 16322
rect 21410 16319 21422 16322
rect 21250 16273 21422 16319
rect 21250 16270 21262 16273
rect 21410 16270 21422 16273
rect 21474 16270 21486 16322
rect 45714 16270 45726 16322
rect 45778 16319 45790 16322
rect 46162 16319 46174 16322
rect 45778 16273 46174 16319
rect 45778 16270 45790 16273
rect 46162 16270 46174 16273
rect 46226 16270 46238 16322
rect 18398 16258 18450 16270
rect 30606 16258 30658 16270
rect 8654 16210 8706 16222
rect 8654 16146 8706 16158
rect 10558 16210 10610 16222
rect 10558 16146 10610 16158
rect 11790 16210 11842 16222
rect 11790 16146 11842 16158
rect 17950 16210 18002 16222
rect 20750 16210 20802 16222
rect 19394 16158 19406 16210
rect 19458 16158 19470 16210
rect 17950 16146 18002 16158
rect 20750 16146 20802 16158
rect 21422 16210 21474 16222
rect 21422 16146 21474 16158
rect 22990 16210 23042 16222
rect 28590 16210 28642 16222
rect 30494 16210 30546 16222
rect 24658 16158 24670 16210
rect 24722 16158 24734 16210
rect 26786 16158 26798 16210
rect 26850 16158 26862 16210
rect 30034 16158 30046 16210
rect 30098 16158 30110 16210
rect 22990 16146 23042 16158
rect 28590 16146 28642 16158
rect 30494 16146 30546 16158
rect 31390 16210 31442 16222
rect 31390 16146 31442 16158
rect 31838 16210 31890 16222
rect 31838 16146 31890 16158
rect 32062 16210 32114 16222
rect 35646 16210 35698 16222
rect 35186 16158 35198 16210
rect 35250 16158 35262 16210
rect 32062 16146 32114 16158
rect 35646 16146 35698 16158
rect 37214 16210 37266 16222
rect 44830 16210 44882 16222
rect 38210 16158 38222 16210
rect 38274 16158 38286 16210
rect 40338 16158 40350 16210
rect 40402 16158 40414 16210
rect 41458 16158 41470 16210
rect 41522 16158 41534 16210
rect 43586 16158 43598 16210
rect 43650 16158 43662 16210
rect 37214 16146 37266 16158
rect 44830 16146 44882 16158
rect 45278 16210 45330 16222
rect 45278 16146 45330 16158
rect 45838 16210 45890 16222
rect 45838 16146 45890 16158
rect 4062 16098 4114 16110
rect 4062 16034 4114 16046
rect 4286 16098 4338 16110
rect 4286 16034 4338 16046
rect 5854 16098 5906 16110
rect 5854 16034 5906 16046
rect 8878 16098 8930 16110
rect 8878 16034 8930 16046
rect 9550 16098 9602 16110
rect 9550 16034 9602 16046
rect 9774 16098 9826 16110
rect 16494 16098 16546 16110
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 9774 16034 9826 16046
rect 16494 16034 16546 16046
rect 16942 16098 16994 16110
rect 16942 16034 16994 16046
rect 17502 16098 17554 16110
rect 22430 16098 22482 16110
rect 27582 16098 27634 16110
rect 18946 16046 18958 16098
rect 19010 16046 19022 16098
rect 19170 16046 19182 16098
rect 19234 16046 19246 16098
rect 23874 16046 23886 16098
rect 23938 16046 23950 16098
rect 17502 16034 17554 16046
rect 22430 16034 22482 16046
rect 27582 16034 27634 16046
rect 27694 16098 27746 16110
rect 29710 16098 29762 16110
rect 29474 16046 29486 16098
rect 29538 16046 29550 16098
rect 27694 16034 27746 16046
rect 29710 16034 29762 16046
rect 29934 16098 29986 16110
rect 29934 16034 29986 16046
rect 32622 16098 32674 16110
rect 36094 16098 36146 16110
rect 33170 16046 33182 16098
rect 33234 16046 33246 16098
rect 33842 16046 33854 16098
rect 33906 16046 33918 16098
rect 35074 16046 35086 16098
rect 35138 16046 35150 16098
rect 37426 16046 37438 16098
rect 37490 16046 37502 16098
rect 40786 16046 40798 16098
rect 40850 16046 40862 16098
rect 32622 16034 32674 16046
rect 36094 16034 36146 16046
rect 4846 15986 4898 15998
rect 4846 15922 4898 15934
rect 5070 15986 5122 15998
rect 5070 15922 5122 15934
rect 9662 15986 9714 15998
rect 9662 15922 9714 15934
rect 10446 15986 10498 15998
rect 10446 15922 10498 15934
rect 15038 15986 15090 15998
rect 15038 15922 15090 15934
rect 15262 15986 15314 15998
rect 15262 15922 15314 15934
rect 16382 15986 16434 15998
rect 16382 15922 16434 15934
rect 20302 15986 20354 15998
rect 20302 15922 20354 15934
rect 27806 15986 27858 15998
rect 27806 15922 27858 15934
rect 30046 15986 30098 15998
rect 44046 15986 44098 15998
rect 36418 15934 36430 15986
rect 36482 15934 36494 15986
rect 30046 15922 30098 15934
rect 44046 15922 44098 15934
rect 3502 15874 3554 15886
rect 5630 15874 5682 15886
rect 3714 15822 3726 15874
rect 3778 15822 3790 15874
rect 3502 15810 3554 15822
rect 5630 15810 5682 15822
rect 5742 15874 5794 15886
rect 5742 15810 5794 15822
rect 6078 15874 6130 15886
rect 10670 15874 10722 15886
rect 9202 15822 9214 15874
rect 9266 15822 9278 15874
rect 6078 15810 6130 15822
rect 10670 15810 10722 15822
rect 15822 15874 15874 15886
rect 15822 15810 15874 15822
rect 16270 15874 16322 15886
rect 21870 15874 21922 15886
rect 28478 15874 28530 15886
rect 43934 15874 43986 15886
rect 18946 15822 18958 15874
rect 19010 15822 19022 15874
rect 27122 15822 27134 15874
rect 27186 15822 27198 15874
rect 32946 15822 32958 15874
rect 33010 15822 33022 15874
rect 33618 15822 33630 15874
rect 33682 15822 33694 15874
rect 16270 15810 16322 15822
rect 21870 15810 21922 15822
rect 28478 15810 28530 15822
rect 43934 15810 43986 15822
rect 44942 15874 44994 15886
rect 44942 15810 44994 15822
rect 45390 15874 45442 15886
rect 45390 15810 45442 15822
rect 1344 15706 46592 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 46592 15706
rect 1344 15620 46592 15654
rect 10110 15538 10162 15550
rect 14702 15538 14754 15550
rect 14354 15486 14366 15538
rect 14418 15486 14430 15538
rect 10110 15474 10162 15486
rect 14702 15474 14754 15486
rect 15038 15538 15090 15550
rect 15038 15474 15090 15486
rect 16830 15538 16882 15550
rect 16830 15474 16882 15486
rect 17614 15538 17666 15550
rect 17614 15474 17666 15486
rect 18062 15538 18114 15550
rect 18062 15474 18114 15486
rect 18174 15538 18226 15550
rect 18174 15474 18226 15486
rect 19182 15538 19234 15550
rect 19182 15474 19234 15486
rect 19294 15538 19346 15550
rect 19294 15474 19346 15486
rect 19406 15538 19458 15550
rect 19406 15474 19458 15486
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 22542 15538 22594 15550
rect 22542 15474 22594 15486
rect 26462 15538 26514 15550
rect 26462 15474 26514 15486
rect 27806 15538 27858 15550
rect 27806 15474 27858 15486
rect 28478 15538 28530 15550
rect 28478 15474 28530 15486
rect 39790 15538 39842 15550
rect 39790 15474 39842 15486
rect 17950 15426 18002 15438
rect 17950 15362 18002 15374
rect 20862 15426 20914 15438
rect 20862 15362 20914 15374
rect 27918 15426 27970 15438
rect 41122 15374 41134 15426
rect 41186 15374 41198 15426
rect 27918 15362 27970 15374
rect 10334 15314 10386 15326
rect 1810 15262 1822 15314
rect 1874 15262 1886 15314
rect 6066 15262 6078 15314
rect 6130 15262 6142 15314
rect 10334 15250 10386 15262
rect 10782 15314 10834 15326
rect 18734 15314 18786 15326
rect 19966 15314 20018 15326
rect 25342 15314 25394 15326
rect 26238 15314 26290 15326
rect 11106 15262 11118 15314
rect 11170 15262 11182 15314
rect 15250 15262 15262 15314
rect 15314 15262 15326 15314
rect 19730 15262 19742 15314
rect 19794 15262 19806 15314
rect 21074 15262 21086 15314
rect 21138 15262 21150 15314
rect 25778 15262 25790 15314
rect 25842 15262 25854 15314
rect 10782 15250 10834 15262
rect 18734 15250 18786 15262
rect 19966 15250 20018 15262
rect 25342 15250 25394 15262
rect 26238 15250 26290 15262
rect 26462 15314 26514 15326
rect 26462 15250 26514 15262
rect 26686 15314 26738 15326
rect 26686 15250 26738 15262
rect 27358 15314 27410 15326
rect 27358 15250 27410 15262
rect 27582 15314 27634 15326
rect 27582 15250 27634 15262
rect 28030 15314 28082 15326
rect 28030 15250 28082 15262
rect 28590 15314 28642 15326
rect 38670 15314 38722 15326
rect 32162 15262 32174 15314
rect 32226 15262 32238 15314
rect 37762 15262 37774 15314
rect 37826 15262 37838 15314
rect 45826 15262 45838 15314
rect 45890 15262 45902 15314
rect 28590 15250 28642 15262
rect 38670 15250 38722 15262
rect 10222 15202 10274 15214
rect 17502 15202 17554 15214
rect 2482 15150 2494 15202
rect 2546 15150 2558 15202
rect 4610 15150 4622 15202
rect 4674 15150 4686 15202
rect 6738 15150 6750 15202
rect 6802 15150 6814 15202
rect 8866 15150 8878 15202
rect 8930 15150 8942 15202
rect 11890 15150 11902 15202
rect 11954 15150 11966 15202
rect 14018 15150 14030 15202
rect 14082 15150 14094 15202
rect 10222 15138 10274 15150
rect 17502 15138 17554 15150
rect 20302 15202 20354 15214
rect 20302 15138 20354 15150
rect 22094 15202 22146 15214
rect 22094 15138 22146 15150
rect 25230 15202 25282 15214
rect 25230 15138 25282 15150
rect 25566 15202 25618 15214
rect 26898 15150 26910 15202
rect 26962 15199 26974 15202
rect 27122 15199 27134 15202
rect 26962 15153 27134 15199
rect 26962 15150 26974 15153
rect 27122 15150 27134 15153
rect 27186 15150 27198 15202
rect 29250 15150 29262 15202
rect 29314 15150 29326 15202
rect 31378 15150 31390 15202
rect 31442 15150 31454 15202
rect 33618 15150 33630 15202
rect 33682 15150 33694 15202
rect 40226 15150 40238 15202
rect 40290 15150 40302 15202
rect 25566 15138 25618 15150
rect 20190 15090 20242 15102
rect 20190 15026 20242 15038
rect 38894 15090 38946 15102
rect 39218 15038 39230 15090
rect 39282 15038 39294 15090
rect 38894 15026 38946 15038
rect 1344 14922 46592 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 46592 14922
rect 1344 14836 46592 14870
rect 3166 14754 3218 14766
rect 3166 14690 3218 14702
rect 22542 14754 22594 14766
rect 22542 14690 22594 14702
rect 26574 14754 26626 14766
rect 26574 14690 26626 14702
rect 27134 14754 27186 14766
rect 27134 14690 27186 14702
rect 4846 14642 4898 14654
rect 12014 14642 12066 14654
rect 7746 14590 7758 14642
rect 7810 14590 7822 14642
rect 9874 14590 9886 14642
rect 9938 14590 9950 14642
rect 10210 14590 10222 14642
rect 10274 14590 10286 14642
rect 4846 14578 4898 14590
rect 12014 14578 12066 14590
rect 13022 14642 13074 14654
rect 30830 14642 30882 14654
rect 15810 14590 15822 14642
rect 15874 14590 15886 14642
rect 16258 14590 16270 14642
rect 16322 14590 16334 14642
rect 18386 14590 18398 14642
rect 18450 14590 18462 14642
rect 20514 14590 20526 14642
rect 20578 14590 20590 14642
rect 23762 14590 23774 14642
rect 23826 14590 23838 14642
rect 25890 14590 25902 14642
rect 25954 14590 25966 14642
rect 30370 14590 30382 14642
rect 30434 14590 30446 14642
rect 13022 14578 13074 14590
rect 30830 14578 30882 14590
rect 30942 14642 30994 14654
rect 30942 14578 30994 14590
rect 33182 14642 33234 14654
rect 33182 14578 33234 14590
rect 36094 14642 36146 14654
rect 42702 14642 42754 14654
rect 38322 14590 38334 14642
rect 38386 14590 38398 14642
rect 36094 14578 36146 14590
rect 42702 14578 42754 14590
rect 4062 14530 4114 14542
rect 10894 14530 10946 14542
rect 4386 14478 4398 14530
rect 4450 14478 4462 14530
rect 7074 14478 7086 14530
rect 7138 14478 7150 14530
rect 4062 14466 4114 14478
rect 10894 14466 10946 14478
rect 11118 14530 11170 14542
rect 11118 14466 11170 14478
rect 11790 14530 11842 14542
rect 11790 14466 11842 14478
rect 12238 14530 12290 14542
rect 12238 14466 12290 14478
rect 13694 14530 13746 14542
rect 13694 14466 13746 14478
rect 14142 14530 14194 14542
rect 28030 14530 28082 14542
rect 29374 14530 29426 14542
rect 30046 14530 30098 14542
rect 14914 14478 14926 14530
rect 14978 14478 14990 14530
rect 15474 14478 15486 14530
rect 15538 14478 15550 14530
rect 19170 14478 19182 14530
rect 19234 14478 19246 14530
rect 21410 14478 21422 14530
rect 21474 14478 21486 14530
rect 23090 14478 23102 14530
rect 23154 14478 23166 14530
rect 28466 14478 28478 14530
rect 28530 14478 28542 14530
rect 29810 14478 29822 14530
rect 29874 14478 29886 14530
rect 14142 14466 14194 14478
rect 28030 14466 28082 14478
rect 29374 14466 29426 14478
rect 30046 14466 30098 14478
rect 32286 14530 32338 14542
rect 34526 14530 34578 14542
rect 32722 14478 32734 14530
rect 32786 14478 32798 14530
rect 32286 14466 32338 14478
rect 34526 14466 34578 14478
rect 34862 14530 34914 14542
rect 34862 14466 34914 14478
rect 35870 14530 35922 14542
rect 37214 14530 37266 14542
rect 36194 14478 36206 14530
rect 36258 14478 36270 14530
rect 35870 14466 35922 14478
rect 37214 14466 37266 14478
rect 37998 14530 38050 14542
rect 41122 14478 41134 14530
rect 41186 14478 41198 14530
rect 37998 14466 38050 14478
rect 3278 14418 3330 14430
rect 3278 14354 3330 14366
rect 3502 14418 3554 14430
rect 3502 14354 3554 14366
rect 5630 14418 5682 14430
rect 5630 14354 5682 14366
rect 5966 14418 6018 14430
rect 10334 14418 10386 14430
rect 6626 14366 6638 14418
rect 6690 14366 6702 14418
rect 5966 14354 6018 14366
rect 10334 14354 10386 14366
rect 10558 14418 10610 14430
rect 10558 14354 10610 14366
rect 12462 14418 12514 14430
rect 12462 14354 12514 14366
rect 13582 14418 13634 14430
rect 13582 14354 13634 14366
rect 19854 14418 19906 14430
rect 19854 14354 19906 14366
rect 20078 14418 20130 14430
rect 22430 14418 22482 14430
rect 21634 14366 21646 14418
rect 21698 14366 21710 14418
rect 20078 14354 20130 14366
rect 22430 14354 22482 14366
rect 27134 14418 27186 14430
rect 27134 14354 27186 14366
rect 27246 14418 27298 14430
rect 27246 14354 27298 14366
rect 27694 14418 27746 14430
rect 27694 14354 27746 14366
rect 30382 14418 30434 14430
rect 33518 14418 33570 14430
rect 31938 14366 31950 14418
rect 32002 14366 32014 14418
rect 30382 14354 30434 14366
rect 33518 14354 33570 14366
rect 33854 14418 33906 14430
rect 41694 14418 41746 14430
rect 37538 14366 37550 14418
rect 37602 14366 37614 14418
rect 37874 14366 37886 14418
rect 37938 14366 37950 14418
rect 40450 14366 40462 14418
rect 40514 14366 40526 14418
rect 33854 14354 33906 14366
rect 41694 14354 41746 14366
rect 43150 14418 43202 14430
rect 43150 14354 43202 14366
rect 43710 14418 43762 14430
rect 43710 14354 43762 14366
rect 3838 14306 3890 14318
rect 3838 14242 3890 14254
rect 3950 14306 4002 14318
rect 3950 14242 4002 14254
rect 6302 14306 6354 14318
rect 13470 14306 13522 14318
rect 11442 14254 11454 14306
rect 11506 14254 11518 14306
rect 6302 14242 6354 14254
rect 13470 14242 13522 14254
rect 14702 14306 14754 14318
rect 14702 14242 14754 14254
rect 22206 14306 22258 14318
rect 22206 14242 22258 14254
rect 22542 14306 22594 14318
rect 22542 14242 22594 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 26462 14306 26514 14318
rect 26462 14242 26514 14254
rect 29038 14306 29090 14318
rect 29038 14242 29090 14254
rect 29262 14306 29314 14318
rect 29262 14242 29314 14254
rect 30270 14306 30322 14318
rect 30270 14242 30322 14254
rect 31726 14306 31778 14318
rect 34974 14306 35026 14318
rect 34178 14254 34190 14306
rect 34242 14254 34254 14306
rect 31726 14242 31778 14254
rect 34974 14242 35026 14254
rect 35086 14306 35138 14318
rect 35086 14242 35138 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 36430 14306 36482 14318
rect 36430 14242 36482 14254
rect 36990 14306 37042 14318
rect 36990 14242 37042 14254
rect 41806 14306 41858 14318
rect 41806 14242 41858 14254
rect 42030 14306 42082 14318
rect 42030 14242 42082 14254
rect 42590 14306 42642 14318
rect 42590 14242 42642 14254
rect 43038 14306 43090 14318
rect 43038 14242 43090 14254
rect 44046 14306 44098 14318
rect 44046 14242 44098 14254
rect 44830 14306 44882 14318
rect 44830 14242 44882 14254
rect 45278 14306 45330 14318
rect 45278 14242 45330 14254
rect 45726 14306 45778 14318
rect 45726 14242 45778 14254
rect 1344 14138 46592 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 46592 14138
rect 1344 14052 46592 14086
rect 6190 13970 6242 13982
rect 7982 13970 8034 13982
rect 5842 13918 5854 13970
rect 5906 13918 5918 13970
rect 6962 13918 6974 13970
rect 7026 13918 7038 13970
rect 6190 13906 6242 13918
rect 7982 13906 8034 13918
rect 8878 13970 8930 13982
rect 10446 13970 10498 13982
rect 9538 13918 9550 13970
rect 9602 13918 9614 13970
rect 8878 13906 8930 13918
rect 10446 13906 10498 13918
rect 10558 13970 10610 13982
rect 10558 13906 10610 13918
rect 10670 13970 10722 13982
rect 10670 13906 10722 13918
rect 11454 13970 11506 13982
rect 11454 13906 11506 13918
rect 13470 13970 13522 13982
rect 13470 13906 13522 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 16158 13970 16210 13982
rect 16158 13906 16210 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 29598 13970 29650 13982
rect 29598 13906 29650 13918
rect 32174 13970 32226 13982
rect 32174 13906 32226 13918
rect 33294 13970 33346 13982
rect 33294 13906 33346 13918
rect 33742 13970 33794 13982
rect 33742 13906 33794 13918
rect 39566 13970 39618 13982
rect 42914 13918 42926 13970
rect 42978 13918 42990 13970
rect 39566 13906 39618 13918
rect 8766 13858 8818 13870
rect 8766 13794 8818 13806
rect 8990 13858 9042 13870
rect 8990 13794 9042 13806
rect 11566 13858 11618 13870
rect 11566 13794 11618 13806
rect 12126 13858 12178 13870
rect 12126 13794 12178 13806
rect 13134 13858 13186 13870
rect 23550 13858 23602 13870
rect 13794 13806 13806 13858
rect 13858 13806 13870 13858
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 15362 13806 15374 13858
rect 15426 13806 15438 13858
rect 22194 13806 22206 13858
rect 22258 13806 22270 13858
rect 13134 13794 13186 13806
rect 23550 13794 23602 13806
rect 23662 13858 23714 13870
rect 23662 13794 23714 13806
rect 26798 13858 26850 13870
rect 26798 13794 26850 13806
rect 26910 13858 26962 13870
rect 34302 13858 34354 13870
rect 38894 13858 38946 13870
rect 27682 13806 27694 13858
rect 27746 13806 27758 13858
rect 28018 13806 28030 13858
rect 28082 13806 28094 13858
rect 30258 13806 30270 13858
rect 30322 13806 30334 13858
rect 35410 13806 35422 13858
rect 35474 13806 35486 13858
rect 26910 13794 26962 13806
rect 34302 13794 34354 13806
rect 38894 13794 38946 13806
rect 39230 13858 39282 13870
rect 39230 13794 39282 13806
rect 40350 13858 40402 13870
rect 40350 13794 40402 13806
rect 41246 13858 41298 13870
rect 41246 13794 41298 13806
rect 42478 13858 42530 13870
rect 45378 13806 45390 13858
rect 45442 13806 45454 13858
rect 42478 13794 42530 13806
rect 5182 13746 5234 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 5182 13682 5234 13694
rect 7534 13746 7586 13758
rect 7534 13682 7586 13694
rect 9886 13746 9938 13758
rect 9886 13682 9938 13694
rect 10110 13746 10162 13758
rect 10110 13682 10162 13694
rect 11118 13746 11170 13758
rect 11118 13682 11170 13694
rect 12014 13746 12066 13758
rect 12014 13682 12066 13694
rect 12238 13746 12290 13758
rect 16718 13746 16770 13758
rect 24222 13746 24274 13758
rect 12562 13694 12574 13746
rect 12626 13694 12638 13746
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 14914 13694 14926 13746
rect 14978 13694 14990 13746
rect 22978 13694 22990 13746
rect 23042 13694 23054 13746
rect 12238 13682 12290 13694
rect 16718 13682 16770 13694
rect 24222 13682 24274 13694
rect 24558 13746 24610 13758
rect 24558 13682 24610 13694
rect 25566 13746 25618 13758
rect 29822 13746 29874 13758
rect 30830 13746 30882 13758
rect 40014 13746 40066 13758
rect 26562 13694 26574 13746
rect 26626 13694 26638 13746
rect 27458 13694 27470 13746
rect 27522 13694 27534 13746
rect 28466 13694 28478 13746
rect 28530 13694 28542 13746
rect 29026 13694 29038 13746
rect 29090 13694 29102 13746
rect 30034 13694 30046 13746
rect 30098 13694 30110 13746
rect 31266 13694 31278 13746
rect 31330 13694 31342 13746
rect 34066 13694 34078 13746
rect 34130 13694 34142 13746
rect 34626 13694 34638 13746
rect 34690 13694 34702 13746
rect 38434 13694 38446 13746
rect 38498 13694 38510 13746
rect 25566 13682 25618 13694
rect 29822 13682 29874 13694
rect 30830 13682 30882 13694
rect 40014 13682 40066 13694
rect 41470 13746 41522 13758
rect 42366 13746 42418 13758
rect 42130 13694 42142 13746
rect 42194 13694 42206 13746
rect 46050 13694 46062 13746
rect 46114 13694 46126 13746
rect 41470 13682 41522 13694
rect 42366 13682 42418 13694
rect 4958 13634 5010 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 4958 13570 5010 13582
rect 6750 13634 6802 13646
rect 6750 13570 6802 13582
rect 18398 13634 18450 13646
rect 25790 13634 25842 13646
rect 20066 13582 20078 13634
rect 20130 13582 20142 13634
rect 18398 13570 18450 13582
rect 25790 13570 25842 13582
rect 32510 13634 32562 13646
rect 41806 13634 41858 13646
rect 37538 13582 37550 13634
rect 37602 13582 37614 13634
rect 37986 13582 37998 13634
rect 38050 13582 38062 13634
rect 43250 13582 43262 13634
rect 43314 13582 43326 13634
rect 32510 13570 32562 13582
rect 41806 13570 41858 13582
rect 7310 13522 7362 13534
rect 5506 13470 5518 13522
rect 5570 13470 5582 13522
rect 7310 13458 7362 13470
rect 11454 13522 11506 13534
rect 11454 13458 11506 13470
rect 12910 13522 12962 13534
rect 12910 13458 12962 13470
rect 18286 13522 18338 13534
rect 18286 13458 18338 13470
rect 24446 13522 24498 13534
rect 25218 13470 25230 13522
rect 25282 13470 25294 13522
rect 24446 13458 24498 13470
rect 1344 13354 46592 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 46592 13354
rect 1344 13268 46592 13302
rect 2942 13186 2994 13198
rect 2942 13122 2994 13134
rect 4734 13186 4786 13198
rect 4734 13122 4786 13134
rect 27022 13186 27074 13198
rect 27022 13122 27074 13134
rect 38446 13186 38498 13198
rect 38446 13122 38498 13134
rect 27918 13074 27970 13086
rect 38334 13074 38386 13086
rect 8418 13022 8430 13074
rect 8482 13022 8494 13074
rect 19170 13022 19182 13074
rect 19234 13022 19246 13074
rect 23538 13022 23550 13074
rect 23602 13022 23614 13074
rect 29698 13022 29710 13074
rect 29762 13022 29774 13074
rect 34290 13022 34302 13074
rect 34354 13022 34366 13074
rect 36418 13022 36430 13074
rect 36482 13022 36494 13074
rect 27918 13010 27970 13022
rect 38334 13010 38386 13022
rect 38782 13074 38834 13086
rect 42354 13022 42366 13074
rect 42418 13022 42430 13074
rect 38782 13010 38834 13022
rect 3838 12962 3890 12974
rect 3838 12898 3890 12910
rect 4510 12962 4562 12974
rect 4510 12898 4562 12910
rect 5630 12962 5682 12974
rect 5630 12898 5682 12910
rect 5854 12962 5906 12974
rect 14254 12962 14306 12974
rect 27358 12962 27410 12974
rect 27806 12962 27858 12974
rect 12898 12910 12910 12962
rect 12962 12910 12974 12962
rect 13682 12910 13694 12962
rect 13746 12910 13758 12962
rect 16370 12910 16382 12962
rect 16434 12910 16446 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 27682 12910 27694 12962
rect 27746 12910 27758 12962
rect 5854 12898 5906 12910
rect 14254 12898 14306 12910
rect 27358 12898 27410 12910
rect 27806 12898 27858 12910
rect 28030 12962 28082 12974
rect 36878 12962 36930 12974
rect 32610 12910 32622 12962
rect 32674 12910 32686 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 28030 12898 28082 12910
rect 36878 12898 36930 12910
rect 37214 12962 37266 12974
rect 37214 12898 37266 12910
rect 37998 12962 38050 12974
rect 37998 12898 38050 12910
rect 40686 12962 40738 12974
rect 43150 12962 43202 12974
rect 41122 12910 41134 12962
rect 41186 12910 41198 12962
rect 41346 12910 41358 12962
rect 41410 12910 41422 12962
rect 42466 12910 42478 12962
rect 42530 12910 42542 12962
rect 40686 12898 40738 12910
rect 43150 12898 43202 12910
rect 43486 12962 43538 12974
rect 43486 12898 43538 12910
rect 43710 12962 43762 12974
rect 46050 12910 46062 12962
rect 46114 12910 46126 12962
rect 43710 12898 43762 12910
rect 3054 12850 3106 12862
rect 3054 12786 3106 12798
rect 3278 12850 3330 12862
rect 3278 12786 3330 12798
rect 3726 12850 3778 12862
rect 3726 12786 3778 12798
rect 6078 12850 6130 12862
rect 19518 12850 19570 12862
rect 17042 12798 17054 12850
rect 17106 12798 17118 12850
rect 6078 12786 6130 12798
rect 19518 12786 19570 12798
rect 26910 12850 26962 12862
rect 26910 12786 26962 12798
rect 28590 12850 28642 12862
rect 28590 12786 28642 12798
rect 29262 12850 29314 12862
rect 29262 12786 29314 12798
rect 29374 12850 29426 12862
rect 37550 12850 37602 12862
rect 31826 12798 31838 12850
rect 31890 12798 31902 12850
rect 29374 12786 29426 12798
rect 37550 12786 37602 12798
rect 39342 12850 39394 12862
rect 39342 12786 39394 12798
rect 39902 12850 39954 12862
rect 39902 12786 39954 12798
rect 40350 12850 40402 12862
rect 40350 12786 40402 12798
rect 40798 12850 40850 12862
rect 40798 12786 40850 12798
rect 45502 12850 45554 12862
rect 45826 12798 45838 12850
rect 45890 12798 45902 12850
rect 45502 12786 45554 12798
rect 3614 12738 3666 12750
rect 3614 12674 3666 12686
rect 4062 12738 4114 12750
rect 5742 12738 5794 12750
rect 5058 12686 5070 12738
rect 5122 12686 5134 12738
rect 4062 12674 4114 12686
rect 5742 12674 5794 12686
rect 13470 12738 13522 12750
rect 13470 12674 13522 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 19854 12738 19906 12750
rect 19854 12674 19906 12686
rect 20750 12738 20802 12750
rect 20750 12674 20802 12686
rect 33182 12738 33234 12750
rect 33182 12674 33234 12686
rect 37214 12738 37266 12750
rect 37214 12674 37266 12686
rect 37886 12738 37938 12750
rect 37886 12674 37938 12686
rect 38894 12738 38946 12750
rect 38894 12674 38946 12686
rect 39230 12738 39282 12750
rect 39230 12674 39282 12686
rect 39790 12738 39842 12750
rect 39790 12674 39842 12686
rect 40238 12738 40290 12750
rect 40238 12674 40290 12686
rect 41582 12738 41634 12750
rect 41582 12674 41634 12686
rect 41694 12738 41746 12750
rect 45166 12738 45218 12750
rect 44034 12686 44046 12738
rect 44098 12686 44110 12738
rect 41694 12674 41746 12686
rect 45166 12674 45218 12686
rect 1344 12570 46592 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 46592 12570
rect 1344 12484 46592 12518
rect 5630 12402 5682 12414
rect 5630 12338 5682 12350
rect 9662 12402 9714 12414
rect 9662 12338 9714 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 15934 12402 15986 12414
rect 15934 12338 15986 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 17838 12402 17890 12414
rect 17838 12338 17890 12350
rect 18174 12402 18226 12414
rect 18174 12338 18226 12350
rect 21086 12402 21138 12414
rect 30158 12402 30210 12414
rect 21634 12350 21646 12402
rect 21698 12350 21710 12402
rect 21086 12338 21138 12350
rect 30158 12338 30210 12350
rect 30270 12402 30322 12414
rect 30270 12338 30322 12350
rect 30494 12402 30546 12414
rect 30494 12338 30546 12350
rect 33518 12402 33570 12414
rect 39118 12402 39170 12414
rect 34402 12350 34414 12402
rect 34466 12350 34478 12402
rect 33518 12338 33570 12350
rect 39118 12338 39170 12350
rect 5518 12290 5570 12302
rect 16270 12290 16322 12302
rect 7298 12238 7310 12290
rect 7362 12238 7374 12290
rect 13458 12238 13470 12290
rect 13522 12238 13534 12290
rect 5518 12226 5570 12238
rect 16270 12226 16322 12238
rect 16606 12290 16658 12302
rect 16606 12226 16658 12238
rect 18398 12290 18450 12302
rect 18398 12226 18450 12238
rect 18846 12290 18898 12302
rect 21982 12290 22034 12302
rect 19282 12238 19294 12290
rect 19346 12238 19358 12290
rect 20402 12238 20414 12290
rect 20466 12238 20478 12290
rect 18846 12226 18898 12238
rect 21982 12226 22034 12238
rect 23998 12290 24050 12302
rect 23998 12226 24050 12238
rect 27134 12290 27186 12302
rect 27134 12226 27186 12238
rect 27246 12290 27298 12302
rect 27246 12226 27298 12238
rect 27694 12290 27746 12302
rect 27694 12226 27746 12238
rect 27806 12290 27858 12302
rect 27806 12226 27858 12238
rect 28926 12290 28978 12302
rect 28926 12226 28978 12238
rect 29150 12290 29202 12302
rect 29150 12226 29202 12238
rect 29934 12290 29986 12302
rect 29934 12226 29986 12238
rect 34862 12290 34914 12302
rect 34862 12226 34914 12238
rect 34974 12290 35026 12302
rect 34974 12226 35026 12238
rect 35086 12290 35138 12302
rect 41358 12290 41410 12302
rect 35746 12238 35758 12290
rect 35810 12238 35822 12290
rect 36642 12238 36654 12290
rect 36706 12238 36718 12290
rect 40114 12238 40126 12290
rect 40178 12238 40190 12290
rect 35086 12226 35138 12238
rect 41358 12226 41410 12238
rect 42366 12290 42418 12302
rect 42366 12226 42418 12238
rect 42814 12290 42866 12302
rect 45378 12238 45390 12290
rect 45442 12238 45454 12290
rect 42814 12226 42866 12238
rect 5742 12178 5794 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 5742 12114 5794 12126
rect 6190 12178 6242 12190
rect 6190 12114 6242 12126
rect 6414 12178 6466 12190
rect 6414 12114 6466 12126
rect 6638 12178 6690 12190
rect 6638 12114 6690 12126
rect 7086 12178 7138 12190
rect 16942 12178 16994 12190
rect 7522 12126 7534 12178
rect 7586 12126 7598 12178
rect 11330 12126 11342 12178
rect 11394 12126 11406 12178
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 7086 12114 7138 12126
rect 16942 12114 16994 12126
rect 17390 12178 17442 12190
rect 17390 12114 17442 12126
rect 17726 12178 17778 12190
rect 17726 12114 17778 12126
rect 18062 12178 18114 12190
rect 18062 12114 18114 12126
rect 18510 12178 18562 12190
rect 22878 12178 22930 12190
rect 23886 12178 23938 12190
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 20066 12126 20078 12178
rect 20130 12126 20142 12178
rect 21410 12126 21422 12178
rect 21474 12126 21486 12178
rect 22418 12126 22430 12178
rect 22482 12126 22494 12178
rect 23650 12126 23662 12178
rect 23714 12126 23726 12178
rect 18510 12114 18562 12126
rect 22878 12114 22930 12126
rect 23886 12114 23938 12126
rect 24110 12178 24162 12190
rect 24110 12114 24162 12126
rect 25342 12178 25394 12190
rect 25342 12114 25394 12126
rect 25566 12178 25618 12190
rect 25566 12114 25618 12126
rect 25790 12178 25842 12190
rect 25790 12114 25842 12126
rect 26462 12178 26514 12190
rect 26462 12114 26514 12126
rect 26910 12178 26962 12190
rect 26910 12114 26962 12126
rect 28030 12178 28082 12190
rect 28030 12114 28082 12126
rect 29374 12178 29426 12190
rect 30382 12178 30434 12190
rect 33294 12178 33346 12190
rect 41134 12178 41186 12190
rect 29586 12126 29598 12178
rect 29650 12126 29662 12178
rect 33058 12126 33070 12178
rect 33122 12126 33134 12178
rect 33730 12126 33742 12178
rect 33794 12126 33806 12178
rect 35970 12126 35982 12178
rect 36034 12126 36046 12178
rect 36418 12126 36430 12178
rect 36482 12126 36494 12178
rect 37314 12126 37326 12178
rect 37378 12126 37390 12178
rect 39442 12126 39454 12178
rect 39506 12126 39518 12178
rect 40002 12126 40014 12178
rect 40066 12126 40078 12178
rect 29374 12114 29426 12126
rect 30382 12114 30434 12126
rect 33294 12114 33346 12126
rect 41134 12114 41186 12126
rect 41246 12178 41298 12190
rect 41246 12114 41298 12126
rect 41806 12178 41858 12190
rect 46050 12126 46062 12178
rect 46114 12126 46126 12178
rect 41806 12114 41858 12126
rect 6862 12066 6914 12078
rect 10334 12066 10386 12078
rect 2482 12014 2494 12066
rect 2546 12014 2558 12066
rect 4610 12014 4622 12066
rect 4674 12014 4686 12066
rect 10098 12014 10110 12066
rect 10162 12014 10174 12066
rect 6862 12002 6914 12014
rect 10334 12002 10386 12014
rect 10670 12066 10722 12078
rect 25678 12066 25730 12078
rect 11442 12014 11454 12066
rect 11506 12014 11518 12066
rect 15586 12014 15598 12066
rect 15650 12014 15662 12066
rect 10670 12002 10722 12014
rect 25678 12002 25730 12014
rect 26126 12066 26178 12078
rect 26126 12002 26178 12014
rect 26686 12066 26738 12078
rect 26686 12002 26738 12014
rect 28478 12066 28530 12078
rect 28478 12002 28530 12014
rect 29262 12066 29314 12078
rect 29262 12002 29314 12014
rect 31054 12066 31106 12078
rect 31054 12002 31106 12014
rect 31502 12066 31554 12078
rect 31502 12002 31554 12014
rect 32174 12066 32226 12078
rect 32174 12002 32226 12014
rect 32398 12066 32450 12078
rect 38110 12066 38162 12078
rect 33170 12014 33182 12066
rect 33234 12014 33246 12066
rect 35634 12014 35646 12066
rect 35698 12014 35710 12066
rect 39666 12014 39678 12066
rect 39730 12014 39742 12066
rect 43250 12014 43262 12066
rect 43314 12014 43326 12066
rect 32398 12002 32450 12014
rect 38110 12002 38162 12014
rect 23214 11954 23266 11966
rect 23214 11890 23266 11902
rect 28590 11954 28642 11966
rect 32510 11954 32562 11966
rect 30818 11902 30830 11954
rect 30882 11951 30894 11954
rect 31266 11951 31278 11954
rect 30882 11905 31278 11951
rect 30882 11902 30894 11905
rect 31266 11902 31278 11905
rect 31330 11951 31342 11954
rect 31490 11951 31502 11954
rect 31330 11905 31502 11951
rect 31330 11902 31342 11905
rect 31490 11902 31502 11905
rect 31554 11951 31566 11954
rect 31714 11951 31726 11954
rect 31554 11905 31726 11951
rect 31554 11902 31566 11905
rect 31714 11902 31726 11905
rect 31778 11902 31790 11954
rect 28590 11890 28642 11902
rect 32510 11890 32562 11902
rect 38222 11954 38274 11966
rect 38222 11890 38274 11902
rect 42030 11954 42082 11966
rect 42030 11890 42082 11902
rect 1344 11786 46592 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 46592 11786
rect 1344 11700 46592 11734
rect 18734 11618 18786 11630
rect 18734 11554 18786 11566
rect 27582 11618 27634 11630
rect 27582 11554 27634 11566
rect 41582 11618 41634 11630
rect 41582 11554 41634 11566
rect 42926 11618 42978 11630
rect 42926 11554 42978 11566
rect 17166 11506 17218 11518
rect 6066 11454 6078 11506
rect 6130 11454 6142 11506
rect 10098 11454 10110 11506
rect 10162 11454 10174 11506
rect 12226 11454 12238 11506
rect 12290 11454 12302 11506
rect 12562 11454 12574 11506
rect 12626 11454 12638 11506
rect 17166 11442 17218 11454
rect 19070 11506 19122 11518
rect 35086 11506 35138 11518
rect 20178 11454 20190 11506
rect 20242 11454 20254 11506
rect 24546 11454 24558 11506
rect 24610 11454 24622 11506
rect 26674 11454 26686 11506
rect 26738 11454 26750 11506
rect 34514 11454 34526 11506
rect 34578 11503 34590 11506
rect 34850 11503 34862 11506
rect 34578 11457 34862 11503
rect 34578 11454 34590 11457
rect 34850 11454 34862 11457
rect 34914 11454 34926 11506
rect 19070 11442 19122 11454
rect 35086 11442 35138 11454
rect 37102 11506 37154 11518
rect 41358 11506 41410 11518
rect 37762 11454 37774 11506
rect 37826 11454 37838 11506
rect 38770 11454 38782 11506
rect 38834 11454 38846 11506
rect 40674 11454 40686 11506
rect 40738 11454 40750 11506
rect 37102 11442 37154 11454
rect 41358 11442 41410 11454
rect 4846 11394 4898 11406
rect 4846 11330 4898 11342
rect 5070 11394 5122 11406
rect 15598 11394 15650 11406
rect 8866 11342 8878 11394
rect 8930 11342 8942 11394
rect 9314 11342 9326 11394
rect 9378 11342 9390 11394
rect 5070 11330 5122 11342
rect 15598 11330 15650 11342
rect 16270 11394 16322 11406
rect 19294 11394 19346 11406
rect 21646 11394 21698 11406
rect 28366 11394 28418 11406
rect 18386 11342 18398 11394
rect 18450 11342 18462 11394
rect 20290 11342 20302 11394
rect 20354 11342 20366 11394
rect 23762 11342 23774 11394
rect 23826 11342 23838 11394
rect 16270 11330 16322 11342
rect 19294 11330 19346 11342
rect 21646 11330 21698 11342
rect 28366 11330 28418 11342
rect 28590 11394 28642 11406
rect 35870 11394 35922 11406
rect 34402 11342 34414 11394
rect 34466 11342 34478 11394
rect 28590 11330 28642 11342
rect 35870 11330 35922 11342
rect 36206 11394 36258 11406
rect 39006 11394 39058 11406
rect 38210 11342 38222 11394
rect 38274 11342 38286 11394
rect 38546 11342 38558 11394
rect 38610 11342 38622 11394
rect 36206 11330 36258 11342
rect 39006 11330 39058 11342
rect 39118 11394 39170 11406
rect 39118 11330 39170 11342
rect 39454 11394 39506 11406
rect 42366 11394 42418 11406
rect 41906 11342 41918 11394
rect 41970 11342 41982 11394
rect 39454 11330 39506 11342
rect 42366 11330 42418 11342
rect 42478 11394 42530 11406
rect 42478 11330 42530 11342
rect 42702 11394 42754 11406
rect 42702 11330 42754 11342
rect 43038 11394 43090 11406
rect 44830 11394 44882 11406
rect 43810 11342 43822 11394
rect 43874 11342 43886 11394
rect 43038 11330 43090 11342
rect 44830 11330 44882 11342
rect 4510 11282 4562 11294
rect 12910 11282 12962 11294
rect 8194 11230 8206 11282
rect 8258 11230 8270 11282
rect 4510 11218 4562 11230
rect 12910 11218 12962 11230
rect 13358 11282 13410 11294
rect 13358 11218 13410 11230
rect 13582 11282 13634 11294
rect 13582 11218 13634 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 15262 11282 15314 11294
rect 15262 11218 15314 11230
rect 15374 11282 15426 11294
rect 15374 11218 15426 11230
rect 19966 11282 20018 11294
rect 19966 11218 20018 11230
rect 27694 11282 27746 11294
rect 35982 11282 36034 11294
rect 31266 11230 31278 11282
rect 31330 11230 31342 11282
rect 27694 11218 27746 11230
rect 35982 11218 36034 11230
rect 40126 11282 40178 11294
rect 40126 11218 40178 11230
rect 41022 11282 41074 11294
rect 41022 11218 41074 11230
rect 4622 11170 4674 11182
rect 4622 11106 4674 11118
rect 12686 11170 12738 11182
rect 12686 11106 12738 11118
rect 14926 11170 14978 11182
rect 14926 11106 14978 11118
rect 15150 11170 15202 11182
rect 15150 11106 15202 11118
rect 16046 11170 16098 11182
rect 16046 11106 16098 11118
rect 16158 11170 16210 11182
rect 16158 11106 16210 11118
rect 18622 11170 18674 11182
rect 22430 11170 22482 11182
rect 19618 11118 19630 11170
rect 19682 11118 19694 11170
rect 21298 11118 21310 11170
rect 21362 11118 21374 11170
rect 18622 11106 18674 11118
rect 22430 11106 22482 11118
rect 27246 11170 27298 11182
rect 35198 11170 35250 11182
rect 28018 11118 28030 11170
rect 28082 11118 28094 11170
rect 27246 11106 27298 11118
rect 35198 11106 35250 11118
rect 37214 11170 37266 11182
rect 37214 11106 37266 11118
rect 37662 11170 37714 11182
rect 37662 11106 37714 11118
rect 37774 11170 37826 11182
rect 37774 11106 37826 11118
rect 37998 11170 38050 11182
rect 37998 11106 38050 11118
rect 38782 11170 38834 11182
rect 38782 11106 38834 11118
rect 39902 11170 39954 11182
rect 39902 11106 39954 11118
rect 40014 11170 40066 11182
rect 40014 11106 40066 11118
rect 40798 11170 40850 11182
rect 40798 11106 40850 11118
rect 43598 11170 43650 11182
rect 43598 11106 43650 11118
rect 45166 11170 45218 11182
rect 46174 11170 46226 11182
rect 45826 11118 45838 11170
rect 45890 11118 45902 11170
rect 45166 11106 45218 11118
rect 46174 11106 46226 11118
rect 1344 11002 46592 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 46592 11002
rect 1344 10916 46592 10950
rect 5406 10834 5458 10846
rect 5406 10770 5458 10782
rect 17390 10834 17442 10846
rect 17390 10770 17442 10782
rect 31950 10834 32002 10846
rect 31950 10770 32002 10782
rect 32062 10834 32114 10846
rect 32062 10770 32114 10782
rect 32286 10834 32338 10846
rect 32286 10770 32338 10782
rect 36430 10834 36482 10846
rect 36430 10770 36482 10782
rect 36542 10834 36594 10846
rect 36542 10770 36594 10782
rect 38334 10834 38386 10846
rect 38334 10770 38386 10782
rect 39454 10834 39506 10846
rect 39454 10770 39506 10782
rect 41470 10834 41522 10846
rect 41470 10770 41522 10782
rect 5630 10722 5682 10734
rect 2818 10670 2830 10722
rect 2882 10670 2894 10722
rect 5630 10658 5682 10670
rect 6414 10722 6466 10734
rect 6414 10658 6466 10670
rect 6526 10722 6578 10734
rect 6526 10658 6578 10670
rect 8094 10722 8146 10734
rect 8094 10658 8146 10670
rect 8542 10722 8594 10734
rect 8542 10658 8594 10670
rect 11230 10722 11282 10734
rect 15486 10722 15538 10734
rect 12562 10670 12574 10722
rect 12626 10670 12638 10722
rect 11230 10658 11282 10670
rect 15486 10658 15538 10670
rect 16046 10722 16098 10734
rect 32510 10722 32562 10734
rect 36654 10722 36706 10734
rect 19058 10670 19070 10722
rect 19122 10670 19134 10722
rect 26002 10670 26014 10722
rect 26066 10670 26078 10722
rect 30594 10670 30606 10722
rect 30658 10670 30670 10722
rect 33842 10670 33854 10722
rect 33906 10670 33918 10722
rect 16046 10658 16098 10670
rect 32510 10658 32562 10670
rect 36654 10658 36706 10670
rect 37438 10722 37490 10734
rect 37438 10658 37490 10670
rect 38222 10722 38274 10734
rect 38222 10658 38274 10670
rect 39230 10722 39282 10734
rect 39230 10658 39282 10670
rect 40014 10722 40066 10734
rect 42354 10670 42366 10722
rect 42418 10670 42430 10722
rect 45378 10670 45390 10722
rect 45442 10670 45454 10722
rect 40014 10658 40066 10670
rect 7758 10610 7810 10622
rect 2034 10558 2046 10610
rect 2098 10558 2110 10610
rect 6178 10558 6190 10610
rect 6242 10558 6254 10610
rect 7758 10546 7810 10558
rect 7982 10610 8034 10622
rect 7982 10546 8034 10558
rect 10894 10610 10946 10622
rect 10894 10546 10946 10558
rect 11454 10610 11506 10622
rect 15822 10610 15874 10622
rect 11890 10558 11902 10610
rect 11954 10558 11966 10610
rect 11454 10546 11506 10558
rect 15822 10546 15874 10558
rect 17502 10610 17554 10622
rect 37102 10610 37154 10622
rect 39566 10610 39618 10622
rect 18386 10558 18398 10610
rect 18450 10558 18462 10610
rect 21634 10558 21646 10610
rect 21698 10558 21710 10610
rect 25330 10558 25342 10610
rect 25394 10558 25406 10610
rect 31266 10558 31278 10610
rect 31330 10558 31342 10610
rect 33058 10558 33070 10610
rect 33122 10558 33134 10610
rect 36754 10558 36766 10610
rect 36818 10558 36830 10610
rect 37762 10558 37774 10610
rect 37826 10558 37838 10610
rect 41234 10558 41246 10610
rect 41298 10558 41310 10610
rect 42578 10558 42590 10610
rect 42642 10558 42654 10610
rect 46050 10558 46062 10610
rect 46114 10558 46126 10610
rect 17502 10546 17554 10558
rect 37102 10546 37154 10558
rect 39566 10546 39618 10558
rect 11006 10498 11058 10510
rect 15038 10498 15090 10510
rect 4946 10446 4958 10498
rect 5010 10446 5022 10498
rect 5282 10446 5294 10498
rect 5346 10446 5358 10498
rect 14690 10446 14702 10498
rect 14754 10446 14766 10498
rect 11006 10434 11058 10446
rect 15038 10434 15090 10446
rect 15598 10498 15650 10510
rect 32174 10498 32226 10510
rect 38894 10498 38946 10510
rect 21186 10446 21198 10498
rect 21250 10446 21262 10498
rect 22306 10446 22318 10498
rect 22370 10446 22382 10498
rect 24434 10446 24446 10498
rect 24498 10446 24510 10498
rect 28130 10446 28142 10498
rect 28194 10446 28206 10498
rect 28466 10446 28478 10498
rect 28530 10446 28542 10498
rect 35970 10446 35982 10498
rect 36034 10446 36046 10498
rect 37650 10446 37662 10498
rect 37714 10446 37726 10498
rect 42018 10446 42030 10498
rect 42082 10446 42094 10498
rect 43250 10446 43262 10498
rect 43314 10446 43326 10498
rect 15598 10434 15650 10446
rect 32174 10434 32226 10446
rect 38894 10434 38946 10446
rect 7646 10386 7698 10398
rect 6962 10334 6974 10386
rect 7026 10334 7038 10386
rect 7646 10322 7698 10334
rect 15150 10386 15202 10398
rect 15150 10322 15202 10334
rect 38334 10386 38386 10398
rect 38334 10322 38386 10334
rect 39006 10386 39058 10398
rect 39006 10322 39058 10334
rect 39902 10386 39954 10398
rect 39902 10322 39954 10334
rect 40238 10386 40290 10398
rect 40238 10322 40290 10334
rect 1344 10218 46592 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 46592 10218
rect 1344 10132 46592 10166
rect 42926 10050 42978 10062
rect 42926 9986 42978 9998
rect 12014 9938 12066 9950
rect 4610 9886 4622 9938
rect 4674 9886 4686 9938
rect 9426 9886 9438 9938
rect 9490 9886 9502 9938
rect 11554 9886 11566 9938
rect 11618 9886 11630 9938
rect 12014 9874 12066 9886
rect 14478 9938 14530 9950
rect 27694 9938 27746 9950
rect 15586 9886 15598 9938
rect 15650 9886 15662 9938
rect 17714 9886 17726 9938
rect 17778 9886 17790 9938
rect 23314 9886 23326 9938
rect 23378 9886 23390 9938
rect 24210 9886 24222 9938
rect 24274 9886 24286 9938
rect 14478 9874 14530 9886
rect 27694 9874 27746 9886
rect 28590 9938 28642 9950
rect 32510 9938 32562 9950
rect 32050 9886 32062 9938
rect 32114 9886 32126 9938
rect 28590 9874 28642 9886
rect 32510 9874 32562 9886
rect 32958 9938 33010 9950
rect 42142 9938 42194 9950
rect 33282 9886 33294 9938
rect 33346 9886 33358 9938
rect 35410 9886 35422 9938
rect 35474 9886 35486 9938
rect 32958 9874 33010 9886
rect 42142 9874 42194 9886
rect 7086 9826 7138 9838
rect 11902 9826 11954 9838
rect 21646 9826 21698 9838
rect 1810 9774 1822 9826
rect 1874 9774 1886 9826
rect 8754 9774 8766 9826
rect 8818 9774 8830 9826
rect 14802 9774 14814 9826
rect 14866 9774 14878 9826
rect 7086 9762 7138 9774
rect 11902 9762 11954 9774
rect 21646 9762 21698 9774
rect 22990 9826 23042 9838
rect 40462 9826 40514 9838
rect 27122 9774 27134 9826
rect 27186 9774 27198 9826
rect 29250 9774 29262 9826
rect 29314 9774 29326 9826
rect 36082 9774 36094 9826
rect 36146 9774 36158 9826
rect 38882 9774 38894 9826
rect 38946 9774 38958 9826
rect 39442 9774 39454 9826
rect 39506 9774 39518 9826
rect 40002 9774 40014 9826
rect 40066 9774 40078 9826
rect 22990 9762 23042 9774
rect 40462 9762 40514 9774
rect 40798 9826 40850 9838
rect 40798 9762 40850 9774
rect 41022 9826 41074 9838
rect 41022 9762 41074 9774
rect 41694 9826 41746 9838
rect 41694 9762 41746 9774
rect 42366 9826 42418 9838
rect 42366 9762 42418 9774
rect 42702 9826 42754 9838
rect 42702 9762 42754 9774
rect 12350 9714 12402 9726
rect 2482 9662 2494 9714
rect 2546 9662 2558 9714
rect 12350 9650 12402 9662
rect 13470 9714 13522 9726
rect 13470 9650 13522 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 18398 9714 18450 9726
rect 18398 9650 18450 9662
rect 20638 9714 20690 9726
rect 20638 9650 20690 9662
rect 22654 9714 22706 9726
rect 22654 9650 22706 9662
rect 23662 9714 23714 9726
rect 38334 9714 38386 9726
rect 26338 9662 26350 9714
rect 26402 9662 26414 9714
rect 29922 9662 29934 9714
rect 29986 9662 29998 9714
rect 23662 9650 23714 9662
rect 38334 9650 38386 9662
rect 38670 9714 38722 9726
rect 45166 9714 45218 9726
rect 38994 9662 39006 9714
rect 39058 9662 39070 9714
rect 43250 9662 43262 9714
rect 43314 9662 43326 9714
rect 38670 9650 38722 9662
rect 45166 9650 45218 9662
rect 46174 9714 46226 9726
rect 46174 9650 46226 9662
rect 7534 9602 7586 9614
rect 7534 9538 7586 9550
rect 7646 9602 7698 9614
rect 7646 9538 7698 9550
rect 7758 9602 7810 9614
rect 7758 9538 7810 9550
rect 12126 9602 12178 9614
rect 12126 9538 12178 9550
rect 18174 9602 18226 9614
rect 18174 9538 18226 9550
rect 18286 9602 18338 9614
rect 18286 9538 18338 9550
rect 20750 9602 20802 9614
rect 20750 9538 20802 9550
rect 22206 9602 22258 9614
rect 22206 9538 22258 9550
rect 23438 9602 23490 9614
rect 23438 9538 23490 9550
rect 28142 9602 28194 9614
rect 28142 9538 28194 9550
rect 37102 9602 37154 9614
rect 37102 9538 37154 9550
rect 37886 9602 37938 9614
rect 37886 9538 37938 9550
rect 38222 9602 38274 9614
rect 38222 9538 38274 9550
rect 40686 9602 40738 9614
rect 40686 9538 40738 9550
rect 41806 9602 41858 9614
rect 41806 9538 41858 9550
rect 41918 9602 41970 9614
rect 43934 9602 43986 9614
rect 43586 9550 43598 9602
rect 43650 9550 43662 9602
rect 41918 9538 41970 9550
rect 43934 9538 43986 9550
rect 44830 9602 44882 9614
rect 44830 9538 44882 9550
rect 45838 9602 45890 9614
rect 45838 9538 45890 9550
rect 1344 9434 46592 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 46592 9434
rect 1344 9348 46592 9382
rect 2270 9266 2322 9278
rect 2270 9202 2322 9214
rect 11230 9266 11282 9278
rect 11230 9202 11282 9214
rect 13022 9266 13074 9278
rect 13022 9202 13074 9214
rect 14702 9266 14754 9278
rect 16606 9266 16658 9278
rect 16034 9214 16046 9266
rect 16098 9214 16110 9266
rect 14702 9202 14754 9214
rect 2718 9154 2770 9166
rect 2718 9090 2770 9102
rect 10110 9154 10162 9166
rect 10110 9090 10162 9102
rect 11342 9154 11394 9166
rect 11342 9090 11394 9102
rect 11902 9154 11954 9166
rect 14030 9154 14082 9166
rect 15150 9154 15202 9166
rect 12114 9102 12126 9154
rect 12178 9102 12190 9154
rect 14354 9102 14366 9154
rect 14418 9102 14430 9154
rect 15698 9102 15710 9154
rect 15762 9151 15774 9154
rect 16049 9151 16095 9214
rect 16606 9202 16658 9214
rect 24782 9266 24834 9278
rect 24782 9202 24834 9214
rect 26574 9266 26626 9278
rect 26574 9202 26626 9214
rect 27134 9266 27186 9278
rect 27134 9202 27186 9214
rect 27470 9266 27522 9278
rect 27470 9202 27522 9214
rect 27918 9266 27970 9278
rect 27918 9202 27970 9214
rect 28814 9266 28866 9278
rect 28814 9202 28866 9214
rect 30494 9266 30546 9278
rect 30494 9202 30546 9214
rect 33630 9266 33682 9278
rect 33630 9202 33682 9214
rect 39342 9266 39394 9278
rect 39342 9202 39394 9214
rect 39566 9266 39618 9278
rect 39566 9202 39618 9214
rect 39902 9266 39954 9278
rect 39902 9202 39954 9214
rect 41134 9266 41186 9278
rect 41134 9202 41186 9214
rect 41358 9266 41410 9278
rect 41358 9202 41410 9214
rect 41470 9266 41522 9278
rect 41470 9202 41522 9214
rect 15762 9105 16095 9151
rect 25790 9154 25842 9166
rect 15762 9102 15774 9105
rect 11902 9090 11954 9102
rect 14030 9090 14082 9102
rect 15150 9090 15202 9102
rect 25790 9090 25842 9102
rect 26014 9154 26066 9166
rect 26014 9090 26066 9102
rect 30158 9154 30210 9166
rect 30158 9090 30210 9102
rect 30606 9154 30658 9166
rect 30606 9090 30658 9102
rect 39118 9154 39170 9166
rect 39118 9090 39170 9102
rect 40910 9154 40962 9166
rect 45378 9102 45390 9154
rect 45442 9102 45454 9154
rect 40910 9090 40962 9102
rect 9438 9042 9490 9054
rect 8530 8990 8542 9042
rect 8594 8990 8606 9042
rect 9438 8978 9490 8990
rect 9774 9042 9826 9054
rect 9774 8978 9826 8990
rect 11790 9042 11842 9054
rect 12686 9042 12738 9054
rect 12226 8990 12238 9042
rect 12290 8990 12302 9042
rect 11790 8978 11842 8990
rect 12686 8978 12738 8990
rect 13694 9042 13746 9054
rect 13694 8978 13746 8990
rect 15486 9042 15538 9054
rect 33406 9042 33458 9054
rect 37550 9042 37602 9054
rect 15698 8990 15710 9042
rect 15762 8990 15774 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 23538 8990 23550 9042
rect 23602 8990 23614 9042
rect 25218 8990 25230 9042
rect 25282 8990 25294 9042
rect 25554 8990 25566 9042
rect 25618 8990 25630 9042
rect 31378 8990 31390 9042
rect 31442 8990 31454 9042
rect 33170 8990 33182 9042
rect 33234 8990 33246 9042
rect 33842 8990 33854 9042
rect 33906 8990 33918 9042
rect 34290 8990 34302 9042
rect 34354 8990 34366 9042
rect 15486 8978 15538 8990
rect 33406 8978 33458 8990
rect 37550 8978 37602 8990
rect 37998 9042 38050 9054
rect 42814 9042 42866 9054
rect 40114 8990 40126 9042
rect 40178 8990 40190 9042
rect 40338 8990 40350 9042
rect 40402 8990 40414 9042
rect 42242 8990 42254 9042
rect 42306 8990 42318 9042
rect 46050 8990 46062 9042
rect 46114 8990 46126 9042
rect 37998 8978 38050 8990
rect 42814 8978 42866 8990
rect 8990 8930 9042 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 3602 8878 3614 8930
rect 3666 8878 3678 8930
rect 8990 8866 9042 8878
rect 9662 8930 9714 8942
rect 9662 8866 9714 8878
rect 10670 8930 10722 8942
rect 10670 8866 10722 8878
rect 16158 8930 16210 8942
rect 16158 8866 16210 8878
rect 16718 8930 16770 8942
rect 23998 8930 24050 8942
rect 28478 8930 28530 8942
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 20626 8878 20638 8930
rect 20690 8878 20702 8930
rect 22754 8878 22766 8930
rect 22818 8878 22830 8930
rect 25666 8878 25678 8930
rect 25730 8878 25742 8930
rect 16718 8866 16770 8878
rect 23998 8866 24050 8878
rect 28478 8866 28530 8878
rect 29262 8930 29314 8942
rect 29262 8866 29314 8878
rect 29710 8930 29762 8942
rect 32398 8930 32450 8942
rect 31490 8878 31502 8930
rect 31554 8878 31566 8930
rect 29710 8866 29762 8878
rect 32398 8866 32450 8878
rect 33518 8930 33570 8942
rect 39454 8930 39506 8942
rect 34962 8878 34974 8930
rect 35026 8878 35038 8930
rect 37090 8878 37102 8930
rect 37154 8878 37166 8930
rect 33518 8866 33570 8878
rect 39454 8866 39506 8878
rect 39790 8930 39842 8942
rect 42926 8930 42978 8942
rect 41346 8878 41358 8930
rect 41410 8878 41422 8930
rect 43250 8878 43262 8930
rect 43314 8878 43326 8930
rect 39790 8866 39842 8878
rect 42926 8866 42978 8878
rect 2942 8818 2994 8830
rect 2942 8754 2994 8766
rect 11230 8818 11282 8830
rect 11230 8754 11282 8766
rect 15262 8818 15314 8830
rect 15262 8754 15314 8766
rect 16830 8818 16882 8830
rect 32286 8818 32338 8830
rect 31826 8766 31838 8818
rect 31890 8766 31902 8818
rect 16830 8754 16882 8766
rect 32286 8754 32338 8766
rect 37774 8818 37826 8830
rect 37774 8754 37826 8766
rect 38446 8818 38498 8830
rect 38446 8754 38498 8766
rect 1344 8650 46592 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 46592 8650
rect 1344 8564 46592 8598
rect 41022 8482 41074 8494
rect 22306 8430 22318 8482
rect 22370 8430 22382 8482
rect 22642 8430 22654 8482
rect 22706 8479 22718 8482
rect 23314 8479 23326 8482
rect 22706 8433 23326 8479
rect 22706 8430 22718 8433
rect 23314 8430 23326 8433
rect 23378 8430 23390 8482
rect 38882 8430 38894 8482
rect 38946 8430 38958 8482
rect 41022 8418 41074 8430
rect 3502 8370 3554 8382
rect 3502 8306 3554 8318
rect 4846 8370 4898 8382
rect 23662 8370 23714 8382
rect 6402 8318 6414 8370
rect 6466 8318 6478 8370
rect 8530 8318 8542 8370
rect 8594 8318 8606 8370
rect 11106 8318 11118 8370
rect 11170 8318 11182 8370
rect 14802 8318 14814 8370
rect 14866 8318 14878 8370
rect 4846 8306 4898 8318
rect 23662 8306 23714 8318
rect 25118 8370 25170 8382
rect 25118 8306 25170 8318
rect 27358 8370 27410 8382
rect 34414 8370 34466 8382
rect 40910 8370 40962 8382
rect 44830 8370 44882 8382
rect 28130 8318 28142 8370
rect 28194 8318 28206 8370
rect 31602 8318 31614 8370
rect 31666 8318 31678 8370
rect 33730 8318 33742 8370
rect 33794 8318 33806 8370
rect 38658 8318 38670 8370
rect 38722 8318 38734 8370
rect 40114 8318 40126 8370
rect 40178 8318 40190 8370
rect 41346 8318 41358 8370
rect 41410 8318 41422 8370
rect 43474 8318 43486 8370
rect 43538 8318 43550 8370
rect 27358 8306 27410 8318
rect 34414 8306 34466 8318
rect 40910 8306 40962 8318
rect 44830 8306 44882 8318
rect 3054 8258 3106 8270
rect 3054 8194 3106 8206
rect 4062 8258 4114 8270
rect 4062 8194 4114 8206
rect 4622 8258 4674 8270
rect 9326 8258 9378 8270
rect 5618 8206 5630 8258
rect 5682 8206 5694 8258
rect 4622 8194 4674 8206
rect 9326 8194 9378 8206
rect 9438 8258 9490 8270
rect 20302 8258 20354 8270
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 11442 8206 11454 8258
rect 11506 8206 11518 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 9438 8194 9490 8206
rect 20302 8194 20354 8206
rect 20638 8258 20690 8270
rect 24110 8258 24162 8270
rect 21970 8206 21982 8258
rect 22034 8206 22046 8258
rect 22418 8206 22430 8258
rect 22482 8206 22494 8258
rect 20638 8194 20690 8206
rect 24110 8194 24162 8206
rect 24334 8258 24386 8270
rect 24334 8194 24386 8206
rect 25006 8258 25058 8270
rect 25006 8194 25058 8206
rect 25566 8258 25618 8270
rect 25566 8194 25618 8206
rect 26126 8258 26178 8270
rect 26126 8194 26178 8206
rect 26350 8258 26402 8270
rect 26350 8194 26402 8206
rect 27470 8258 27522 8270
rect 27470 8194 27522 8206
rect 27806 8258 27858 8270
rect 27806 8194 27858 8206
rect 29038 8258 29090 8270
rect 29038 8194 29090 8206
rect 29374 8258 29426 8270
rect 29374 8194 29426 8206
rect 29598 8258 29650 8270
rect 29598 8194 29650 8206
rect 30494 8258 30546 8270
rect 34526 8258 34578 8270
rect 36990 8258 37042 8270
rect 30930 8206 30942 8258
rect 30994 8206 31006 8258
rect 34066 8206 34078 8258
rect 34130 8206 34142 8258
rect 34738 8206 34750 8258
rect 34802 8206 34814 8258
rect 35298 8206 35310 8258
rect 35362 8206 35374 8258
rect 30494 8194 30546 8206
rect 34526 8194 34578 8206
rect 36990 8194 37042 8206
rect 37214 8258 37266 8270
rect 37214 8194 37266 8206
rect 37438 8258 37490 8270
rect 37998 8258 38050 8270
rect 45054 8258 45106 8270
rect 37650 8206 37662 8258
rect 37714 8206 37726 8258
rect 38546 8206 38558 8258
rect 38610 8206 38622 8258
rect 38770 8206 38782 8258
rect 38834 8206 38846 8258
rect 40002 8206 40014 8258
rect 40066 8206 40078 8258
rect 44258 8206 44270 8258
rect 44322 8206 44334 8258
rect 45378 8206 45390 8258
rect 45442 8206 45454 8258
rect 45938 8206 45950 8258
rect 46002 8206 46014 8258
rect 37438 8194 37490 8206
rect 37998 8194 38050 8206
rect 45054 8194 45106 8206
rect 10222 8146 10274 8158
rect 4274 8094 4286 8146
rect 4338 8094 4350 8146
rect 10222 8082 10274 8094
rect 10446 8146 10498 8158
rect 10446 8082 10498 8094
rect 10782 8146 10834 8158
rect 10782 8082 10834 8094
rect 12910 8146 12962 8158
rect 12910 8082 12962 8094
rect 14142 8146 14194 8158
rect 14142 8082 14194 8094
rect 21758 8146 21810 8158
rect 21758 8082 21810 8094
rect 25342 8146 25394 8158
rect 25342 8082 25394 8094
rect 25902 8146 25954 8158
rect 25902 8082 25954 8094
rect 28478 8146 28530 8158
rect 28478 8082 28530 8094
rect 29262 8146 29314 8158
rect 36094 8146 36146 8158
rect 35074 8094 35086 8146
rect 35138 8094 35150 8146
rect 29262 8082 29314 8094
rect 36094 8082 36146 8094
rect 2270 8034 2322 8046
rect 2270 7970 2322 7982
rect 2606 8034 2658 8046
rect 2606 7970 2658 7982
rect 2830 8034 2882 8046
rect 2830 7970 2882 7982
rect 2942 8034 2994 8046
rect 2942 7970 2994 7982
rect 3390 8034 3442 8046
rect 3390 7970 3442 7982
rect 3614 8034 3666 8046
rect 10334 8034 10386 8046
rect 20190 8034 20242 8046
rect 8866 7982 8878 8034
rect 8930 7982 8942 8034
rect 13794 7982 13806 8034
rect 13858 7982 13870 8034
rect 3614 7970 3666 7982
rect 10334 7970 10386 7982
rect 20190 7970 20242 7982
rect 20414 8034 20466 8046
rect 20414 7970 20466 7982
rect 20526 8034 20578 8046
rect 20526 7970 20578 7982
rect 21422 8034 21474 8046
rect 21422 7970 21474 7982
rect 22542 8034 22594 8046
rect 22542 7970 22594 7982
rect 23214 8034 23266 8046
rect 23214 7970 23266 7982
rect 24446 8034 24498 8046
rect 24446 7970 24498 7982
rect 24670 8034 24722 8046
rect 24670 7970 24722 7982
rect 26014 8034 26066 8046
rect 26014 7970 26066 7982
rect 27694 8034 27746 8046
rect 27694 7970 27746 7982
rect 28254 8034 28306 8046
rect 34302 8034 34354 8046
rect 30146 7982 30158 8034
rect 30210 7982 30222 8034
rect 28254 7970 28306 7982
rect 34302 7970 34354 7982
rect 36206 8034 36258 8046
rect 36206 7970 36258 7982
rect 37102 8034 37154 8046
rect 37102 7970 37154 7982
rect 45726 8034 45778 8046
rect 45726 7970 45778 7982
rect 1344 7866 46592 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 46592 7866
rect 1344 7780 46592 7814
rect 16606 7698 16658 7710
rect 16606 7634 16658 7646
rect 20638 7698 20690 7710
rect 20638 7634 20690 7646
rect 22990 7698 23042 7710
rect 22990 7634 23042 7646
rect 23662 7698 23714 7710
rect 23662 7634 23714 7646
rect 30830 7698 30882 7710
rect 30830 7634 30882 7646
rect 32062 7698 32114 7710
rect 32062 7634 32114 7646
rect 32174 7698 32226 7710
rect 32174 7634 32226 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 34078 7698 34130 7710
rect 34078 7634 34130 7646
rect 34526 7698 34578 7710
rect 34526 7634 34578 7646
rect 38558 7698 38610 7710
rect 38558 7634 38610 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 4958 7586 5010 7598
rect 4958 7522 5010 7534
rect 5182 7586 5234 7598
rect 16830 7586 16882 7598
rect 10322 7534 10334 7586
rect 10386 7534 10398 7586
rect 13906 7534 13918 7586
rect 13970 7534 13982 7586
rect 5182 7522 5234 7534
rect 16830 7522 16882 7534
rect 20302 7586 20354 7598
rect 20302 7522 20354 7534
rect 22206 7586 22258 7598
rect 22206 7522 22258 7534
rect 22878 7586 22930 7598
rect 22878 7522 22930 7534
rect 25230 7586 25282 7598
rect 26238 7586 26290 7598
rect 25554 7534 25566 7586
rect 25618 7534 25630 7586
rect 25230 7522 25282 7534
rect 26238 7522 26290 7534
rect 26350 7586 26402 7598
rect 32510 7586 32562 7598
rect 28018 7534 28030 7586
rect 28082 7534 28094 7586
rect 31490 7534 31502 7586
rect 31554 7534 31566 7586
rect 26350 7522 26402 7534
rect 32510 7522 32562 7534
rect 33630 7586 33682 7598
rect 33630 7522 33682 7534
rect 33966 7586 34018 7598
rect 39678 7586 39730 7598
rect 36978 7534 36990 7586
rect 37042 7534 37054 7586
rect 33966 7522 34018 7534
rect 39678 7522 39730 7534
rect 39902 7586 39954 7598
rect 39902 7522 39954 7534
rect 40238 7586 40290 7598
rect 44146 7534 44158 7586
rect 44210 7534 44222 7586
rect 40238 7522 40290 7534
rect 20526 7474 20578 7486
rect 4498 7422 4510 7474
rect 4562 7422 4574 7474
rect 5618 7422 5630 7474
rect 5682 7422 5694 7474
rect 9538 7422 9550 7474
rect 9602 7422 9614 7474
rect 13122 7422 13134 7474
rect 13186 7422 13198 7474
rect 17378 7422 17390 7474
rect 17442 7422 17454 7474
rect 20526 7410 20578 7422
rect 20750 7474 20802 7486
rect 22654 7474 22706 7486
rect 20962 7422 20974 7474
rect 21026 7422 21038 7474
rect 21858 7422 21870 7474
rect 21922 7422 21934 7474
rect 20750 7410 20802 7422
rect 22654 7410 22706 7422
rect 22766 7474 22818 7486
rect 24334 7474 24386 7486
rect 23202 7422 23214 7474
rect 23266 7422 23278 7474
rect 22766 7410 22818 7422
rect 24334 7410 24386 7422
rect 24558 7474 24610 7486
rect 24558 7410 24610 7422
rect 26126 7474 26178 7486
rect 32286 7474 32338 7486
rect 27346 7422 27358 7474
rect 27410 7422 27422 7474
rect 31266 7422 31278 7474
rect 31330 7422 31342 7474
rect 31826 7422 31838 7474
rect 31890 7422 31902 7474
rect 26126 7410 26178 7422
rect 32286 7410 32338 7422
rect 34414 7474 34466 7486
rect 38334 7474 38386 7486
rect 37650 7422 37662 7474
rect 37714 7422 37726 7474
rect 34414 7410 34466 7422
rect 38334 7410 38386 7422
rect 38446 7474 38498 7486
rect 38446 7410 38498 7422
rect 38670 7474 38722 7486
rect 38882 7422 38894 7474
rect 38946 7422 38958 7474
rect 44706 7422 44718 7474
rect 44770 7422 44782 7474
rect 38670 7410 38722 7422
rect 5070 7362 5122 7374
rect 8990 7362 9042 7374
rect 21646 7362 21698 7374
rect 1698 7310 1710 7362
rect 1762 7310 1774 7362
rect 3826 7310 3838 7362
rect 3890 7310 3902 7362
rect 6402 7310 6414 7362
rect 6466 7310 6478 7362
rect 8530 7310 8542 7362
rect 8594 7310 8606 7362
rect 12450 7310 12462 7362
rect 12514 7310 12526 7362
rect 16034 7310 16046 7362
rect 16098 7310 16110 7362
rect 16482 7310 16494 7362
rect 16546 7310 16558 7362
rect 18498 7310 18510 7362
rect 18562 7310 18574 7362
rect 5070 7298 5122 7310
rect 8990 7298 9042 7310
rect 21646 7298 21698 7310
rect 22094 7362 22146 7374
rect 22094 7298 22146 7310
rect 24222 7362 24274 7374
rect 39342 7362 39394 7374
rect 26786 7310 26798 7362
rect 26850 7310 26862 7362
rect 30146 7310 30158 7362
rect 30210 7310 30222 7362
rect 34850 7310 34862 7362
rect 34914 7310 34926 7362
rect 24222 7298 24274 7310
rect 39342 7298 39394 7310
rect 24670 7250 24722 7262
rect 24670 7186 24722 7198
rect 39230 7250 39282 7262
rect 39230 7186 39282 7198
rect 1344 7082 46592 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 46592 7082
rect 1344 6996 46592 7030
rect 3838 6914 3890 6926
rect 3838 6850 3890 6862
rect 12238 6914 12290 6926
rect 12238 6850 12290 6862
rect 12910 6914 12962 6926
rect 22654 6914 22706 6926
rect 21858 6862 21870 6914
rect 21922 6862 21934 6914
rect 12910 6850 12962 6862
rect 22654 6850 22706 6862
rect 23438 6914 23490 6926
rect 23438 6850 23490 6862
rect 43598 6914 43650 6926
rect 43598 6850 43650 6862
rect 43710 6914 43762 6926
rect 43710 6850 43762 6862
rect 43934 6914 43986 6926
rect 43934 6850 43986 6862
rect 44158 6914 44210 6926
rect 44158 6850 44210 6862
rect 45278 6914 45330 6926
rect 45278 6850 45330 6862
rect 45502 6914 45554 6926
rect 45502 6850 45554 6862
rect 3278 6802 3330 6814
rect 3278 6738 3330 6750
rect 4958 6802 5010 6814
rect 4958 6738 5010 6750
rect 5630 6802 5682 6814
rect 5630 6738 5682 6750
rect 5742 6802 5794 6814
rect 5742 6738 5794 6750
rect 6414 6802 6466 6814
rect 15598 6802 15650 6814
rect 19854 6802 19906 6814
rect 10994 6750 11006 6802
rect 11058 6750 11070 6802
rect 12562 6750 12574 6802
rect 12626 6750 12638 6802
rect 19170 6750 19182 6802
rect 19234 6750 19246 6802
rect 6414 6738 6466 6750
rect 15598 6738 15650 6750
rect 19854 6738 19906 6750
rect 23214 6802 23266 6814
rect 44942 6802 44994 6814
rect 24658 6750 24670 6802
rect 24722 6750 24734 6802
rect 26786 6750 26798 6802
rect 26850 6750 26862 6802
rect 29138 6750 29150 6802
rect 29202 6750 29214 6802
rect 23214 6738 23266 6750
rect 44942 6738 44994 6750
rect 45054 6802 45106 6814
rect 45054 6738 45106 6750
rect 3614 6690 3666 6702
rect 4398 6690 4450 6702
rect 4162 6638 4174 6690
rect 4226 6638 4238 6690
rect 3614 6626 3666 6638
rect 4398 6626 4450 6638
rect 5070 6690 5122 6702
rect 6190 6690 6242 6702
rect 5954 6638 5966 6690
rect 6018 6638 6030 6690
rect 5070 6626 5122 6638
rect 6190 6626 6242 6638
rect 6862 6690 6914 6702
rect 6862 6626 6914 6638
rect 7310 6690 7362 6702
rect 7310 6626 7362 6638
rect 7870 6690 7922 6702
rect 15374 6690 15426 6702
rect 19630 6690 19682 6702
rect 28366 6690 28418 6702
rect 40462 6690 40514 6702
rect 8194 6638 8206 6690
rect 8258 6638 8270 6690
rect 16370 6638 16382 6690
rect 16434 6638 16446 6690
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 20178 6638 20190 6690
rect 20242 6638 20254 6690
rect 21858 6638 21870 6690
rect 21922 6638 21934 6690
rect 23986 6638 23998 6690
rect 24050 6638 24062 6690
rect 28130 6638 28142 6690
rect 28194 6638 28206 6690
rect 31938 6638 31950 6690
rect 32002 6638 32014 6690
rect 32722 6638 32734 6690
rect 32786 6638 32798 6690
rect 36194 6638 36206 6690
rect 36258 6638 36270 6690
rect 39442 6638 39454 6690
rect 39506 6638 39518 6690
rect 7870 6626 7922 6638
rect 15374 6626 15426 6638
rect 19630 6626 19682 6638
rect 28366 6626 28418 6638
rect 40462 6626 40514 6638
rect 40686 6690 40738 6702
rect 45614 6690 45666 6702
rect 40898 6638 40910 6690
rect 40962 6638 40974 6690
rect 41906 6638 41918 6690
rect 41970 6638 41982 6690
rect 42802 6638 42814 6690
rect 42866 6638 42878 6690
rect 40686 6626 40738 6638
rect 45614 6626 45666 6638
rect 6638 6578 6690 6590
rect 12014 6578 12066 6590
rect 8866 6526 8878 6578
rect 8930 6526 8942 6578
rect 6638 6514 6690 6526
rect 12014 6514 12066 6526
rect 12686 6578 12738 6590
rect 12686 6514 12738 6526
rect 14254 6578 14306 6590
rect 14254 6514 14306 6526
rect 15710 6578 15762 6590
rect 15710 6514 15762 6526
rect 21310 6578 21362 6590
rect 22878 6578 22930 6590
rect 21522 6526 21534 6578
rect 21586 6526 21598 6578
rect 21310 6514 21362 6526
rect 22878 6514 22930 6526
rect 28590 6578 28642 6590
rect 35646 6578 35698 6590
rect 31266 6526 31278 6578
rect 31330 6526 31342 6578
rect 28590 6514 28642 6526
rect 35646 6514 35698 6526
rect 36430 6578 36482 6590
rect 40014 6578 40066 6590
rect 37762 6526 37774 6578
rect 37826 6526 37838 6578
rect 36430 6514 36482 6526
rect 40014 6514 40066 6526
rect 40238 6578 40290 6590
rect 42130 6526 42142 6578
rect 42194 6526 42206 6578
rect 42914 6526 42926 6578
rect 42978 6526 42990 6578
rect 40238 6514 40290 6526
rect 4846 6466 4898 6478
rect 4846 6402 4898 6414
rect 7198 6466 7250 6478
rect 7198 6402 7250 6414
rect 7422 6466 7474 6478
rect 7422 6402 7474 6414
rect 11566 6466 11618 6478
rect 11566 6402 11618 6414
rect 12126 6466 12178 6478
rect 12126 6402 12178 6414
rect 13582 6466 13634 6478
rect 14478 6466 14530 6478
rect 13906 6414 13918 6466
rect 13970 6414 13982 6466
rect 13582 6402 13634 6414
rect 14478 6402 14530 6414
rect 14590 6466 14642 6478
rect 14590 6402 14642 6414
rect 14702 6466 14754 6478
rect 14702 6402 14754 6414
rect 14814 6466 14866 6478
rect 14814 6402 14866 6414
rect 15486 6466 15538 6478
rect 15486 6402 15538 6414
rect 15822 6466 15874 6478
rect 15822 6402 15874 6414
rect 19742 6466 19794 6478
rect 19742 6402 19794 6414
rect 19966 6466 20018 6478
rect 19966 6402 20018 6414
rect 20750 6466 20802 6478
rect 23550 6466 23602 6478
rect 21746 6414 21758 6466
rect 21810 6414 21822 6466
rect 20750 6402 20802 6414
rect 23550 6402 23602 6414
rect 33742 6466 33794 6478
rect 33742 6402 33794 6414
rect 35758 6466 35810 6478
rect 35758 6402 35810 6414
rect 40798 6466 40850 6478
rect 40798 6402 40850 6414
rect 44046 6466 44098 6478
rect 44046 6402 44098 6414
rect 46062 6466 46114 6478
rect 46062 6402 46114 6414
rect 1344 6298 46592 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 46592 6298
rect 1344 6212 46592 6246
rect 6190 6130 6242 6142
rect 6190 6066 6242 6078
rect 8542 6130 8594 6142
rect 8542 6066 8594 6078
rect 15262 6130 15314 6142
rect 15262 6066 15314 6078
rect 15374 6130 15426 6142
rect 15374 6066 15426 6078
rect 15598 6130 15650 6142
rect 15598 6066 15650 6078
rect 16382 6130 16434 6142
rect 16382 6066 16434 6078
rect 17726 6130 17778 6142
rect 18622 6130 18674 6142
rect 33294 6130 33346 6142
rect 18050 6078 18062 6130
rect 18114 6078 18126 6130
rect 26226 6078 26238 6130
rect 26290 6078 26302 6130
rect 17726 6066 17778 6078
rect 18622 6066 18674 6078
rect 33294 6066 33346 6078
rect 33518 6130 33570 6142
rect 33518 6066 33570 6078
rect 40238 6130 40290 6142
rect 40238 6066 40290 6078
rect 41022 6130 41074 6142
rect 41022 6066 41074 6078
rect 41134 6130 41186 6142
rect 41134 6066 41186 6078
rect 41246 6130 41298 6142
rect 41246 6066 41298 6078
rect 9102 6018 9154 6030
rect 2482 5966 2494 6018
rect 2546 5966 2558 6018
rect 9102 5954 9154 5966
rect 15822 6018 15874 6030
rect 33742 6018 33794 6030
rect 21634 5966 21646 6018
rect 21698 5966 21710 6018
rect 25554 5966 25566 6018
rect 25618 5966 25630 6018
rect 27346 5966 27358 6018
rect 27410 5966 27422 6018
rect 15822 5954 15874 5966
rect 33742 5954 33794 5966
rect 40350 6018 40402 6030
rect 40350 5954 40402 5966
rect 42254 6018 42306 6030
rect 42254 5954 42306 5966
rect 42366 6018 42418 6030
rect 45378 5966 45390 6018
rect 45442 5966 45454 6018
rect 42366 5954 42418 5966
rect 4958 5906 5010 5918
rect 1810 5854 1822 5906
rect 1874 5854 1886 5906
rect 4958 5842 5010 5854
rect 5182 5906 5234 5918
rect 7086 5906 7138 5918
rect 5954 5854 5966 5906
rect 6018 5854 6030 5906
rect 5182 5842 5234 5854
rect 7086 5842 7138 5854
rect 7198 5906 7250 5918
rect 7198 5842 7250 5854
rect 7310 5906 7362 5918
rect 7982 5906 8034 5918
rect 7522 5854 7534 5906
rect 7586 5854 7598 5906
rect 7310 5842 7362 5854
rect 7982 5842 8034 5854
rect 8206 5906 8258 5918
rect 16606 5906 16658 5918
rect 10098 5854 10110 5906
rect 10162 5854 10174 5906
rect 16146 5854 16158 5906
rect 16210 5854 16222 5906
rect 8206 5842 8258 5854
rect 16606 5842 16658 5854
rect 16718 5906 16770 5918
rect 18846 5906 18898 5918
rect 18386 5854 18398 5906
rect 18450 5854 18462 5906
rect 16718 5842 16770 5854
rect 18846 5842 18898 5854
rect 18958 5906 19010 5918
rect 25230 5906 25282 5918
rect 23650 5854 23662 5906
rect 23714 5854 23726 5906
rect 18958 5842 19010 5854
rect 25230 5842 25282 5854
rect 26574 5906 26626 5918
rect 33182 5906 33234 5918
rect 41470 5906 41522 5918
rect 31154 5854 31166 5906
rect 31218 5854 31230 5906
rect 39554 5854 39566 5906
rect 39618 5854 39630 5906
rect 40002 5854 40014 5906
rect 40066 5854 40078 5906
rect 26574 5842 26626 5854
rect 33182 5842 33234 5854
rect 41470 5842 41522 5854
rect 41694 5906 41746 5918
rect 41694 5842 41746 5854
rect 42142 5906 42194 5918
rect 46162 5854 46174 5906
rect 46226 5854 46238 5906
rect 42142 5842 42194 5854
rect 16494 5794 16546 5806
rect 4610 5742 4622 5794
rect 4674 5742 4686 5794
rect 13122 5742 13134 5794
rect 13186 5742 13198 5794
rect 15362 5742 15374 5794
rect 15426 5742 15438 5794
rect 16494 5730 16546 5742
rect 18734 5794 18786 5806
rect 18734 5730 18786 5742
rect 33406 5794 33458 5806
rect 34626 5742 34638 5794
rect 34690 5742 34702 5794
rect 42802 5742 42814 5794
rect 42866 5742 42878 5794
rect 43250 5742 43262 5794
rect 43314 5742 43326 5794
rect 33406 5730 33458 5742
rect 5506 5630 5518 5682
rect 5570 5630 5582 5682
rect 1344 5514 46592 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 46592 5514
rect 1344 5428 46592 5462
rect 9662 5346 9714 5358
rect 9662 5282 9714 5294
rect 25678 5346 25730 5358
rect 25678 5282 25730 5294
rect 26350 5346 26402 5358
rect 26350 5282 26402 5294
rect 26798 5346 26850 5358
rect 29486 5346 29538 5358
rect 29138 5294 29150 5346
rect 29202 5294 29214 5346
rect 26798 5282 26850 5294
rect 29486 5282 29538 5294
rect 30046 5346 30098 5358
rect 30046 5282 30098 5294
rect 30382 5346 30434 5358
rect 30382 5282 30434 5294
rect 40798 5346 40850 5358
rect 45378 5294 45390 5346
rect 45442 5294 45454 5346
rect 40798 5282 40850 5294
rect 8206 5234 8258 5246
rect 8206 5170 8258 5182
rect 8542 5234 8594 5246
rect 8542 5170 8594 5182
rect 9550 5234 9602 5246
rect 24558 5234 24610 5246
rect 10770 5182 10782 5234
rect 10834 5182 10846 5234
rect 12898 5182 12910 5234
rect 12962 5182 12974 5234
rect 16930 5182 16942 5234
rect 16994 5182 17006 5234
rect 19058 5182 19070 5234
rect 19122 5182 19134 5234
rect 22082 5182 22094 5234
rect 22146 5182 22158 5234
rect 24210 5182 24222 5234
rect 24274 5182 24286 5234
rect 9550 5170 9602 5182
rect 24558 5170 24610 5182
rect 24782 5234 24834 5246
rect 26462 5234 26514 5246
rect 26002 5182 26014 5234
rect 26066 5182 26078 5234
rect 24782 5170 24834 5182
rect 26462 5170 26514 5182
rect 27470 5234 27522 5246
rect 34526 5234 34578 5246
rect 36318 5234 36370 5246
rect 41022 5234 41074 5246
rect 44830 5234 44882 5246
rect 33842 5182 33854 5234
rect 33906 5182 33918 5234
rect 35410 5182 35422 5234
rect 35474 5182 35486 5234
rect 37762 5182 37774 5234
rect 37826 5182 37838 5234
rect 39890 5182 39902 5234
rect 39954 5182 39966 5234
rect 41346 5182 41358 5234
rect 41410 5182 41422 5234
rect 43474 5182 43486 5234
rect 43538 5182 43550 5234
rect 27470 5170 27522 5182
rect 34526 5170 34578 5182
rect 36318 5170 36370 5182
rect 41022 5170 41074 5182
rect 44830 5170 44882 5182
rect 4846 5122 4898 5134
rect 4846 5058 4898 5070
rect 5182 5122 5234 5134
rect 5182 5058 5234 5070
rect 6078 5122 6130 5134
rect 27806 5122 27858 5134
rect 6290 5070 6302 5122
rect 6354 5070 6366 5122
rect 10098 5070 10110 5122
rect 10162 5070 10174 5122
rect 15922 5070 15934 5122
rect 15986 5070 15998 5122
rect 19842 5070 19854 5122
rect 19906 5070 19918 5122
rect 20626 5070 20638 5122
rect 20690 5070 20702 5122
rect 21410 5070 21422 5122
rect 21474 5070 21486 5122
rect 25106 5070 25118 5122
rect 25170 5070 25182 5122
rect 27570 5070 27582 5122
rect 27634 5070 27646 5122
rect 6078 5058 6130 5070
rect 27806 5058 27858 5070
rect 29710 5122 29762 5134
rect 34302 5122 34354 5134
rect 30370 5070 30382 5122
rect 30434 5070 30446 5122
rect 30930 5070 30942 5122
rect 30994 5070 31006 5122
rect 29710 5058 29762 5070
rect 34302 5058 34354 5070
rect 34414 5122 34466 5134
rect 34414 5058 34466 5070
rect 34750 5122 34802 5134
rect 45054 5122 45106 5134
rect 35186 5070 35198 5122
rect 35250 5070 35262 5122
rect 36978 5070 36990 5122
rect 37042 5070 37054 5122
rect 44258 5070 44270 5122
rect 44322 5070 44334 5122
rect 45938 5070 45950 5122
rect 46002 5070 46014 5122
rect 34750 5058 34802 5070
rect 45054 5058 45106 5070
rect 4958 5010 5010 5022
rect 4958 4946 5010 4958
rect 6974 5010 7026 5022
rect 6974 4946 7026 4958
rect 9438 5010 9490 5022
rect 25902 5010 25954 5022
rect 20402 4958 20414 5010
rect 20466 4958 20478 5010
rect 9438 4946 9490 4958
rect 25902 4946 25954 4958
rect 27022 5010 27074 5022
rect 35646 5010 35698 5022
rect 31714 4958 31726 5010
rect 31778 4958 31790 5010
rect 27022 4946 27074 4958
rect 35646 4946 35698 4958
rect 35870 5010 35922 5022
rect 35870 4946 35922 4958
rect 8990 4898 9042 4910
rect 8990 4834 9042 4846
rect 15374 4898 15426 4910
rect 15374 4834 15426 4846
rect 26910 4898 26962 4910
rect 26910 4834 26962 4846
rect 34638 4898 34690 4910
rect 34638 4834 34690 4846
rect 35422 4898 35474 4910
rect 35422 4834 35474 4846
rect 36430 4898 36482 4910
rect 45726 4898 45778 4910
rect 40450 4846 40462 4898
rect 40514 4846 40526 4898
rect 36430 4834 36482 4846
rect 45726 4834 45778 4846
rect 1344 4730 46592 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 46592 4730
rect 1344 4644 46592 4678
rect 8654 4562 8706 4574
rect 8654 4498 8706 4510
rect 17726 4562 17778 4574
rect 17726 4498 17778 4510
rect 31838 4562 31890 4574
rect 31838 4498 31890 4510
rect 32286 4562 32338 4574
rect 32286 4498 32338 4510
rect 41022 4562 41074 4574
rect 41022 4498 41074 4510
rect 7422 4450 7474 4462
rect 7422 4386 7474 4398
rect 9662 4450 9714 4462
rect 13582 4450 13634 4462
rect 24446 4450 24498 4462
rect 31950 4450 32002 4462
rect 10770 4398 10782 4450
rect 10834 4398 10846 4450
rect 14690 4398 14702 4450
rect 14754 4398 14766 4450
rect 21970 4398 21982 4450
rect 22034 4398 22046 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 9662 4386 9714 4398
rect 13582 4386 13634 4398
rect 24446 4386 24498 4398
rect 31950 4386 32002 4398
rect 32398 4450 32450 4462
rect 40126 4450 40178 4462
rect 33842 4398 33854 4450
rect 33906 4398 33918 4450
rect 37090 4398 37102 4450
rect 37154 4398 37166 4450
rect 32398 4386 32450 4398
rect 40126 4386 40178 4398
rect 42478 4450 42530 4462
rect 45378 4398 45390 4450
rect 45442 4398 45454 4450
rect 42478 4386 42530 4398
rect 31614 4338 31666 4350
rect 40014 4338 40066 4350
rect 40798 4338 40850 4350
rect 7074 4286 7086 4338
rect 7138 4286 7150 4338
rect 7746 4286 7758 4338
rect 7810 4286 7822 4338
rect 8418 4286 8430 4338
rect 8482 4286 8494 4338
rect 10098 4286 10110 4338
rect 10162 4286 10174 4338
rect 13234 4286 13246 4338
rect 13298 4286 13310 4338
rect 14018 4286 14030 4338
rect 14082 4286 14094 4338
rect 18050 4286 18062 4338
rect 18114 4286 18126 4338
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 28578 4286 28590 4338
rect 28642 4286 28654 4338
rect 33058 4286 33070 4338
rect 33122 4286 33134 4338
rect 36306 4286 36318 4338
rect 36370 4286 36382 4338
rect 40338 4286 40350 4338
rect 40402 4286 40414 4338
rect 31614 4274 31666 4286
rect 40014 4274 40066 4286
rect 40798 4274 40850 4286
rect 41134 4338 41186 4350
rect 42018 4286 42030 4338
rect 42082 4286 42094 4338
rect 46162 4286 46174 4338
rect 46226 4286 46238 4338
rect 41134 4274 41186 4286
rect 7534 4226 7586 4238
rect 42814 4226 42866 4238
rect 4162 4174 4174 4226
rect 4226 4174 4238 4226
rect 6290 4174 6302 4226
rect 6354 4174 6366 4226
rect 12898 4174 12910 4226
rect 12962 4174 12974 4226
rect 13346 4174 13358 4226
rect 13410 4174 13422 4226
rect 16818 4174 16830 4226
rect 16882 4174 16894 4226
rect 18722 4174 18734 4226
rect 18786 4174 18798 4226
rect 20850 4174 20862 4226
rect 20914 4174 20926 4226
rect 24098 4174 24110 4226
rect 24162 4174 24174 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 29250 4174 29262 4226
rect 29314 4174 29326 4226
rect 31378 4174 31390 4226
rect 31442 4174 31454 4226
rect 35970 4174 35982 4226
rect 36034 4174 36046 4226
rect 39218 4174 39230 4226
rect 39282 4174 39294 4226
rect 41570 4174 41582 4226
rect 41634 4174 41646 4226
rect 43250 4174 43262 4226
rect 43314 4174 43326 4226
rect 7534 4162 7586 4174
rect 42814 4162 42866 4174
rect 42926 4114 42978 4126
rect 39554 4062 39566 4114
rect 39618 4062 39630 4114
rect 42926 4050 42978 4062
rect 1344 3946 46592 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 46592 3946
rect 1344 3860 46592 3894
rect 8766 3778 8818 3790
rect 8766 3714 8818 3726
rect 23662 3778 23714 3790
rect 23662 3714 23714 3726
rect 27470 3778 27522 3790
rect 27470 3714 27522 3726
rect 38894 3778 38946 3790
rect 38894 3714 38946 3726
rect 39230 3778 39282 3790
rect 39230 3714 39282 3726
rect 44606 3778 44658 3790
rect 44606 3714 44658 3726
rect 18622 3666 18674 3678
rect 23774 3666 23826 3678
rect 12562 3614 12574 3666
rect 12626 3614 12638 3666
rect 13906 3614 13918 3666
rect 13970 3614 13982 3666
rect 16034 3614 16046 3666
rect 16098 3614 16110 3666
rect 21858 3614 21870 3666
rect 21922 3614 21934 3666
rect 18622 3602 18674 3614
rect 23774 3602 23826 3614
rect 27582 3666 27634 3678
rect 36990 3666 37042 3678
rect 29474 3614 29486 3666
rect 29538 3614 29550 3666
rect 31602 3614 31614 3666
rect 31666 3614 31678 3666
rect 40114 3614 40126 3666
rect 40178 3614 40190 3666
rect 42242 3614 42254 3666
rect 42306 3614 42318 3666
rect 27582 3602 27634 3614
rect 36990 3602 37042 3614
rect 17278 3554 17330 3566
rect 26686 3554 26738 3566
rect 9762 3502 9774 3554
rect 9826 3502 9838 3554
rect 13122 3502 13134 3554
rect 13186 3502 13198 3554
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 20962 3502 20974 3554
rect 21026 3502 21038 3554
rect 23986 3502 23998 3554
rect 24050 3502 24062 3554
rect 28690 3502 28702 3554
rect 28754 3502 28766 3554
rect 32162 3502 32174 3554
rect 32226 3502 32238 3554
rect 35186 3502 35198 3554
rect 35250 3502 35262 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 43026 3502 43038 3554
rect 43090 3502 43102 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 17278 3490 17330 3502
rect 26686 3490 26738 3502
rect 8542 3442 8594 3454
rect 8542 3378 8594 3390
rect 8654 3442 8706 3454
rect 35422 3442 35474 3454
rect 10434 3390 10446 3442
rect 10498 3390 10510 3442
rect 16930 3390 16942 3442
rect 16994 3390 17006 3442
rect 26338 3390 26350 3442
rect 26402 3390 26414 3442
rect 33730 3390 33742 3442
rect 33794 3390 33806 3442
rect 8654 3378 8706 3390
rect 35422 3378 35474 3390
rect 39118 3442 39170 3454
rect 39118 3378 39170 3390
rect 2942 3330 2994 3342
rect 2942 3266 2994 3278
rect 4510 3330 4562 3342
rect 4510 3266 4562 3278
rect 6078 3330 6130 3342
rect 6078 3266 6130 3278
rect 7534 3330 7586 3342
rect 7534 3266 7586 3278
rect 8094 3330 8146 3342
rect 8094 3266 8146 3278
rect 24894 3330 24946 3342
rect 24894 3266 24946 3278
rect 25342 3330 25394 3342
rect 25342 3266 25394 3278
rect 26014 3330 26066 3342
rect 26014 3266 26066 3278
rect 27022 3330 27074 3342
rect 27022 3266 27074 3278
rect 1344 3162 46592 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 46592 3162
rect 1344 3076 46592 3110
<< via1 >>
rect 13582 44830 13634 44882
rect 14478 44830 14530 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 31278 44494 31330 44546
rect 10110 44382 10162 44434
rect 14478 44382 14530 44434
rect 14590 44382 14642 44434
rect 15598 44382 15650 44434
rect 15822 44382 15874 44434
rect 20078 44382 20130 44434
rect 23102 44382 23154 44434
rect 23550 44382 23602 44434
rect 27806 44382 27858 44434
rect 29150 44382 29202 44434
rect 32510 44382 32562 44434
rect 39230 44382 39282 44434
rect 43038 44382 43090 44434
rect 13582 44270 13634 44322
rect 14142 44270 14194 44322
rect 17502 44270 17554 44322
rect 18174 44270 18226 44322
rect 18734 44270 18786 44322
rect 21758 44270 21810 44322
rect 22766 44270 22818 44322
rect 25006 44270 25058 44322
rect 30046 44270 30098 44322
rect 30606 44270 30658 44322
rect 34526 44270 34578 44322
rect 34862 44270 34914 44322
rect 36430 44270 36482 44322
rect 40126 44270 40178 44322
rect 45166 44270 45218 44322
rect 9774 44158 9826 44210
rect 13694 44158 13746 44210
rect 16158 44158 16210 44210
rect 20190 44158 20242 44210
rect 20750 44158 20802 44210
rect 21534 44158 21586 44210
rect 21870 44158 21922 44210
rect 22542 44158 22594 44210
rect 25678 44158 25730 44210
rect 29710 44158 29762 44210
rect 30942 44158 30994 44210
rect 32174 44158 32226 44210
rect 33406 44158 33458 44210
rect 33518 44158 33570 44210
rect 33854 44158 33906 44210
rect 35422 44158 35474 44210
rect 37102 44158 37154 44210
rect 40910 44158 40962 44210
rect 43598 44158 43650 44210
rect 44270 44158 44322 44210
rect 44942 44158 44994 44210
rect 9550 44046 9602 44098
rect 9998 44046 10050 44098
rect 13806 44046 13858 44098
rect 15150 44046 15202 44098
rect 15934 44046 15986 44098
rect 17950 44046 18002 44098
rect 19294 44046 19346 44098
rect 19854 44046 19906 44098
rect 20862 44046 20914 44098
rect 21086 44046 21138 44098
rect 21982 44046 22034 44098
rect 22094 44046 22146 44098
rect 22990 44046 23042 44098
rect 23102 44046 23154 44098
rect 23662 44046 23714 44098
rect 28702 44046 28754 44098
rect 29486 44046 29538 44098
rect 29598 44046 29650 44098
rect 31166 44046 31218 44098
rect 32398 44046 32450 44098
rect 33182 44046 33234 44098
rect 33966 44046 34018 44098
rect 34190 44046 34242 44098
rect 43710 44046 43762 44098
rect 44382 44046 44434 44098
rect 44494 44046 44546 44098
rect 45614 44046 45666 44098
rect 45950 44046 46002 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 8878 43710 8930 43762
rect 29486 43710 29538 43762
rect 19070 43598 19122 43650
rect 23886 43598 23938 43650
rect 29150 43598 29202 43650
rect 30158 43598 30210 43650
rect 31054 43598 31106 43650
rect 32622 43598 32674 43650
rect 39902 43598 39954 43650
rect 5966 43486 6018 43538
rect 10110 43486 10162 43538
rect 10782 43486 10834 43538
rect 14030 43486 14082 43538
rect 17614 43486 17666 43538
rect 18398 43486 18450 43538
rect 24558 43486 24610 43538
rect 25230 43486 25282 43538
rect 25678 43486 25730 43538
rect 29822 43486 29874 43538
rect 30718 43486 30770 43538
rect 31726 43486 31778 43538
rect 31838 43486 31890 43538
rect 35982 43486 36034 43538
rect 36430 43486 36482 43538
rect 39454 43486 39506 43538
rect 40014 43486 40066 43538
rect 41022 43486 41074 43538
rect 41134 43486 41186 43538
rect 41246 43486 41298 43538
rect 42142 43486 42194 43538
rect 42366 43486 42418 43538
rect 43262 43486 43314 43538
rect 6638 43374 6690 43426
rect 11454 43374 11506 43426
rect 13582 43374 13634 43426
rect 14702 43374 14754 43426
rect 16830 43374 16882 43426
rect 17838 43374 17890 43426
rect 21198 43374 21250 43426
rect 21646 43374 21698 43426
rect 26462 43374 26514 43426
rect 28590 43374 28642 43426
rect 30494 43374 30546 43426
rect 31390 43374 31442 43426
rect 33070 43374 33122 43426
rect 35198 43374 35250 43426
rect 37102 43374 37154 43426
rect 39230 43374 39282 43426
rect 39678 43374 39730 43426
rect 44046 43374 44098 43426
rect 46174 43374 46226 43426
rect 9550 43262 9602 43314
rect 9886 43262 9938 43314
rect 17950 43262 18002 43314
rect 25342 43262 25394 43314
rect 31502 43262 31554 43314
rect 41694 43262 41746 43314
rect 42030 43262 42082 43314
rect 42478 43262 42530 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 9998 42926 10050 42978
rect 10670 42926 10722 42978
rect 11006 42926 11058 42978
rect 11342 42926 11394 42978
rect 11678 42926 11730 42978
rect 13470 42926 13522 42978
rect 14814 42926 14866 42978
rect 20078 42926 20130 42978
rect 31054 42926 31106 42978
rect 32510 42926 32562 42978
rect 32846 42926 32898 42978
rect 35310 42926 35362 42978
rect 35646 42926 35698 42978
rect 38446 42926 38498 42978
rect 39118 42926 39170 42978
rect 9214 42814 9266 42866
rect 18622 42814 18674 42866
rect 19294 42814 19346 42866
rect 21758 42814 21810 42866
rect 24782 42814 24834 42866
rect 26462 42814 26514 42866
rect 29262 42814 29314 42866
rect 30494 42814 30546 42866
rect 33518 42814 33570 42866
rect 39454 42814 39506 42866
rect 41582 42814 41634 42866
rect 42814 42814 42866 42866
rect 9662 42702 9714 42754
rect 9886 42702 9938 42754
rect 10558 42702 10610 42754
rect 10894 42702 10946 42754
rect 11454 42702 11506 42754
rect 11902 42702 11954 42754
rect 13918 42702 13970 42754
rect 14142 42702 14194 42754
rect 14926 42702 14978 42754
rect 15150 42702 15202 42754
rect 15374 42702 15426 42754
rect 15822 42702 15874 42754
rect 19182 42702 19234 42754
rect 20414 42702 20466 42754
rect 20638 42702 20690 42754
rect 21870 42702 21922 42754
rect 22878 42702 22930 42754
rect 23550 42702 23602 42754
rect 24334 42702 24386 42754
rect 26350 42702 26402 42754
rect 26686 42702 26738 42754
rect 29486 42702 29538 42754
rect 30046 42702 30098 42754
rect 30718 42702 30770 42754
rect 32398 42702 32450 42754
rect 32734 42702 32786 42754
rect 35646 42702 35698 42754
rect 36094 42702 36146 42754
rect 37550 42702 37602 42754
rect 37774 42702 37826 42754
rect 37998 42702 38050 42754
rect 38558 42702 38610 42754
rect 38782 42702 38834 42754
rect 39006 42702 39058 42754
rect 42366 42702 42418 42754
rect 43038 42702 43090 42754
rect 45278 42702 45330 42754
rect 9550 42590 9602 42642
rect 12910 42590 12962 42642
rect 14030 42590 14082 42642
rect 16494 42590 16546 42642
rect 26126 42590 26178 42642
rect 29598 42590 29650 42642
rect 33182 42590 33234 42642
rect 33406 42590 33458 42642
rect 34414 42590 34466 42642
rect 34638 42590 34690 42642
rect 43710 42590 43762 42642
rect 44270 42590 44322 42642
rect 44830 42590 44882 42642
rect 45390 42590 45442 42642
rect 45502 42590 45554 42642
rect 46062 42590 46114 42642
rect 12798 42478 12850 42530
rect 26574 42478 26626 42530
rect 27358 42478 27410 42530
rect 27806 42478 27858 42530
rect 28142 42478 28194 42530
rect 28702 42478 28754 42530
rect 30270 42478 30322 42530
rect 31502 42478 31554 42530
rect 31950 42478 32002 42530
rect 34974 42478 35026 42530
rect 36318 42478 36370 42530
rect 37214 42478 37266 42530
rect 37886 42478 37938 42530
rect 43934 42478 43986 42530
rect 44158 42478 44210 42530
rect 45950 42478 46002 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 15822 42142 15874 42194
rect 16382 42142 16434 42194
rect 18846 42142 18898 42194
rect 31054 42142 31106 42194
rect 36654 42142 36706 42194
rect 17502 42030 17554 42082
rect 32174 42030 32226 42082
rect 5966 41918 6018 41970
rect 6638 41918 6690 41970
rect 13694 41918 13746 41970
rect 15486 41918 15538 41970
rect 15710 41918 15762 41970
rect 15934 41918 15986 41970
rect 16494 41918 16546 41970
rect 18062 41918 18114 41970
rect 18398 41918 18450 41970
rect 19406 41918 19458 41970
rect 30158 41918 30210 41970
rect 30942 41918 30994 41970
rect 31166 41918 31218 41970
rect 31838 41918 31890 41970
rect 35982 41918 36034 41970
rect 36318 41918 36370 41970
rect 37102 41918 37154 41970
rect 37438 41918 37490 41970
rect 44718 41918 44770 41970
rect 8766 41806 8818 41858
rect 10110 41806 10162 41858
rect 18174 41806 18226 41858
rect 21982 41806 22034 41858
rect 28030 41806 28082 41858
rect 33070 41806 33122 41858
rect 35198 41806 35250 41858
rect 36990 41806 37042 41858
rect 38222 41806 38274 41858
rect 40350 41806 40402 41858
rect 42702 41806 42754 41858
rect 16382 41694 16434 41746
rect 16718 41694 16770 41746
rect 31390 41694 31442 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 9326 41358 9378 41410
rect 9662 41358 9714 41410
rect 30830 41358 30882 41410
rect 33182 41358 33234 41410
rect 33294 41358 33346 41410
rect 33630 41358 33682 41410
rect 35310 41358 35362 41410
rect 35646 41358 35698 41410
rect 36094 41358 36146 41410
rect 45166 41358 45218 41410
rect 12910 41246 12962 41298
rect 14926 41246 14978 41298
rect 15262 41246 15314 41298
rect 16270 41246 16322 41298
rect 21310 41246 21362 41298
rect 24670 41246 24722 41298
rect 28142 41246 28194 41298
rect 30270 41246 30322 41298
rect 32398 41246 32450 41298
rect 35086 41246 35138 41298
rect 37214 41246 37266 41298
rect 43934 41246 43986 41298
rect 45838 41246 45890 41298
rect 9102 41134 9154 41186
rect 10110 41134 10162 41186
rect 14702 41134 14754 41186
rect 15598 41134 15650 41186
rect 17278 41134 17330 41186
rect 18062 41134 18114 41186
rect 18398 41134 18450 41186
rect 20414 41134 20466 41186
rect 24222 41134 24274 41186
rect 25342 41134 25394 41186
rect 30046 41134 30098 41186
rect 30494 41134 30546 41186
rect 33518 41134 33570 41186
rect 36430 41134 36482 41186
rect 41918 41134 41970 41186
rect 42590 41134 42642 41186
rect 43486 41134 43538 41186
rect 43710 41134 43762 41186
rect 44830 41134 44882 41186
rect 44942 41134 44994 41186
rect 45278 41134 45330 41186
rect 10782 41022 10834 41074
rect 14030 41022 14082 41074
rect 15822 41022 15874 41074
rect 16158 41022 16210 41074
rect 20638 41022 20690 41074
rect 23438 41022 23490 41074
rect 26014 41022 26066 41074
rect 28590 41022 28642 41074
rect 31166 41022 31218 41074
rect 31950 41022 32002 41074
rect 44046 41022 44098 41074
rect 45726 41022 45778 41074
rect 13694 40910 13746 40962
rect 20862 40910 20914 40962
rect 24558 40910 24610 40962
rect 28478 40910 28530 40962
rect 29374 40910 29426 40962
rect 29486 40910 29538 40962
rect 29598 40910 29650 40962
rect 31278 40910 31330 40962
rect 31390 40910 31442 40962
rect 31838 40910 31890 40962
rect 32286 40910 32338 40962
rect 32846 40910 32898 40962
rect 34190 40910 34242 40962
rect 34750 40910 34802 40962
rect 36206 40910 36258 40962
rect 43150 40910 43202 40962
rect 45950 40910 46002 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 16270 40574 16322 40626
rect 16718 40574 16770 40626
rect 22206 40574 22258 40626
rect 23550 40574 23602 40626
rect 24446 40574 24498 40626
rect 28590 40574 28642 40626
rect 30606 40574 30658 40626
rect 32174 40574 32226 40626
rect 33182 40574 33234 40626
rect 33854 40574 33906 40626
rect 35198 40574 35250 40626
rect 36766 40574 36818 40626
rect 40350 40574 40402 40626
rect 45614 40574 45666 40626
rect 11230 40462 11282 40514
rect 15038 40462 15090 40514
rect 15710 40462 15762 40514
rect 15822 40462 15874 40514
rect 17502 40462 17554 40514
rect 18958 40462 19010 40514
rect 21646 40462 21698 40514
rect 22878 40462 22930 40514
rect 23214 40462 23266 40514
rect 29374 40462 29426 40514
rect 30494 40462 30546 40514
rect 30718 40462 30770 40514
rect 35086 40462 35138 40514
rect 35534 40462 35586 40514
rect 35870 40462 35922 40514
rect 41694 40462 41746 40514
rect 45838 40462 45890 40514
rect 6078 40350 6130 40402
rect 9774 40350 9826 40402
rect 10110 40350 10162 40402
rect 11790 40350 11842 40402
rect 15486 40350 15538 40402
rect 16830 40350 16882 40402
rect 18734 40350 18786 40402
rect 20190 40350 20242 40402
rect 21870 40350 21922 40402
rect 23662 40350 23714 40402
rect 24110 40350 24162 40402
rect 27358 40350 27410 40402
rect 28030 40350 28082 40402
rect 30382 40350 30434 40402
rect 30942 40350 30994 40402
rect 31278 40350 31330 40402
rect 31838 40350 31890 40402
rect 31950 40350 32002 40402
rect 32398 40350 32450 40402
rect 33406 40350 33458 40402
rect 34302 40350 34354 40402
rect 37886 40350 37938 40402
rect 38894 40350 38946 40402
rect 39118 40350 39170 40402
rect 39342 40350 39394 40402
rect 39454 40350 39506 40402
rect 40126 40350 40178 40402
rect 41022 40350 41074 40402
rect 44718 40350 44770 40402
rect 45054 40350 45106 40402
rect 45166 40350 45218 40402
rect 45390 40350 45442 40402
rect 45950 40350 46002 40402
rect 6862 40238 6914 40290
rect 8990 40238 9042 40290
rect 10670 40238 10722 40290
rect 11118 40238 11170 40290
rect 11454 40238 11506 40290
rect 12574 40238 12626 40290
rect 14702 40238 14754 40290
rect 17614 40238 17666 40290
rect 22542 40238 22594 40290
rect 25230 40238 25282 40290
rect 29710 40238 29762 40290
rect 29822 40238 29874 40290
rect 31390 40238 31442 40290
rect 32286 40238 32338 40290
rect 34862 40238 34914 40290
rect 36878 40238 36930 40290
rect 37214 40238 37266 40290
rect 38110 40238 38162 40290
rect 43822 40238 43874 40290
rect 15150 40126 15202 40178
rect 16718 40126 16770 40178
rect 17726 40126 17778 40178
rect 28590 40126 28642 40178
rect 28702 40126 28754 40178
rect 28926 40126 28978 40178
rect 29486 40126 29538 40178
rect 33070 40126 33122 40178
rect 33630 40126 33682 40178
rect 34190 40126 34242 40178
rect 39006 40126 39058 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 10222 39790 10274 39842
rect 10558 39790 10610 39842
rect 11006 39790 11058 39842
rect 11790 39790 11842 39842
rect 13470 39790 13522 39842
rect 18286 39790 18338 39842
rect 21422 39790 21474 39842
rect 30270 39790 30322 39842
rect 31166 39790 31218 39842
rect 34078 39790 34130 39842
rect 36990 39790 37042 39842
rect 37326 39790 37378 39842
rect 4622 39678 4674 39730
rect 11118 39678 11170 39730
rect 15710 39678 15762 39730
rect 17278 39678 17330 39730
rect 18398 39678 18450 39730
rect 24670 39678 24722 39730
rect 25006 39678 25058 39730
rect 27134 39678 27186 39730
rect 29710 39678 29762 39730
rect 32958 39678 33010 39730
rect 34190 39678 34242 39730
rect 37774 39678 37826 39730
rect 41918 39678 41970 39730
rect 1822 39566 1874 39618
rect 8094 39566 8146 39618
rect 8318 39566 8370 39618
rect 9662 39566 9714 39618
rect 11902 39566 11954 39618
rect 12910 39566 12962 39618
rect 13470 39566 13522 39618
rect 14142 39566 14194 39618
rect 15486 39566 15538 39618
rect 17166 39566 17218 39618
rect 18174 39566 18226 39618
rect 19070 39566 19122 39618
rect 19294 39566 19346 39618
rect 20078 39566 20130 39618
rect 20526 39566 20578 39618
rect 21870 39566 21922 39618
rect 27918 39566 27970 39618
rect 28254 39566 28306 39618
rect 29822 39566 29874 39618
rect 29934 39566 29986 39618
rect 31166 39566 31218 39618
rect 31614 39566 31666 39618
rect 32510 39566 32562 39618
rect 32734 39566 32786 39618
rect 33070 39566 33122 39618
rect 33518 39566 33570 39618
rect 34974 39566 35026 39618
rect 35758 39566 35810 39618
rect 38670 39566 38722 39618
rect 40686 39566 40738 39618
rect 43038 39566 43090 39618
rect 43374 39566 43426 39618
rect 44270 39566 44322 39618
rect 44830 39566 44882 39618
rect 45614 39566 45666 39618
rect 2494 39454 2546 39506
rect 7758 39454 7810 39506
rect 10334 39454 10386 39506
rect 11230 39454 11282 39506
rect 13806 39454 13858 39506
rect 14814 39454 14866 39506
rect 16158 39454 16210 39506
rect 19630 39454 19682 39506
rect 21310 39454 21362 39506
rect 22542 39454 22594 39506
rect 30606 39454 30658 39506
rect 31726 39454 31778 39506
rect 32286 39454 32338 39506
rect 33182 39454 33234 39506
rect 33630 39454 33682 39506
rect 35198 39454 35250 39506
rect 35534 39454 35586 39506
rect 38782 39454 38834 39506
rect 41246 39454 41298 39506
rect 42814 39454 42866 39506
rect 44046 39454 44098 39506
rect 7086 39342 7138 39394
rect 7422 39342 7474 39394
rect 7870 39342 7922 39394
rect 8654 39342 8706 39394
rect 8766 39342 8818 39394
rect 8878 39342 8930 39394
rect 9438 39342 9490 39394
rect 9774 39342 9826 39394
rect 9998 39342 10050 39394
rect 12574 39342 12626 39394
rect 14478 39342 14530 39394
rect 16494 39342 16546 39394
rect 28590 39342 28642 39394
rect 29598 39342 29650 39394
rect 30830 39342 30882 39394
rect 31054 39342 31106 39394
rect 31950 39342 32002 39394
rect 33854 39342 33906 39394
rect 34638 39342 34690 39394
rect 36094 39342 36146 39394
rect 37102 39342 37154 39394
rect 38334 39342 38386 39394
rect 45166 39342 45218 39394
rect 46174 39342 46226 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 13134 39006 13186 39058
rect 14142 39006 14194 39058
rect 17390 39006 17442 39058
rect 23102 39006 23154 39058
rect 23214 39006 23266 39058
rect 23438 39006 23490 39058
rect 24334 39006 24386 39058
rect 26686 39006 26738 39058
rect 27358 39006 27410 39058
rect 27470 39006 27522 39058
rect 27582 39006 27634 39058
rect 29822 39006 29874 39058
rect 32174 39006 32226 39058
rect 33070 39006 33122 39058
rect 33630 39006 33682 39058
rect 35086 39006 35138 39058
rect 40014 39006 40066 39058
rect 41022 39006 41074 39058
rect 45054 39006 45106 39058
rect 2830 38894 2882 38946
rect 3502 38894 3554 38946
rect 4174 38894 4226 38946
rect 6078 38894 6130 38946
rect 8990 38894 9042 38946
rect 13806 38894 13858 38946
rect 16606 38894 16658 38946
rect 22878 38894 22930 38946
rect 23326 38894 23378 38946
rect 24110 38894 24162 38946
rect 24670 38894 24722 38946
rect 28030 38894 28082 38946
rect 29374 38894 29426 38946
rect 31726 38894 31778 38946
rect 34302 38894 34354 38946
rect 36542 38894 36594 38946
rect 40238 38894 40290 38946
rect 40350 38894 40402 38946
rect 43486 38894 43538 38946
rect 44942 38894 44994 38946
rect 45950 38894 46002 38946
rect 3726 38782 3778 38834
rect 3950 38782 4002 38834
rect 4286 38782 4338 38834
rect 5294 38782 5346 38834
rect 8654 38782 8706 38834
rect 9886 38782 9938 38834
rect 13022 38782 13074 38834
rect 13470 38782 13522 38834
rect 14478 38782 14530 38834
rect 15710 38782 15762 38834
rect 16046 38782 16098 38834
rect 17726 38782 17778 38834
rect 19182 38782 19234 38834
rect 20190 38782 20242 38834
rect 20862 38782 20914 38834
rect 21310 38782 21362 38834
rect 24446 38782 24498 38834
rect 25902 38782 25954 38834
rect 27022 38782 27074 38834
rect 27246 38782 27298 38834
rect 28366 38782 28418 38834
rect 28702 38782 28754 38834
rect 28926 38782 28978 38834
rect 29262 38782 29314 38834
rect 30494 38782 30546 38834
rect 30718 38782 30770 38834
rect 30942 38782 30994 38834
rect 33854 38782 33906 38834
rect 34414 38782 34466 38834
rect 34638 38782 34690 38834
rect 34974 38782 35026 38834
rect 35758 38782 35810 38834
rect 39118 38782 39170 38834
rect 39342 38782 39394 38834
rect 40910 38782 40962 38834
rect 44158 38782 44210 38834
rect 45166 38782 45218 38834
rect 45614 38782 45666 38834
rect 2718 38670 2770 38722
rect 3054 38670 3106 38722
rect 8206 38670 8258 38722
rect 10558 38670 10610 38722
rect 12686 38670 12738 38722
rect 15150 38670 15202 38722
rect 15262 38670 15314 38722
rect 15486 38670 15538 38722
rect 16494 38670 16546 38722
rect 16830 38670 16882 38722
rect 18734 38670 18786 38722
rect 20638 38670 20690 38722
rect 25230 38670 25282 38722
rect 26126 38670 26178 38722
rect 29150 38670 29202 38722
rect 33182 38670 33234 38722
rect 38670 38670 38722 38722
rect 39230 38670 39282 38722
rect 39566 38670 39618 38722
rect 39790 38670 39842 38722
rect 41358 38670 41410 38722
rect 3390 38558 3442 38610
rect 16158 38558 16210 38610
rect 28142 38558 28194 38610
rect 31390 38558 31442 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 4398 38222 4450 38274
rect 21758 38222 21810 38274
rect 27246 38222 27298 38274
rect 32510 38222 32562 38274
rect 35198 38222 35250 38274
rect 3614 38110 3666 38162
rect 11342 38110 11394 38162
rect 20078 38110 20130 38162
rect 25118 38110 25170 38162
rect 25454 38110 25506 38162
rect 27358 38110 27410 38162
rect 29486 38110 29538 38162
rect 34526 38110 34578 38162
rect 39790 38110 39842 38162
rect 41918 38110 41970 38162
rect 43374 38110 43426 38162
rect 44942 38110 44994 38162
rect 45950 38110 46002 38162
rect 3390 37998 3442 38050
rect 4286 37998 4338 38050
rect 10110 37998 10162 38050
rect 11118 37998 11170 38050
rect 11566 37998 11618 38050
rect 11790 37998 11842 38050
rect 18062 37998 18114 38050
rect 19070 37998 19122 38050
rect 20302 37998 20354 38050
rect 21310 37998 21362 38050
rect 22542 37998 22594 38050
rect 24446 37998 24498 38050
rect 25790 37998 25842 38050
rect 26686 37998 26738 38050
rect 27694 37998 27746 38050
rect 28030 37998 28082 38050
rect 29374 37998 29426 38050
rect 29598 37998 29650 38050
rect 29822 37998 29874 38050
rect 30158 37998 30210 38050
rect 30494 37998 30546 38050
rect 30718 37998 30770 38050
rect 31054 37998 31106 38050
rect 31390 37998 31442 38050
rect 31838 37998 31890 38050
rect 32734 37998 32786 38050
rect 34414 37998 34466 38050
rect 34974 37998 35026 38050
rect 35982 37998 36034 38050
rect 36094 37998 36146 38050
rect 37886 37998 37938 38050
rect 38334 37998 38386 38050
rect 38894 37998 38946 38050
rect 39342 37998 39394 38050
rect 42702 37998 42754 38050
rect 43038 37998 43090 38050
rect 43486 37998 43538 38050
rect 43710 37998 43762 38050
rect 45054 37998 45106 38050
rect 45278 37998 45330 38050
rect 45390 37998 45442 38050
rect 3950 37886 4002 37938
rect 5854 37886 5906 37938
rect 12574 37886 12626 37938
rect 12798 37886 12850 37938
rect 13694 37886 13746 37938
rect 20414 37886 20466 37938
rect 23886 37886 23938 37938
rect 26798 37886 26850 37938
rect 28254 37886 28306 37938
rect 29150 37886 29202 37938
rect 33966 37886 34018 37938
rect 35534 37886 35586 37938
rect 35870 37886 35922 37938
rect 36430 37886 36482 37938
rect 37326 37886 37378 37938
rect 38558 37886 38610 37938
rect 44046 37886 44098 37938
rect 44158 37886 44210 37938
rect 45838 37886 45890 37938
rect 46062 37886 46114 37938
rect 4398 37774 4450 37826
rect 12350 37774 12402 37826
rect 12686 37774 12738 37826
rect 19294 37774 19346 37826
rect 26014 37774 26066 37826
rect 28142 37774 28194 37826
rect 28366 37774 28418 37826
rect 30270 37774 30322 37826
rect 30830 37774 30882 37826
rect 33182 37774 33234 37826
rect 33518 37774 33570 37826
rect 34190 37774 34242 37826
rect 34526 37774 34578 37826
rect 37214 37774 37266 37826
rect 43262 37774 43314 37826
rect 44382 37774 44434 37826
rect 44942 37774 44994 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5070 37438 5122 37490
rect 5182 37438 5234 37490
rect 8990 37438 9042 37490
rect 12910 37438 12962 37490
rect 17502 37438 17554 37490
rect 22878 37438 22930 37490
rect 23662 37438 23714 37490
rect 27806 37438 27858 37490
rect 30830 37438 30882 37490
rect 31390 37438 31442 37490
rect 38894 37438 38946 37490
rect 6414 37326 6466 37378
rect 8878 37326 8930 37378
rect 9550 37326 9602 37378
rect 10446 37326 10498 37378
rect 14254 37326 14306 37378
rect 18398 37326 18450 37378
rect 24110 37326 24162 37378
rect 24222 37326 24274 37378
rect 26686 37326 26738 37378
rect 29934 37326 29986 37378
rect 39790 37326 39842 37378
rect 4622 37214 4674 37266
rect 5742 37214 5794 37266
rect 9886 37214 9938 37266
rect 10782 37214 10834 37266
rect 11790 37214 11842 37266
rect 12574 37214 12626 37266
rect 13470 37214 13522 37266
rect 16942 37214 16994 37266
rect 17726 37214 17778 37266
rect 18174 37214 18226 37266
rect 21982 37214 22034 37266
rect 22654 37214 22706 37266
rect 23326 37214 23378 37266
rect 24670 37214 24722 37266
rect 26126 37214 26178 37266
rect 28142 37214 28194 37266
rect 31278 37214 31330 37266
rect 35310 37214 35362 37266
rect 39006 37214 39058 37266
rect 39566 37214 39618 37266
rect 41806 37214 41858 37266
rect 1710 37102 1762 37154
rect 3838 37102 3890 37154
rect 8542 37102 8594 37154
rect 10110 37102 10162 37154
rect 12014 37102 12066 37154
rect 12350 37102 12402 37154
rect 16382 37102 16434 37154
rect 18510 37102 18562 37154
rect 19182 37102 19234 37154
rect 21310 37102 21362 37154
rect 25454 37102 25506 37154
rect 30270 37102 30322 37154
rect 30382 37102 30434 37154
rect 31838 37102 31890 37154
rect 32398 37102 32450 37154
rect 33294 37102 33346 37154
rect 33742 37102 33794 37154
rect 34078 37102 34130 37154
rect 34526 37102 34578 37154
rect 35982 37102 36034 37154
rect 38110 37102 38162 37154
rect 39454 37102 39506 37154
rect 43374 37102 43426 37154
rect 4958 36990 5010 37042
rect 11454 36990 11506 37042
rect 24110 36990 24162 37042
rect 31726 36990 31778 37042
rect 32510 36990 32562 37042
rect 33966 36990 34018 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 3614 36654 3666 36706
rect 8878 36654 8930 36706
rect 3838 36542 3890 36594
rect 5630 36542 5682 36594
rect 12462 36542 12514 36594
rect 14254 36542 14306 36594
rect 16382 36542 16434 36594
rect 19854 36542 19906 36594
rect 20190 36542 20242 36594
rect 21422 36542 21474 36594
rect 21870 36542 21922 36594
rect 22094 36542 22146 36594
rect 27246 36542 27298 36594
rect 29262 36542 29314 36594
rect 31502 36542 31554 36594
rect 33630 36542 33682 36594
rect 36206 36542 36258 36594
rect 37998 36542 38050 36594
rect 40238 36542 40290 36594
rect 42366 36542 42418 36594
rect 2830 36430 2882 36482
rect 3054 36430 3106 36482
rect 3278 36430 3330 36482
rect 4958 36430 5010 36482
rect 8542 36430 8594 36482
rect 9662 36430 9714 36482
rect 13470 36430 13522 36482
rect 16718 36430 16770 36482
rect 17054 36430 17106 36482
rect 17390 36430 17442 36482
rect 18286 36430 18338 36482
rect 20750 36430 20802 36482
rect 21870 36430 21922 36482
rect 22318 36430 22370 36482
rect 23214 36430 23266 36482
rect 23550 36430 23602 36482
rect 23886 36430 23938 36482
rect 26910 36430 26962 36482
rect 30830 36430 30882 36482
rect 34974 36430 35026 36482
rect 38446 36430 38498 36482
rect 39454 36430 39506 36482
rect 40574 36430 40626 36482
rect 41470 36430 41522 36482
rect 42478 36430 42530 36482
rect 2718 36318 2770 36370
rect 7758 36318 7810 36370
rect 9102 36318 9154 36370
rect 10334 36318 10386 36370
rect 18398 36318 18450 36370
rect 18510 36318 18562 36370
rect 18958 36318 19010 36370
rect 19182 36318 19234 36370
rect 19518 36318 19570 36370
rect 20638 36318 20690 36370
rect 22654 36318 22706 36370
rect 23662 36318 23714 36370
rect 26014 36318 26066 36370
rect 29598 36318 29650 36370
rect 29822 36318 29874 36370
rect 30270 36318 30322 36370
rect 34414 36318 34466 36370
rect 35310 36318 35362 36370
rect 36430 36318 36482 36370
rect 41918 36318 41970 36370
rect 43598 36542 43650 36594
rect 45502 36542 45554 36594
rect 42814 36430 42866 36482
rect 43934 36430 43986 36482
rect 45166 36430 45218 36482
rect 42814 36318 42866 36370
rect 43822 36318 43874 36370
rect 44830 36318 44882 36370
rect 46174 36318 46226 36370
rect 3838 36206 3890 36258
rect 4734 36206 4786 36258
rect 8990 36206 9042 36258
rect 13022 36206 13074 36258
rect 17166 36206 17218 36258
rect 17278 36206 17330 36258
rect 17838 36206 17890 36258
rect 19406 36206 19458 36258
rect 20414 36206 20466 36258
rect 21310 36206 21362 36258
rect 21534 36206 21586 36258
rect 22542 36206 22594 36258
rect 22878 36206 22930 36258
rect 23102 36206 23154 36258
rect 24446 36206 24498 36258
rect 25230 36206 25282 36258
rect 26910 36206 26962 36258
rect 28702 36206 28754 36258
rect 29262 36206 29314 36258
rect 29374 36206 29426 36258
rect 30158 36206 30210 36258
rect 34302 36206 34354 36258
rect 34638 36206 34690 36258
rect 34862 36206 34914 36258
rect 35422 36206 35474 36258
rect 35646 36206 35698 36258
rect 41806 36206 41858 36258
rect 42030 36206 42082 36258
rect 43038 36206 43090 36258
rect 44942 36206 44994 36258
rect 45390 36206 45442 36258
rect 45838 36206 45890 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 5854 35870 5906 35922
rect 6974 35870 7026 35922
rect 15710 35870 15762 35922
rect 16494 35870 16546 35922
rect 25230 35870 25282 35922
rect 27134 35870 27186 35922
rect 31054 35870 31106 35922
rect 31278 35870 31330 35922
rect 32174 35870 32226 35922
rect 36990 35870 37042 35922
rect 41022 35870 41074 35922
rect 2494 35758 2546 35810
rect 5742 35758 5794 35810
rect 7870 35758 7922 35810
rect 16830 35758 16882 35810
rect 17502 35758 17554 35810
rect 28254 35758 28306 35810
rect 30718 35758 30770 35810
rect 31166 35758 31218 35810
rect 32510 35758 32562 35810
rect 33854 35758 33906 35810
rect 40910 35758 40962 35810
rect 1822 35646 1874 35698
rect 6750 35646 6802 35698
rect 7758 35646 7810 35698
rect 8430 35646 8482 35698
rect 8990 35646 9042 35698
rect 14702 35646 14754 35698
rect 15374 35646 15426 35698
rect 15598 35646 15650 35698
rect 15710 35646 15762 35698
rect 17614 35646 17666 35698
rect 17950 35646 18002 35698
rect 20414 35646 20466 35698
rect 25342 35646 25394 35698
rect 26238 35646 26290 35698
rect 26686 35646 26738 35698
rect 27470 35646 27522 35698
rect 30942 35646 30994 35698
rect 31838 35646 31890 35698
rect 32062 35646 32114 35698
rect 32286 35646 32338 35698
rect 33070 35646 33122 35698
rect 36654 35646 36706 35698
rect 36878 35646 36930 35698
rect 37214 35646 37266 35698
rect 37550 35646 37602 35698
rect 41246 35646 41298 35698
rect 42254 35646 42306 35698
rect 42926 35646 42978 35698
rect 43374 35646 43426 35698
rect 4622 35534 4674 35586
rect 5294 35534 5346 35586
rect 5966 35534 6018 35586
rect 6526 35534 6578 35586
rect 6862 35534 6914 35586
rect 7646 35534 7698 35586
rect 9774 35534 9826 35586
rect 21870 35534 21922 35586
rect 25902 35534 25954 35586
rect 30382 35534 30434 35586
rect 35982 35534 36034 35586
rect 38222 35534 38274 35586
rect 40350 35534 40402 35586
rect 42142 35534 42194 35586
rect 44046 35534 44098 35586
rect 46174 35534 46226 35586
rect 5182 35422 5234 35474
rect 6302 35422 6354 35474
rect 42030 35422 42082 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 7198 35086 7250 35138
rect 29374 35086 29426 35138
rect 35534 35086 35586 35138
rect 36094 35086 36146 35138
rect 37550 35086 37602 35138
rect 43150 35086 43202 35138
rect 44942 35086 44994 35138
rect 3054 34974 3106 35026
rect 4846 34974 4898 35026
rect 8094 34974 8146 35026
rect 9662 34974 9714 35026
rect 13694 34974 13746 35026
rect 15822 34974 15874 35026
rect 17838 34974 17890 35026
rect 24670 34974 24722 35026
rect 27918 34974 27970 35026
rect 30270 34974 30322 35026
rect 35870 34974 35922 35026
rect 36318 34974 36370 35026
rect 38446 34974 38498 35026
rect 39566 34974 39618 35026
rect 46174 34974 46226 35026
rect 3278 34862 3330 34914
rect 3950 34862 4002 34914
rect 4062 34862 4114 34914
rect 4398 34862 4450 34914
rect 7646 34862 7698 34914
rect 7870 34862 7922 34914
rect 8766 34862 8818 34914
rect 12574 34862 12626 34914
rect 16606 34862 16658 34914
rect 16942 34862 16994 34914
rect 20638 34862 20690 34914
rect 21870 34862 21922 34914
rect 25118 34862 25170 34914
rect 34750 34862 34802 34914
rect 35646 34862 35698 34914
rect 37214 34862 37266 34914
rect 37774 34862 37826 34914
rect 39006 34862 39058 34914
rect 41134 34862 41186 34914
rect 43710 34862 43762 34914
rect 43934 34862 43986 34914
rect 45390 34862 45442 34914
rect 45614 34862 45666 34914
rect 2942 34750 2994 34802
rect 3502 34750 3554 34802
rect 4286 34750 4338 34802
rect 7198 34750 7250 34802
rect 7310 34750 7362 34802
rect 9326 34750 9378 34802
rect 11790 34750 11842 34802
rect 19966 34750 20018 34802
rect 22542 34750 22594 34802
rect 25790 34750 25842 34802
rect 29262 34750 29314 34802
rect 36990 34750 37042 34802
rect 37326 34750 37378 34802
rect 38670 34750 38722 34802
rect 39678 34750 39730 34802
rect 42702 34750 42754 34802
rect 43374 34750 43426 34802
rect 43486 34750 43538 34802
rect 44830 34750 44882 34802
rect 45054 34750 45106 34802
rect 17278 34638 17330 34690
rect 21534 34638 21586 34690
rect 28590 34638 28642 34690
rect 46062 34638 46114 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2830 34302 2882 34354
rect 2942 34302 2994 34354
rect 3950 34302 4002 34354
rect 5070 34302 5122 34354
rect 7870 34302 7922 34354
rect 9102 34302 9154 34354
rect 9886 34302 9938 34354
rect 9998 34302 10050 34354
rect 10446 34302 10498 34354
rect 11118 34302 11170 34354
rect 11902 34302 11954 34354
rect 12014 34302 12066 34354
rect 12574 34302 12626 34354
rect 13022 34302 13074 34354
rect 13806 34302 13858 34354
rect 14926 34302 14978 34354
rect 16494 34302 16546 34354
rect 17390 34302 17442 34354
rect 19070 34302 19122 34354
rect 19294 34302 19346 34354
rect 20414 34302 20466 34354
rect 21422 34302 21474 34354
rect 22654 34302 22706 34354
rect 22990 34302 23042 34354
rect 25342 34302 25394 34354
rect 26350 34302 26402 34354
rect 26910 34302 26962 34354
rect 27358 34302 27410 34354
rect 27806 34302 27858 34354
rect 32174 34302 32226 34354
rect 33294 34302 33346 34354
rect 33406 34302 33458 34354
rect 35534 34302 35586 34354
rect 40238 34302 40290 34354
rect 44830 34302 44882 34354
rect 4398 34190 4450 34242
rect 4622 34190 4674 34242
rect 6302 34190 6354 34242
rect 6862 34190 6914 34242
rect 7422 34190 7474 34242
rect 8206 34190 8258 34242
rect 11454 34190 11506 34242
rect 11678 34190 11730 34242
rect 18958 34190 19010 34242
rect 20750 34190 20802 34242
rect 20862 34190 20914 34242
rect 24334 34190 24386 34242
rect 24446 34190 24498 34242
rect 25230 34190 25282 34242
rect 26462 34190 26514 34242
rect 32510 34190 32562 34242
rect 33518 34190 33570 34242
rect 34078 34190 34130 34242
rect 34862 34190 34914 34242
rect 35198 34190 35250 34242
rect 35310 34190 35362 34242
rect 36542 34190 36594 34242
rect 39006 34190 39058 34242
rect 39342 34190 39394 34242
rect 40350 34190 40402 34242
rect 41694 34190 41746 34242
rect 44270 34190 44322 34242
rect 46174 34190 46226 34242
rect 1934 34078 1986 34130
rect 2158 34078 2210 34130
rect 2494 34078 2546 34130
rect 2718 34078 2770 34130
rect 3278 34078 3330 34130
rect 4510 34078 4562 34130
rect 5294 34078 5346 34130
rect 5854 34078 5906 34130
rect 6414 34078 6466 34130
rect 6974 34078 7026 34130
rect 7198 34078 7250 34130
rect 7758 34078 7810 34130
rect 7982 34078 8034 34130
rect 9438 34078 9490 34130
rect 10110 34078 10162 34130
rect 10558 34078 10610 34130
rect 13358 34078 13410 34130
rect 13582 34078 13634 34130
rect 13918 34078 13970 34130
rect 21086 34078 21138 34130
rect 21310 34078 21362 34130
rect 21534 34078 21586 34130
rect 21982 34078 22034 34130
rect 22318 34078 22370 34130
rect 23326 34078 23378 34130
rect 23774 34078 23826 34130
rect 24110 34078 24162 34130
rect 31166 34078 31218 34130
rect 31838 34078 31890 34130
rect 32062 34078 32114 34130
rect 32286 34078 32338 34130
rect 33070 34078 33122 34130
rect 33630 34078 33682 34130
rect 34414 34078 34466 34130
rect 35870 34078 35922 34130
rect 39118 34078 39170 34130
rect 39566 34078 39618 34130
rect 40910 34078 40962 34130
rect 44158 34078 44210 34130
rect 44494 34078 44546 34130
rect 45166 34078 45218 34130
rect 45614 34078 45666 34130
rect 2270 33966 2322 34018
rect 6078 33966 6130 34018
rect 11006 33966 11058 34018
rect 11790 33966 11842 34018
rect 13694 33966 13746 34018
rect 14590 33966 14642 34018
rect 15486 33966 15538 34018
rect 15934 33966 15986 34018
rect 16942 33966 16994 34018
rect 17502 33966 17554 34018
rect 18062 33966 18114 34018
rect 18622 33966 18674 34018
rect 19966 33966 20018 34018
rect 26014 33966 26066 34018
rect 28366 33966 28418 34018
rect 30494 33966 30546 34018
rect 38670 33966 38722 34018
rect 43822 33966 43874 34018
rect 45502 33966 45554 34018
rect 17950 33854 18002 33906
rect 23102 33854 23154 33906
rect 23886 33854 23938 33906
rect 25342 33854 25394 33906
rect 25902 33854 25954 33906
rect 34750 33854 34802 33906
rect 39790 33854 39842 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 10782 33518 10834 33570
rect 21646 33518 21698 33570
rect 2494 33406 2546 33458
rect 4622 33406 4674 33458
rect 6414 33406 6466 33458
rect 8542 33406 8594 33458
rect 9438 33406 9490 33458
rect 1822 33294 1874 33346
rect 5630 33294 5682 33346
rect 9998 33294 10050 33346
rect 10334 33294 10386 33346
rect 21982 33518 22034 33570
rect 44830 33518 44882 33570
rect 44942 33518 44994 33570
rect 45390 33518 45442 33570
rect 45614 33518 45666 33570
rect 46062 33518 46114 33570
rect 11790 33406 11842 33458
rect 12798 33406 12850 33458
rect 16382 33406 16434 33458
rect 17502 33406 17554 33458
rect 19630 33406 19682 33458
rect 25454 33406 25506 33458
rect 27582 33406 27634 33458
rect 28254 33406 28306 33458
rect 30046 33406 30098 33458
rect 32734 33406 32786 33458
rect 34862 33406 34914 33458
rect 40462 33406 40514 33458
rect 46174 33406 46226 33458
rect 13470 33294 13522 33346
rect 16830 33294 16882 33346
rect 21982 33294 22034 33346
rect 22430 33294 22482 33346
rect 22990 33294 23042 33346
rect 24782 33294 24834 33346
rect 27918 33294 27970 33346
rect 28366 33294 28418 33346
rect 28590 33294 28642 33346
rect 29486 33294 29538 33346
rect 30158 33294 30210 33346
rect 31502 33294 31554 33346
rect 31950 33294 32002 33346
rect 35422 33294 35474 33346
rect 37214 33294 37266 33346
rect 42814 33294 42866 33346
rect 14254 33182 14306 33234
rect 20414 33182 20466 33234
rect 22766 33182 22818 33234
rect 23326 33182 23378 33234
rect 24222 33182 24274 33234
rect 28142 33182 28194 33234
rect 29710 33182 29762 33234
rect 30494 33182 30546 33234
rect 31166 33182 31218 33234
rect 35198 33182 35250 33234
rect 36206 33182 36258 33234
rect 36990 33182 37042 33234
rect 38670 33182 38722 33234
rect 45054 33182 45106 33234
rect 10894 33070 10946 33122
rect 11118 33070 11170 33122
rect 12238 33070 12290 33122
rect 12910 33070 12962 33122
rect 20862 33070 20914 33122
rect 22542 33070 22594 33122
rect 23662 33070 23714 33122
rect 23886 33070 23938 33122
rect 24110 33070 24162 33122
rect 29934 33070 29986 33122
rect 30830 33070 30882 33122
rect 36094 33070 36146 33122
rect 37662 33070 37714 33122
rect 37998 33070 38050 33122
rect 38334 33070 38386 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 11342 32734 11394 32786
rect 15374 32734 15426 32786
rect 16494 32734 16546 32786
rect 17502 32734 17554 32786
rect 18286 32734 18338 32786
rect 19406 32734 19458 32786
rect 23326 32734 23378 32786
rect 23886 32734 23938 32786
rect 29150 32734 29202 32786
rect 30382 32734 30434 32786
rect 31278 32734 31330 32786
rect 31950 32734 32002 32786
rect 39790 32734 39842 32786
rect 41918 32734 41970 32786
rect 42142 32734 42194 32786
rect 14030 32622 14082 32674
rect 15598 32622 15650 32674
rect 16046 32622 16098 32674
rect 17390 32622 17442 32674
rect 18622 32622 18674 32674
rect 19070 32622 19122 32674
rect 26350 32622 26402 32674
rect 29598 32622 29650 32674
rect 33742 32622 33794 32674
rect 37886 32622 37938 32674
rect 41806 32622 41858 32674
rect 7534 32510 7586 32562
rect 10894 32510 10946 32562
rect 11118 32510 11170 32562
rect 11566 32510 11618 32562
rect 14814 32510 14866 32562
rect 15486 32510 15538 32562
rect 16270 32510 16322 32562
rect 16382 32510 16434 32562
rect 16606 32510 16658 32562
rect 16718 32510 16770 32562
rect 17950 32510 18002 32562
rect 18174 32510 18226 32562
rect 18398 32510 18450 32562
rect 19742 32510 19794 32562
rect 22990 32510 23042 32562
rect 23326 32510 23378 32562
rect 23550 32510 23602 32562
rect 24222 32510 24274 32562
rect 24558 32510 24610 32562
rect 25454 32510 25506 32562
rect 26574 32510 26626 32562
rect 27358 32510 27410 32562
rect 27582 32510 27634 32562
rect 27806 32510 27858 32562
rect 30942 32510 30994 32562
rect 31726 32510 31778 32562
rect 32174 32510 32226 32562
rect 32398 32510 32450 32562
rect 33406 32510 33458 32562
rect 34078 32510 34130 32562
rect 34750 32510 34802 32562
rect 38110 32510 38162 32562
rect 38446 32510 38498 32562
rect 38894 32510 38946 32562
rect 39006 32510 39058 32562
rect 39454 32510 39506 32562
rect 42478 32510 42530 32562
rect 43374 32510 43426 32562
rect 7982 32398 8034 32450
rect 10558 32398 10610 32450
rect 11006 32398 11058 32450
rect 11902 32398 11954 32450
rect 20526 32398 20578 32450
rect 22654 32398 22706 32450
rect 25902 32398 25954 32450
rect 27694 32398 27746 32450
rect 28254 32398 28306 32450
rect 28814 32398 28866 32450
rect 30494 32398 30546 32450
rect 32286 32398 32338 32450
rect 35422 32398 35474 32450
rect 37550 32398 37602 32450
rect 37998 32398 38050 32450
rect 39230 32398 39282 32450
rect 40238 32398 40290 32450
rect 41022 32398 41074 32450
rect 41470 32398 41522 32450
rect 42814 32398 42866 32450
rect 44046 32398 44098 32450
rect 46174 32398 46226 32450
rect 8766 32286 8818 32338
rect 10446 32286 10498 32338
rect 24670 32286 24722 32338
rect 30158 32286 30210 32338
rect 33070 32286 33122 32338
rect 33406 32286 33458 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 16830 31950 16882 32002
rect 18286 31950 18338 32002
rect 28030 31950 28082 32002
rect 4622 31838 4674 31890
rect 9550 31838 9602 31890
rect 11678 31838 11730 31890
rect 16270 31838 16322 31890
rect 16830 31838 16882 31890
rect 19854 31838 19906 31890
rect 27358 31838 27410 31890
rect 29262 31838 29314 31890
rect 29710 31838 29762 31890
rect 31054 31838 31106 31890
rect 33182 31838 33234 31890
rect 35646 31838 35698 31890
rect 37102 31838 37154 31890
rect 42142 31838 42194 31890
rect 43822 31838 43874 31890
rect 44942 31838 44994 31890
rect 45390 31838 45442 31890
rect 1822 31726 1874 31778
rect 8430 31726 8482 31778
rect 8878 31726 8930 31778
rect 13918 31726 13970 31778
rect 14142 31726 14194 31778
rect 17278 31726 17330 31778
rect 20190 31726 20242 31778
rect 20862 31726 20914 31778
rect 21310 31726 21362 31778
rect 27246 31726 27298 31778
rect 27470 31726 27522 31778
rect 33966 31726 34018 31778
rect 34302 31726 34354 31778
rect 34862 31726 34914 31778
rect 35534 31726 35586 31778
rect 36094 31726 36146 31778
rect 37326 31726 37378 31778
rect 37662 31726 37714 31778
rect 37886 31726 37938 31778
rect 39342 31726 39394 31778
rect 42478 31726 42530 31778
rect 43038 31726 43090 31778
rect 2494 31614 2546 31666
rect 5854 31614 5906 31666
rect 6302 31614 6354 31666
rect 6638 31614 6690 31666
rect 6862 31614 6914 31666
rect 7198 31614 7250 31666
rect 7422 31614 7474 31666
rect 7758 31614 7810 31666
rect 13470 31614 13522 31666
rect 14478 31614 14530 31666
rect 15822 31614 15874 31666
rect 18510 31614 18562 31666
rect 19406 31614 19458 31666
rect 20414 31614 20466 31666
rect 23326 31614 23378 31666
rect 27022 31614 27074 31666
rect 28142 31614 28194 31666
rect 28590 31614 28642 31666
rect 30382 31614 30434 31666
rect 30718 31614 30770 31666
rect 35870 31614 35922 31666
rect 37550 31614 37602 31666
rect 38670 31614 38722 31666
rect 40014 31614 40066 31666
rect 5518 31502 5570 31554
rect 5742 31502 5794 31554
rect 6414 31502 6466 31554
rect 6974 31502 7026 31554
rect 7870 31502 7922 31554
rect 8094 31502 8146 31554
rect 12574 31502 12626 31554
rect 13022 31502 13074 31554
rect 13694 31502 13746 31554
rect 13806 31502 13858 31554
rect 14814 31502 14866 31554
rect 15486 31502 15538 31554
rect 15710 31502 15762 31554
rect 17838 31502 17890 31554
rect 18174 31502 18226 31554
rect 18622 31502 18674 31554
rect 20526 31502 20578 31554
rect 28366 31502 28418 31554
rect 38334 31502 38386 31554
rect 43374 31502 43426 31554
rect 45950 31502 46002 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 9550 31166 9602 31218
rect 21422 31166 21474 31218
rect 34078 31166 34130 31218
rect 41022 31166 41074 31218
rect 41806 31166 41858 31218
rect 42590 31166 42642 31218
rect 44494 31166 44546 31218
rect 44942 31166 44994 31218
rect 45838 31166 45890 31218
rect 5630 31054 5682 31106
rect 8206 31054 8258 31106
rect 8430 31054 8482 31106
rect 14702 31054 14754 31106
rect 19518 31054 19570 31106
rect 21086 31054 21138 31106
rect 22542 31054 22594 31106
rect 26686 31054 26738 31106
rect 27918 31054 27970 31106
rect 29598 31054 29650 31106
rect 33294 31054 33346 31106
rect 42366 31054 42418 31106
rect 43934 31054 43986 31106
rect 45950 31054 46002 31106
rect 7646 30942 7698 30994
rect 8542 30942 8594 30994
rect 9102 30942 9154 30994
rect 9886 30942 9938 30994
rect 13358 30942 13410 30994
rect 14030 30942 14082 30994
rect 20302 30942 20354 30994
rect 21758 30942 21810 30994
rect 25230 30942 25282 30994
rect 28366 30942 28418 30994
rect 28926 30942 28978 30994
rect 32398 30942 32450 30994
rect 33518 30942 33570 30994
rect 39790 30942 39842 30994
rect 41358 30942 41410 30994
rect 41582 30942 41634 30994
rect 42030 30942 42082 30994
rect 43038 30942 43090 30994
rect 43486 30942 43538 30994
rect 10446 30830 10498 30882
rect 12574 30830 12626 30882
rect 16830 30830 16882 30882
rect 17390 30830 17442 30882
rect 20862 30830 20914 30882
rect 24670 30830 24722 30882
rect 26574 30830 26626 30882
rect 31726 30830 31778 30882
rect 32174 30830 32226 30882
rect 35982 30830 36034 30882
rect 40238 30830 40290 30882
rect 40910 30830 40962 30882
rect 41694 30830 41746 30882
rect 45390 30830 45442 30882
rect 32062 30718 32114 30770
rect 40126 30718 40178 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 12014 30382 12066 30434
rect 30830 30382 30882 30434
rect 1710 30270 1762 30322
rect 7422 30270 7474 30322
rect 14030 30270 14082 30322
rect 19406 30270 19458 30322
rect 26798 30270 26850 30322
rect 35198 30270 35250 30322
rect 40462 30270 40514 30322
rect 41582 30270 41634 30322
rect 43710 30270 43762 30322
rect 4622 30158 4674 30210
rect 5854 30158 5906 30210
rect 6190 30158 6242 30210
rect 6414 30158 6466 30210
rect 7086 30158 7138 30210
rect 10334 30158 10386 30210
rect 11230 30158 11282 30210
rect 11902 30158 11954 30210
rect 17278 30158 17330 30210
rect 19070 30158 19122 30210
rect 19294 30158 19346 30210
rect 20414 30158 20466 30210
rect 21310 30158 21362 30210
rect 21982 30158 22034 30210
rect 22766 30158 22818 30210
rect 22990 30158 23042 30210
rect 23326 30158 23378 30210
rect 23886 30158 23938 30210
rect 24558 30158 24610 30210
rect 25902 30158 25954 30210
rect 26686 30158 26738 30210
rect 27246 30158 27298 30210
rect 27582 30158 27634 30210
rect 27806 30158 27858 30210
rect 28478 30158 28530 30210
rect 30158 30158 30210 30210
rect 31838 30158 31890 30210
rect 32398 30158 32450 30210
rect 33742 30158 33794 30210
rect 34302 30158 34354 30210
rect 34862 30158 34914 30210
rect 37550 30158 37602 30210
rect 38334 30158 38386 30210
rect 40798 30158 40850 30210
rect 44046 30158 44098 30210
rect 44942 30158 44994 30210
rect 45390 30158 45442 30210
rect 46174 30158 46226 30210
rect 3838 30046 3890 30098
rect 5630 30046 5682 30098
rect 5742 30046 5794 30098
rect 6862 30046 6914 30098
rect 9550 30046 9602 30098
rect 24894 30046 24946 30098
rect 25230 30046 25282 30098
rect 25454 30046 25506 30098
rect 28142 30046 28194 30098
rect 29598 30046 29650 30098
rect 30270 30046 30322 30098
rect 30382 30046 30434 30098
rect 35758 30046 35810 30098
rect 36094 30046 36146 30098
rect 44158 30046 44210 30098
rect 45838 30046 45890 30098
rect 6638 29934 6690 29986
rect 10670 29934 10722 29986
rect 12462 29934 12514 29986
rect 19518 29934 19570 29986
rect 19630 29934 19682 29986
rect 20078 29934 20130 29986
rect 21422 29934 21474 29986
rect 21534 29934 21586 29986
rect 22430 29934 22482 29986
rect 25678 29934 25730 29986
rect 26462 29934 26514 29986
rect 26910 29934 26962 29986
rect 27694 29934 27746 29986
rect 28254 29934 28306 29986
rect 29486 29934 29538 29986
rect 31278 29934 31330 29986
rect 32958 29934 33010 29986
rect 33406 29934 33458 29986
rect 35646 29934 35698 29986
rect 36430 29934 36482 29986
rect 37214 29934 37266 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 3166 29598 3218 29650
rect 8094 29598 8146 29650
rect 8654 29598 8706 29650
rect 16382 29598 16434 29650
rect 17614 29598 17666 29650
rect 17726 29598 17778 29650
rect 17838 29598 17890 29650
rect 17950 29598 18002 29650
rect 18510 29598 18562 29650
rect 23214 29598 23266 29650
rect 23662 29598 23714 29650
rect 24558 29598 24610 29650
rect 24670 29598 24722 29650
rect 31390 29598 31442 29650
rect 33182 29598 33234 29650
rect 33406 29598 33458 29650
rect 33518 29598 33570 29650
rect 2046 29486 2098 29538
rect 2606 29486 2658 29538
rect 4398 29486 4450 29538
rect 7422 29486 7474 29538
rect 7870 29486 7922 29538
rect 8430 29486 8482 29538
rect 8878 29486 8930 29538
rect 14142 29486 14194 29538
rect 17390 29486 17442 29538
rect 20974 29486 21026 29538
rect 23774 29486 23826 29538
rect 36094 29486 36146 29538
rect 43822 29486 43874 29538
rect 2158 29374 2210 29426
rect 2494 29374 2546 29426
rect 2830 29374 2882 29426
rect 3054 29374 3106 29426
rect 3726 29374 3778 29426
rect 7310 29374 7362 29426
rect 7646 29374 7698 29426
rect 8094 29374 8146 29426
rect 8990 29374 9042 29426
rect 10894 29374 10946 29426
rect 14478 29374 14530 29426
rect 14926 29374 14978 29426
rect 15374 29374 15426 29426
rect 21646 29374 21698 29426
rect 22430 29374 22482 29426
rect 22878 29374 22930 29426
rect 23998 29374 24050 29426
rect 24446 29374 24498 29426
rect 30494 29374 30546 29426
rect 31054 29374 31106 29426
rect 32286 29374 32338 29426
rect 33294 29374 33346 29426
rect 33742 29374 33794 29426
rect 34078 29374 34130 29426
rect 39790 29374 39842 29426
rect 39902 29374 39954 29426
rect 40014 29374 40066 29426
rect 40126 29374 40178 29426
rect 40350 29374 40402 29426
rect 42254 29374 42306 29426
rect 6526 29262 6578 29314
rect 11566 29262 11618 29314
rect 13694 29262 13746 29314
rect 15822 29262 15874 29314
rect 16942 29262 16994 29314
rect 18846 29262 18898 29314
rect 22654 29262 22706 29314
rect 25566 29262 25618 29314
rect 30830 29262 30882 29314
rect 31838 29262 31890 29314
rect 2046 29150 2098 29202
rect 3166 29150 3218 29202
rect 23662 29150 23714 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 6862 28814 6914 28866
rect 25454 28814 25506 28866
rect 26910 28814 26962 28866
rect 1710 28702 1762 28754
rect 6638 28702 6690 28754
rect 7422 28702 7474 28754
rect 11118 28702 11170 28754
rect 13022 28702 13074 28754
rect 20190 28702 20242 28754
rect 21646 28702 21698 28754
rect 22766 28702 22818 28754
rect 24894 28702 24946 28754
rect 25342 28702 25394 28754
rect 28478 28702 28530 28754
rect 29934 28702 29986 28754
rect 32062 28702 32114 28754
rect 33182 28702 33234 28754
rect 35310 28702 35362 28754
rect 36990 28702 37042 28754
rect 40910 28702 40962 28754
rect 41358 28702 41410 28754
rect 44942 28702 44994 28754
rect 45390 28702 45442 28754
rect 4622 28590 4674 28642
rect 6414 28590 6466 28642
rect 6974 28590 7026 28642
rect 9550 28590 9602 28642
rect 10334 28590 10386 28642
rect 10782 28590 10834 28642
rect 11006 28590 11058 28642
rect 11342 28590 11394 28642
rect 12238 28590 12290 28642
rect 19630 28590 19682 28642
rect 20638 28590 20690 28642
rect 21982 28590 22034 28642
rect 26126 28590 26178 28642
rect 26462 28590 26514 28642
rect 26686 28590 26738 28642
rect 27806 28590 27858 28642
rect 28142 28590 28194 28642
rect 29150 28590 29202 28642
rect 32734 28590 32786 28642
rect 35982 28590 36034 28642
rect 39118 28590 39170 28642
rect 39902 28590 39954 28642
rect 40350 28590 40402 28642
rect 41022 28590 41074 28642
rect 43486 28590 43538 28642
rect 44158 28590 44210 28642
rect 44830 28590 44882 28642
rect 45838 28590 45890 28642
rect 3838 28478 3890 28530
rect 5630 28478 5682 28530
rect 11678 28478 11730 28530
rect 16382 28478 16434 28530
rect 25790 28478 25842 28530
rect 32398 28478 32450 28530
rect 40798 28478 40850 28530
rect 5966 28366 6018 28418
rect 6526 28366 6578 28418
rect 11566 28366 11618 28418
rect 11790 28366 11842 28418
rect 13470 28366 13522 28418
rect 13806 28366 13858 28418
rect 20078 28366 20130 28418
rect 20190 28366 20242 28418
rect 20414 28366 20466 28418
rect 26238 28366 26290 28418
rect 27246 28366 27298 28418
rect 32510 28366 32562 28418
rect 40574 28366 40626 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 3838 28030 3890 28082
rect 5742 28030 5794 28082
rect 6302 28030 6354 28082
rect 7198 28030 7250 28082
rect 7422 28030 7474 28082
rect 7758 28030 7810 28082
rect 8318 28030 8370 28082
rect 9662 28030 9714 28082
rect 10446 28030 10498 28082
rect 11790 28030 11842 28082
rect 18846 28030 18898 28082
rect 23214 28030 23266 28082
rect 24558 28030 24610 28082
rect 24670 28030 24722 28082
rect 26798 28030 26850 28082
rect 27246 28030 27298 28082
rect 31614 28030 31666 28082
rect 31950 28030 32002 28082
rect 32062 28030 32114 28082
rect 32286 28030 32338 28082
rect 39566 28030 39618 28082
rect 3166 27918 3218 27970
rect 5294 27918 5346 27970
rect 6414 27918 6466 27970
rect 8766 27918 8818 27970
rect 12126 27918 12178 27970
rect 14702 27918 14754 27970
rect 17838 27918 17890 27970
rect 17950 27918 18002 27970
rect 19518 27918 19570 27970
rect 28254 27918 28306 27970
rect 29710 27918 29762 27970
rect 38334 27918 38386 27970
rect 38894 27918 38946 27970
rect 41246 27918 41298 27970
rect 3054 27806 3106 27858
rect 3502 27806 3554 27858
rect 3950 27806 4002 27858
rect 4174 27806 4226 27858
rect 4622 27806 4674 27858
rect 4958 27806 5010 27858
rect 5182 27806 5234 27858
rect 5518 27806 5570 27858
rect 5854 27806 5906 27858
rect 7086 27806 7138 27858
rect 7646 27806 7698 27858
rect 7982 27806 8034 27858
rect 8094 27806 8146 27858
rect 8542 27806 8594 27858
rect 12462 27806 12514 27858
rect 13246 27806 13298 27858
rect 13358 27806 13410 27858
rect 13582 27806 13634 27858
rect 14030 27806 14082 27858
rect 18398 27806 18450 27858
rect 18622 27806 18674 27858
rect 19070 27806 19122 27858
rect 22654 27806 22706 27858
rect 22990 27806 23042 27858
rect 23326 27806 23378 27858
rect 23662 27806 23714 27858
rect 23998 27806 24050 27858
rect 24446 27806 24498 27858
rect 26126 27806 26178 27858
rect 26350 27806 26402 27858
rect 28702 27806 28754 27858
rect 30942 27806 30994 27858
rect 32510 27806 32562 27858
rect 33182 27806 33234 27858
rect 37326 27806 37378 27858
rect 37662 27806 37714 27858
rect 38782 27806 38834 27858
rect 39454 27806 39506 27858
rect 39790 27806 39842 27858
rect 39902 27806 39954 27858
rect 41022 27806 41074 27858
rect 42142 27806 42194 27858
rect 46062 27806 46114 27858
rect 10334 27694 10386 27746
rect 16830 27694 16882 27746
rect 17502 27694 17554 27746
rect 18734 27694 18786 27746
rect 19854 27694 19906 27746
rect 21982 27694 22034 27746
rect 26014 27694 26066 27746
rect 32174 27694 32226 27746
rect 33854 27694 33906 27746
rect 35982 27694 36034 27746
rect 36430 27694 36482 27746
rect 37774 27694 37826 27746
rect 38110 27694 38162 27746
rect 38334 27694 38386 27746
rect 39678 27694 39730 27746
rect 41918 27694 41970 27746
rect 42702 27694 42754 27746
rect 43262 27694 43314 27746
rect 45390 27694 45442 27746
rect 3166 27582 3218 27634
rect 4734 27582 4786 27634
rect 6302 27582 6354 27634
rect 10222 27582 10274 27634
rect 12798 27582 12850 27634
rect 17390 27582 17442 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 13806 27246 13858 27298
rect 14142 27246 14194 27298
rect 27582 27246 27634 27298
rect 27918 27246 27970 27298
rect 28254 27246 28306 27298
rect 29486 27246 29538 27298
rect 29822 27246 29874 27298
rect 30382 27246 30434 27298
rect 30718 27246 30770 27298
rect 33294 27246 33346 27298
rect 38894 27246 38946 27298
rect 39902 27246 39954 27298
rect 40462 27246 40514 27298
rect 44718 27246 44770 27298
rect 4622 27134 4674 27186
rect 12238 27134 12290 27186
rect 13918 27134 13970 27186
rect 16270 27134 16322 27186
rect 18398 27134 18450 27186
rect 19070 27134 19122 27186
rect 19742 27134 19794 27186
rect 24222 27134 24274 27186
rect 29262 27134 29314 27186
rect 30158 27134 30210 27186
rect 31614 27134 31666 27186
rect 32510 27134 32562 27186
rect 33182 27134 33234 27186
rect 34190 27134 34242 27186
rect 35310 27134 35362 27186
rect 35982 27134 36034 27186
rect 37886 27134 37938 27186
rect 38446 27134 38498 27186
rect 38782 27134 38834 27186
rect 42590 27134 42642 27186
rect 43822 27134 43874 27186
rect 1822 27022 1874 27074
rect 7086 27022 7138 27074
rect 9438 27022 9490 27074
rect 14142 27022 14194 27074
rect 14254 27022 14306 27074
rect 15486 27022 15538 27074
rect 18958 27022 19010 27074
rect 20078 27022 20130 27074
rect 21422 27022 21474 27074
rect 24782 27022 24834 27074
rect 26462 27022 26514 27074
rect 28366 27022 28418 27074
rect 33742 27022 33794 27074
rect 34862 27022 34914 27074
rect 37102 27022 37154 27074
rect 39230 27022 39282 27074
rect 40014 27022 40066 27074
rect 40798 27022 40850 27074
rect 41022 27022 41074 27074
rect 41246 27022 41298 27074
rect 41358 27022 41410 27074
rect 42478 27022 42530 27074
rect 42926 27022 42978 27074
rect 43150 27022 43202 27074
rect 44046 27022 44098 27074
rect 45054 27022 45106 27074
rect 45614 27022 45666 27074
rect 46062 27022 46114 27074
rect 2494 26910 2546 26962
rect 10110 26910 10162 26962
rect 19630 26910 19682 26962
rect 22094 26910 22146 26962
rect 25678 26910 25730 26962
rect 27694 26910 27746 26962
rect 31166 26910 31218 26962
rect 37438 26910 37490 26962
rect 40350 26910 40402 26962
rect 6862 26798 6914 26850
rect 13694 26798 13746 26850
rect 26126 26798 26178 26850
rect 31054 26798 31106 26850
rect 36094 26798 36146 26850
rect 39566 26798 39618 26850
rect 41134 26798 41186 26850
rect 41806 26854 41858 26906
rect 41918 26910 41970 26962
rect 42702 26910 42754 26962
rect 44830 26910 44882 26962
rect 45278 26910 45330 26962
rect 42142 26798 42194 26850
rect 43486 26798 43538 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 3166 26462 3218 26514
rect 3950 26462 4002 26514
rect 4622 26462 4674 26514
rect 10334 26462 10386 26514
rect 17614 26462 17666 26514
rect 22990 26462 23042 26514
rect 24110 26462 24162 26514
rect 24782 26462 24834 26514
rect 28478 26462 28530 26514
rect 37774 26462 37826 26514
rect 38446 26462 38498 26514
rect 39902 26462 39954 26514
rect 40350 26462 40402 26514
rect 3054 26350 3106 26402
rect 3838 26350 3890 26402
rect 4398 26350 4450 26402
rect 9886 26350 9938 26402
rect 17950 26350 18002 26402
rect 21198 26350 21250 26402
rect 23662 26350 23714 26402
rect 26238 26350 26290 26402
rect 30270 26350 30322 26402
rect 39454 26350 39506 26402
rect 42254 26350 42306 26402
rect 3726 26238 3778 26290
rect 4286 26238 4338 26290
rect 4734 26238 4786 26290
rect 5742 26238 5794 26290
rect 9662 26238 9714 26290
rect 10782 26238 10834 26290
rect 13918 26238 13970 26290
rect 18286 26238 18338 26290
rect 19630 26238 19682 26290
rect 21758 26238 21810 26290
rect 22878 26238 22930 26290
rect 23102 26238 23154 26290
rect 23550 26238 23602 26290
rect 25454 26238 25506 26290
rect 29598 26238 29650 26290
rect 33406 26238 33458 26290
rect 36878 26238 36930 26290
rect 37326 26238 37378 26290
rect 37550 26238 37602 26290
rect 37998 26238 38050 26290
rect 38782 26238 38834 26290
rect 45502 26238 45554 26290
rect 6414 26126 6466 26178
rect 8542 26126 8594 26178
rect 11454 26126 11506 26178
rect 13582 26126 13634 26178
rect 14702 26126 14754 26178
rect 16830 26126 16882 26178
rect 20526 26126 20578 26178
rect 22654 26126 22706 26178
rect 32398 26126 32450 26178
rect 34190 26126 34242 26178
rect 36318 26126 36370 26178
rect 36766 26126 36818 26178
rect 37662 26126 37714 26178
rect 40238 26126 40290 26178
rect 3166 26014 3218 26066
rect 22430 26014 22482 26066
rect 39342 26014 39394 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6414 25678 6466 25730
rect 21422 25678 21474 25730
rect 29486 25678 29538 25730
rect 35982 25678 36034 25730
rect 36318 25678 36370 25730
rect 37326 25678 37378 25730
rect 44830 25678 44882 25730
rect 45166 25678 45218 25730
rect 1710 25566 1762 25618
rect 12798 25566 12850 25618
rect 17502 25566 17554 25618
rect 19294 25566 19346 25618
rect 20414 25566 20466 25618
rect 21310 25566 21362 25618
rect 24670 25566 24722 25618
rect 29710 25566 29762 25618
rect 30718 25566 30770 25618
rect 31166 25566 31218 25618
rect 32174 25566 32226 25618
rect 33182 25566 33234 25618
rect 35310 25566 35362 25618
rect 37102 25566 37154 25618
rect 40798 25566 40850 25618
rect 45614 25566 45666 25618
rect 46174 25566 46226 25618
rect 4510 25454 4562 25506
rect 5854 25454 5906 25506
rect 8318 25454 8370 25506
rect 13582 25454 13634 25506
rect 18062 25454 18114 25506
rect 18398 25454 18450 25506
rect 18510 25454 18562 25506
rect 18734 25454 18786 25506
rect 18958 25454 19010 25506
rect 19406 25454 19458 25506
rect 19854 25454 19906 25506
rect 20078 25454 20130 25506
rect 20302 25454 20354 25506
rect 21870 25454 21922 25506
rect 25118 25454 25170 25506
rect 25230 25454 25282 25506
rect 26238 25454 26290 25506
rect 31278 25454 31330 25506
rect 31502 25454 31554 25506
rect 32062 25454 32114 25506
rect 32510 25454 32562 25506
rect 32734 25454 32786 25506
rect 35758 25454 35810 25506
rect 36206 25454 36258 25506
rect 38558 25454 38610 25506
rect 38894 25454 38946 25506
rect 39230 25454 39282 25506
rect 39678 25454 39730 25506
rect 41470 25454 41522 25506
rect 41582 25454 41634 25506
rect 41694 25454 41746 25506
rect 42030 25454 42082 25506
rect 43262 25454 43314 25506
rect 44270 25454 44322 25506
rect 46062 25454 46114 25506
rect 3838 25342 3890 25394
rect 5630 25342 5682 25394
rect 6750 25342 6802 25394
rect 11006 25342 11058 25394
rect 14254 25342 14306 25394
rect 22542 25342 22594 25394
rect 25454 25342 25506 25394
rect 25566 25342 25618 25394
rect 26014 25342 26066 25394
rect 26798 25342 26850 25394
rect 27134 25342 27186 25394
rect 30606 25342 30658 25394
rect 31166 25342 31218 25394
rect 31726 25342 31778 25394
rect 35422 25342 35474 25394
rect 40126 25342 40178 25394
rect 40350 25342 40402 25394
rect 42814 25342 42866 25394
rect 6526 25230 6578 25282
rect 16494 25230 16546 25282
rect 18622 25230 18674 25282
rect 20526 25230 20578 25282
rect 25342 25230 25394 25282
rect 27246 25230 27298 25282
rect 29150 25230 29202 25282
rect 32286 25230 32338 25282
rect 33630 25230 33682 25282
rect 35198 25230 35250 25282
rect 37662 25230 37714 25282
rect 38334 25230 38386 25282
rect 38894 25230 38946 25282
rect 39902 25230 39954 25282
rect 40686 25230 40738 25282
rect 42366 25230 42418 25282
rect 43150 25230 43202 25282
rect 44158 25230 44210 25282
rect 45054 25230 45106 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 3278 24894 3330 24946
rect 3838 24894 3890 24946
rect 5406 24894 5458 24946
rect 7198 24894 7250 24946
rect 7310 24894 7362 24946
rect 7422 24894 7474 24946
rect 9774 24894 9826 24946
rect 23998 24894 24050 24946
rect 25230 24894 25282 24946
rect 37550 24894 37602 24946
rect 38222 24894 38274 24946
rect 4622 24782 4674 24834
rect 5518 24782 5570 24834
rect 6526 24782 6578 24834
rect 7982 24782 8034 24834
rect 8094 24782 8146 24834
rect 8542 24782 8594 24834
rect 8654 24782 8706 24834
rect 16830 24782 16882 24834
rect 23326 24782 23378 24834
rect 24110 24782 24162 24834
rect 28366 24782 28418 24834
rect 30382 24782 30434 24834
rect 34862 24782 34914 24834
rect 36766 24782 36818 24834
rect 36990 24782 37042 24834
rect 39902 24782 39954 24834
rect 40014 24782 40066 24834
rect 41022 24782 41074 24834
rect 41134 24782 41186 24834
rect 41470 24782 41522 24834
rect 3166 24670 3218 24722
rect 3502 24670 3554 24722
rect 3726 24670 3778 24722
rect 3950 24670 4002 24722
rect 4174 24670 4226 24722
rect 4958 24670 5010 24722
rect 6190 24670 6242 24722
rect 6750 24670 6802 24722
rect 8318 24670 8370 24722
rect 8878 24670 8930 24722
rect 9438 24670 9490 24722
rect 9774 24670 9826 24722
rect 10110 24670 10162 24722
rect 11006 24670 11058 24722
rect 14478 24670 14530 24722
rect 14814 24670 14866 24722
rect 15038 24670 15090 24722
rect 16382 24670 16434 24722
rect 17726 24670 17778 24722
rect 23662 24670 23714 24722
rect 25566 24670 25618 24722
rect 29150 24670 29202 24722
rect 29710 24670 29762 24722
rect 35422 24670 35474 24722
rect 36654 24670 36706 24722
rect 37102 24670 37154 24722
rect 37662 24670 37714 24722
rect 38110 24670 38162 24722
rect 38334 24670 38386 24722
rect 39454 24670 39506 24722
rect 40238 24670 40290 24722
rect 41582 24670 41634 24722
rect 42254 24670 42306 24722
rect 43374 24670 43426 24722
rect 11790 24558 11842 24610
rect 13918 24558 13970 24610
rect 14702 24558 14754 24610
rect 22318 24558 22370 24610
rect 24558 24558 24610 24610
rect 26238 24558 26290 24610
rect 32510 24558 32562 24610
rect 34190 24558 34242 24610
rect 34974 24558 35026 24610
rect 39006 24558 39058 24610
rect 42478 24558 42530 24610
rect 42926 24558 42978 24610
rect 44046 24558 44098 24610
rect 46174 24558 46226 24610
rect 5406 24446 5458 24498
rect 16718 24446 16770 24498
rect 24446 24446 24498 24498
rect 34302 24446 34354 24498
rect 34638 24446 34690 24498
rect 35534 24446 35586 24498
rect 35758 24446 35810 24498
rect 35870 24446 35922 24498
rect 39230 24446 39282 24498
rect 41022 24446 41074 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12350 24110 12402 24162
rect 12686 24110 12738 24162
rect 29486 24110 29538 24162
rect 30270 24110 30322 24162
rect 40350 24110 40402 24162
rect 43374 24110 43426 24162
rect 43710 24110 43762 24162
rect 44830 24110 44882 24162
rect 46062 24110 46114 24162
rect 7198 23998 7250 24050
rect 7646 23998 7698 24050
rect 7758 23998 7810 24050
rect 8654 23998 8706 24050
rect 13918 23998 13970 24050
rect 14702 23998 14754 24050
rect 14814 23998 14866 24050
rect 16382 23998 16434 24050
rect 18510 23998 18562 24050
rect 30046 23998 30098 24050
rect 31838 23998 31890 24050
rect 33966 23998 34018 24050
rect 34414 23998 34466 24050
rect 39566 23998 39618 24050
rect 40462 23998 40514 24050
rect 40910 23998 40962 24050
rect 41470 23998 41522 24050
rect 42478 23998 42530 24050
rect 45166 23998 45218 24050
rect 45838 23998 45890 24050
rect 46174 23998 46226 24050
rect 3838 23886 3890 23938
rect 4062 23886 4114 23938
rect 6862 23886 6914 23938
rect 7086 23886 7138 23938
rect 7982 23886 8034 23938
rect 11454 23886 11506 23938
rect 12462 23886 12514 23938
rect 12910 23886 12962 23938
rect 13806 23886 13858 23938
rect 15710 23886 15762 23938
rect 19182 23886 19234 23938
rect 19406 23886 19458 23938
rect 19630 23886 19682 23938
rect 19854 23886 19906 23938
rect 20078 23886 20130 23938
rect 20302 23886 20354 23938
rect 21198 23886 21250 23938
rect 21534 23886 21586 23938
rect 22206 23886 22258 23938
rect 23550 23886 23602 23938
rect 29710 23886 29762 23938
rect 31166 23886 31218 23938
rect 34638 23886 34690 23938
rect 35310 23886 35362 23938
rect 35646 23886 35698 23938
rect 36206 23886 36258 23938
rect 37214 23886 37266 23938
rect 37550 23886 37602 23938
rect 37886 23886 37938 23938
rect 39454 23886 39506 23938
rect 39678 23886 39730 23938
rect 40126 23886 40178 23938
rect 42254 23886 42306 23938
rect 42366 23886 42418 23938
rect 42814 23886 42866 23938
rect 43150 23886 43202 23938
rect 43598 23886 43650 23938
rect 3502 23774 3554 23826
rect 6078 23774 6130 23826
rect 6414 23774 6466 23826
rect 7310 23774 7362 23826
rect 10782 23774 10834 23826
rect 12014 23774 12066 23826
rect 19070 23774 19122 23826
rect 22430 23774 22482 23826
rect 22542 23774 22594 23826
rect 25342 23774 25394 23826
rect 36094 23774 36146 23826
rect 36318 23774 36370 23826
rect 36990 23774 37042 23826
rect 38334 23774 38386 23826
rect 44158 23774 44210 23826
rect 45054 23774 45106 23826
rect 3614 23662 3666 23714
rect 4398 23662 4450 23714
rect 4734 23662 4786 23714
rect 5742 23662 5794 23714
rect 14030 23662 14082 23714
rect 14254 23662 14306 23714
rect 14926 23662 14978 23714
rect 20414 23662 20466 23714
rect 20526 23662 20578 23714
rect 21422 23662 21474 23714
rect 22094 23662 22146 23714
rect 22990 23662 23042 23714
rect 29150 23662 29202 23714
rect 30606 23662 30658 23714
rect 37438 23662 37490 23714
rect 37998 23662 38050 23714
rect 38110 23662 38162 23714
rect 41806 23662 41858 23714
rect 42590 23662 42642 23714
rect 44046 23662 44098 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 4958 23326 5010 23378
rect 5518 23326 5570 23378
rect 8990 23326 9042 23378
rect 9774 23326 9826 23378
rect 13582 23326 13634 23378
rect 22542 23326 22594 23378
rect 25790 23326 25842 23378
rect 25902 23326 25954 23378
rect 26126 23326 26178 23378
rect 27358 23326 27410 23378
rect 27470 23326 27522 23378
rect 27582 23326 27634 23378
rect 28142 23326 28194 23378
rect 28702 23326 28754 23378
rect 35646 23326 35698 23378
rect 36878 23326 36930 23378
rect 40350 23326 40402 23378
rect 41358 23326 41410 23378
rect 2494 23214 2546 23266
rect 5742 23214 5794 23266
rect 7646 23214 7698 23266
rect 8654 23214 8706 23266
rect 8766 23214 8818 23266
rect 10558 23214 10610 23266
rect 14702 23214 14754 23266
rect 17950 23214 18002 23266
rect 20190 23214 20242 23266
rect 22990 23214 23042 23266
rect 23102 23214 23154 23266
rect 24222 23214 24274 23266
rect 26014 23214 26066 23266
rect 26686 23214 26738 23266
rect 33742 23214 33794 23266
rect 39118 23214 39170 23266
rect 40238 23214 40290 23266
rect 41582 23214 41634 23266
rect 42254 23214 42306 23266
rect 42366 23214 42418 23266
rect 42478 23214 42530 23266
rect 45390 23214 45442 23266
rect 1822 23102 1874 23154
rect 5294 23102 5346 23154
rect 5854 23102 5906 23154
rect 6414 23102 6466 23154
rect 6638 23102 6690 23154
rect 6862 23102 6914 23154
rect 7198 23102 7250 23154
rect 7534 23102 7586 23154
rect 7758 23102 7810 23154
rect 8206 23102 8258 23154
rect 9438 23102 9490 23154
rect 9886 23102 9938 23154
rect 10110 23102 10162 23154
rect 10334 23102 10386 23154
rect 10670 23102 10722 23154
rect 13022 23102 13074 23154
rect 13246 23102 13298 23154
rect 14030 23102 14082 23154
rect 18286 23102 18338 23154
rect 19630 23102 19682 23154
rect 20638 23102 20690 23154
rect 21758 23102 21810 23154
rect 22654 23102 22706 23154
rect 23662 23102 23714 23154
rect 23998 23102 24050 23154
rect 24334 23102 24386 23154
rect 25566 23102 25618 23154
rect 27022 23102 27074 23154
rect 27246 23102 27298 23154
rect 29486 23102 29538 23154
rect 29710 23102 29762 23154
rect 30494 23102 30546 23154
rect 31166 23102 31218 23154
rect 31614 23102 31666 23154
rect 31838 23102 31890 23154
rect 32398 23102 32450 23154
rect 33518 23102 33570 23154
rect 34190 23102 34242 23154
rect 34638 23102 34690 23154
rect 35422 23102 35474 23154
rect 35758 23102 35810 23154
rect 35870 23102 35922 23154
rect 38222 23102 38274 23154
rect 38558 23102 38610 23154
rect 39006 23102 39058 23154
rect 39230 23102 39282 23154
rect 39454 23102 39506 23154
rect 41022 23102 41074 23154
rect 41134 23102 41186 23154
rect 41246 23102 41298 23154
rect 46062 23102 46114 23154
rect 4622 22990 4674 23042
rect 16830 22990 16882 23042
rect 17726 22990 17778 23042
rect 26574 22990 26626 23042
rect 29150 22990 29202 23042
rect 30830 22990 30882 23042
rect 31726 22990 31778 23042
rect 35086 22990 35138 23042
rect 36094 22990 36146 23042
rect 36430 22990 36482 23042
rect 43262 22990 43314 23042
rect 7086 22878 7138 22930
rect 8094 22878 8146 22930
rect 22542 22878 22594 22930
rect 23102 22878 23154 22930
rect 23774 22878 23826 22930
rect 30046 22878 30098 22930
rect 36430 22878 36482 22930
rect 38110 22878 38162 22930
rect 38446 22878 38498 22930
rect 39902 22878 39954 22930
rect 42926 22878 42978 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19630 22542 19682 22594
rect 21310 22542 21362 22594
rect 21534 22542 21586 22594
rect 27246 22542 27298 22594
rect 27582 22542 27634 22594
rect 41022 22542 41074 22594
rect 42366 22542 42418 22594
rect 43822 22542 43874 22594
rect 4734 22430 4786 22482
rect 6750 22430 6802 22482
rect 12910 22430 12962 22482
rect 17950 22430 18002 22482
rect 18510 22430 18562 22482
rect 19294 22430 19346 22482
rect 23102 22430 23154 22482
rect 25230 22430 25282 22482
rect 26798 22430 26850 22482
rect 39230 22430 39282 22482
rect 43150 22430 43202 22482
rect 43710 22430 43762 22482
rect 45054 22430 45106 22482
rect 45614 22430 45666 22482
rect 4062 22318 4114 22370
rect 4398 22318 4450 22370
rect 9662 22318 9714 22370
rect 9998 22318 10050 22370
rect 13694 22318 13746 22370
rect 15710 22318 15762 22370
rect 18622 22318 18674 22370
rect 19742 22318 19794 22370
rect 21870 22318 21922 22370
rect 22318 22318 22370 22370
rect 25790 22318 25842 22370
rect 28030 22318 28082 22370
rect 29374 22318 29426 22370
rect 30046 22318 30098 22370
rect 35982 22318 36034 22370
rect 37662 22318 37714 22370
rect 39342 22318 39394 22370
rect 40014 22318 40066 22370
rect 42702 22318 42754 22370
rect 43038 22318 43090 22370
rect 44046 22318 44098 22370
rect 3390 22206 3442 22258
rect 4958 22206 5010 22258
rect 5742 22206 5794 22258
rect 5854 22206 5906 22258
rect 8878 22206 8930 22258
rect 10782 22206 10834 22258
rect 14814 22206 14866 22258
rect 16270 22206 16322 22258
rect 20414 22206 20466 22258
rect 25678 22206 25730 22258
rect 27358 22206 27410 22258
rect 29150 22206 29202 22258
rect 29598 22206 29650 22258
rect 33854 22206 33906 22258
rect 37326 22206 37378 22258
rect 37998 22206 38050 22258
rect 39566 22206 39618 22258
rect 40910 22206 40962 22258
rect 41806 22206 41858 22258
rect 43262 22206 43314 22258
rect 44158 22206 44210 22258
rect 45838 22206 45890 22258
rect 46174 22206 46226 22258
rect 5518 22094 5570 22146
rect 6302 22094 6354 22146
rect 13806 22094 13858 22146
rect 20526 22094 20578 22146
rect 21534 22094 21586 22146
rect 21982 22094 22034 22146
rect 25454 22094 25506 22146
rect 26350 22094 26402 22146
rect 28590 22094 28642 22146
rect 29038 22094 29090 22146
rect 35982 22094 36034 22146
rect 36206 22094 36258 22146
rect 36430 22094 36482 22146
rect 36990 22094 37042 22146
rect 38894 22094 38946 22146
rect 42142 22094 42194 22146
rect 42254 22094 42306 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 5966 21758 6018 21810
rect 6974 21758 7026 21810
rect 7870 21758 7922 21810
rect 8430 21758 8482 21810
rect 9662 21758 9714 21810
rect 14142 21758 14194 21810
rect 15934 21758 15986 21810
rect 17726 21758 17778 21810
rect 23214 21758 23266 21810
rect 24334 21758 24386 21810
rect 26126 21758 26178 21810
rect 29710 21758 29762 21810
rect 32062 21758 32114 21810
rect 33742 21758 33794 21810
rect 37774 21758 37826 21810
rect 38894 21758 38946 21810
rect 39678 21758 39730 21810
rect 39790 21758 39842 21810
rect 39902 21758 39954 21810
rect 40238 21758 40290 21810
rect 4958 21646 5010 21698
rect 5854 21646 5906 21698
rect 7086 21646 7138 21698
rect 7758 21646 7810 21698
rect 8318 21646 8370 21698
rect 10110 21646 10162 21698
rect 13358 21646 13410 21698
rect 13918 21646 13970 21698
rect 17390 21646 17442 21698
rect 18846 21646 18898 21698
rect 22990 21646 23042 21698
rect 24110 21646 24162 21698
rect 25230 21646 25282 21698
rect 28702 21646 28754 21698
rect 32398 21646 32450 21698
rect 35310 21646 35362 21698
rect 38110 21646 38162 21698
rect 45390 21646 45442 21698
rect 1822 21534 1874 21586
rect 5294 21534 5346 21586
rect 6190 21534 6242 21586
rect 6750 21534 6802 21586
rect 8094 21534 8146 21586
rect 8654 21534 8706 21586
rect 9438 21534 9490 21586
rect 9774 21534 9826 21586
rect 14478 21534 14530 21586
rect 14814 21534 14866 21586
rect 15038 21534 15090 21586
rect 16718 21534 16770 21586
rect 18398 21534 18450 21586
rect 22094 21534 22146 21586
rect 22542 21534 22594 21586
rect 22878 21534 22930 21586
rect 23998 21534 24050 21586
rect 25566 21534 25618 21586
rect 29486 21534 29538 21586
rect 30158 21534 30210 21586
rect 31166 21534 31218 21586
rect 31502 21534 31554 21586
rect 34526 21534 34578 21586
rect 38558 21534 38610 21586
rect 39230 21534 39282 21586
rect 42366 21534 42418 21586
rect 46062 21534 46114 21586
rect 2494 21422 2546 21474
rect 4622 21422 4674 21474
rect 13246 21422 13298 21474
rect 14030 21422 14082 21474
rect 16382 21422 16434 21474
rect 19182 21422 19234 21474
rect 21310 21422 21362 21474
rect 23102 21422 23154 21474
rect 24222 21422 24274 21474
rect 25342 21422 25394 21474
rect 26238 21422 26290 21474
rect 26574 21422 26626 21474
rect 30606 21422 30658 21474
rect 31726 21422 31778 21474
rect 33182 21422 33234 21474
rect 37438 21422 37490 21474
rect 39006 21422 39058 21474
rect 40350 21422 40402 21474
rect 41806 21422 41858 21474
rect 42142 21422 42194 21474
rect 43262 21422 43314 21474
rect 13582 21310 13634 21362
rect 15374 21310 15426 21362
rect 18734 21310 18786 21362
rect 23662 21310 23714 21362
rect 30382 21310 30434 21362
rect 33070 21310 33122 21362
rect 41246 21310 41298 21362
rect 41582 21310 41634 21362
rect 42702 21310 42754 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 20526 20974 20578 21026
rect 20862 20974 20914 21026
rect 21310 20974 21362 21026
rect 35310 20974 35362 21026
rect 35646 20974 35698 21026
rect 35870 20974 35922 21026
rect 36430 20974 36482 21026
rect 44942 20974 44994 21026
rect 45166 20974 45218 21026
rect 45278 20974 45330 21026
rect 8766 20862 8818 20914
rect 10894 20862 10946 20914
rect 12910 20862 12962 20914
rect 18174 20862 18226 20914
rect 21534 20862 21586 20914
rect 21870 20862 21922 20914
rect 29598 20862 29650 20914
rect 34190 20862 34242 20914
rect 35086 20862 35138 20914
rect 36206 20862 36258 20914
rect 39566 20862 39618 20914
rect 40350 20862 40402 20914
rect 41022 20862 41074 20914
rect 41358 20862 41410 20914
rect 45950 20862 46002 20914
rect 2382 20750 2434 20802
rect 2718 20750 2770 20802
rect 3950 20750 4002 20802
rect 4622 20750 4674 20802
rect 5966 20750 6018 20802
rect 12686 20750 12738 20802
rect 14030 20750 14082 20802
rect 14254 20750 14306 20802
rect 15262 20750 15314 20802
rect 19070 20750 19122 20802
rect 19182 20750 19234 20802
rect 19854 20750 19906 20802
rect 21758 20750 21810 20802
rect 21982 20750 22034 20802
rect 22542 20750 22594 20802
rect 23998 20750 24050 20802
rect 25006 20750 25058 20802
rect 26350 20750 26402 20802
rect 27022 20750 27074 20802
rect 29038 20750 29090 20802
rect 29710 20750 29762 20802
rect 31390 20750 31442 20802
rect 32062 20750 32114 20802
rect 37326 20750 37378 20802
rect 37774 20750 37826 20802
rect 39678 20750 39730 20802
rect 44270 20750 44322 20802
rect 2830 20638 2882 20690
rect 3054 20638 3106 20690
rect 3278 20638 3330 20690
rect 3502 20638 3554 20690
rect 4174 20638 4226 20690
rect 4510 20638 4562 20690
rect 6638 20638 6690 20690
rect 9438 20638 9490 20690
rect 11230 20638 11282 20690
rect 16046 20638 16098 20690
rect 18958 20638 19010 20690
rect 25790 20638 25842 20690
rect 27246 20638 27298 20690
rect 27358 20638 27410 20690
rect 30718 20638 30770 20690
rect 36990 20638 37042 20690
rect 37998 20638 38050 20690
rect 38782 20638 38834 20690
rect 39902 20638 39954 20690
rect 40686 20638 40738 20690
rect 40910 20638 40962 20690
rect 43486 20638 43538 20690
rect 44830 20638 44882 20690
rect 2046 20526 2098 20578
rect 2270 20526 2322 20578
rect 3614 20526 3666 20578
rect 4286 20526 4338 20578
rect 9102 20526 9154 20578
rect 11006 20526 11058 20578
rect 11790 20526 11842 20578
rect 12350 20526 12402 20578
rect 14142 20526 14194 20578
rect 14478 20526 14530 20578
rect 18510 20526 18562 20578
rect 20302 20526 20354 20578
rect 20750 20526 20802 20578
rect 22766 20526 22818 20578
rect 27806 20526 27858 20578
rect 28142 20526 28194 20578
rect 28478 20526 28530 20578
rect 29486 20526 29538 20578
rect 30046 20526 30098 20578
rect 30382 20526 30434 20578
rect 30830 20526 30882 20578
rect 34750 20526 34802 20578
rect 38558 20526 38610 20578
rect 38894 20526 38946 20578
rect 39342 20526 39394 20578
rect 39454 20526 39506 20578
rect 40238 20526 40290 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 17614 20190 17666 20242
rect 23662 20190 23714 20242
rect 27806 20190 27858 20242
rect 30046 20190 30098 20242
rect 30718 20190 30770 20242
rect 31726 20190 31778 20242
rect 33406 20190 33458 20242
rect 38894 20190 38946 20242
rect 2046 20078 2098 20130
rect 2270 20078 2322 20130
rect 8542 20078 8594 20130
rect 8878 20078 8930 20130
rect 15262 20078 15314 20130
rect 17838 20078 17890 20130
rect 18174 20078 18226 20130
rect 19294 20078 19346 20130
rect 20078 20078 20130 20130
rect 21198 20078 21250 20130
rect 24334 20078 24386 20130
rect 27358 20078 27410 20130
rect 34190 20078 34242 20130
rect 36094 20078 36146 20130
rect 38446 20078 38498 20130
rect 39006 20078 39058 20130
rect 39118 20078 39170 20130
rect 2606 19966 2658 20018
rect 8206 19966 8258 20018
rect 13022 19966 13074 20018
rect 18286 19966 18338 20018
rect 20526 19966 20578 20018
rect 23774 19966 23826 20018
rect 26462 19966 26514 20018
rect 26686 19966 26738 20018
rect 26798 19966 26850 20018
rect 27022 19966 27074 20018
rect 27582 19966 27634 20018
rect 33070 19966 33122 20018
rect 33294 19966 33346 20018
rect 33518 19966 33570 20018
rect 33630 19966 33682 20018
rect 34302 19966 34354 20018
rect 34526 19966 34578 20018
rect 34750 19966 34802 20018
rect 38782 19966 38834 20018
rect 39566 19966 39618 20018
rect 40014 19966 40066 20018
rect 40238 19966 40290 20018
rect 40910 19966 40962 20018
rect 2494 19854 2546 19906
rect 3390 19854 3442 19906
rect 9774 19854 9826 19906
rect 17950 19854 18002 19906
rect 18846 19854 18898 19906
rect 23326 19854 23378 19906
rect 24670 19854 24722 19906
rect 26014 19854 26066 19906
rect 27694 19854 27746 19906
rect 28254 19854 28306 19906
rect 28702 19854 28754 19906
rect 29150 19854 29202 19906
rect 29598 19854 29650 19906
rect 31278 19854 31330 19906
rect 34414 19854 34466 19906
rect 35086 19854 35138 19906
rect 35646 19854 35698 19906
rect 36654 19854 36706 19906
rect 37102 19854 37154 19906
rect 37550 19854 37602 19906
rect 37886 19854 37938 19906
rect 44718 19854 44770 19906
rect 31166 19742 31218 19794
rect 35198 19742 35250 19794
rect 35534 19742 35586 19794
rect 38222 19742 38274 19794
rect 39902 19742 39954 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 8094 19406 8146 19458
rect 8542 19406 8594 19458
rect 16158 19406 16210 19458
rect 16270 19406 16322 19458
rect 16494 19406 16546 19458
rect 2494 19294 2546 19346
rect 4622 19294 4674 19346
rect 6638 19294 6690 19346
rect 12910 19294 12962 19346
rect 13806 19294 13858 19346
rect 18174 19294 18226 19346
rect 21534 19294 21586 19346
rect 22430 19294 22482 19346
rect 29598 19406 29650 19458
rect 45278 19406 45330 19458
rect 45726 19406 45778 19458
rect 23102 19294 23154 19346
rect 25342 19294 25394 19346
rect 29038 19294 29090 19346
rect 30718 19294 30770 19346
rect 32846 19294 32898 19346
rect 33518 19294 33570 19346
rect 35646 19294 35698 19346
rect 38670 19294 38722 19346
rect 39678 19294 39730 19346
rect 41022 19294 41074 19346
rect 41358 19294 41410 19346
rect 1822 19182 1874 19234
rect 5518 19182 5570 19234
rect 6190 19182 6242 19234
rect 6414 19182 6466 19234
rect 6750 19182 6802 19234
rect 7534 19182 7586 19234
rect 7758 19182 7810 19234
rect 8654 19182 8706 19234
rect 10110 19182 10162 19234
rect 13582 19182 13634 19234
rect 14478 19182 14530 19234
rect 15038 19182 15090 19234
rect 15262 19182 15314 19234
rect 16718 19182 16770 19234
rect 17054 19182 17106 19234
rect 17390 19182 17442 19234
rect 17838 19182 17890 19234
rect 19518 19182 19570 19234
rect 21982 19182 22034 19234
rect 24670 19182 24722 19234
rect 29934 19182 29986 19234
rect 36430 19182 36482 19234
rect 39006 19182 39058 19234
rect 40462 19182 40514 19234
rect 40798 19182 40850 19234
rect 44270 19182 44322 19234
rect 44942 19182 44994 19234
rect 45166 19182 45218 19234
rect 45838 19182 45890 19234
rect 5742 19070 5794 19122
rect 5854 19070 5906 19122
rect 10782 19070 10834 19122
rect 17166 19070 17218 19122
rect 19966 19070 20018 19122
rect 20414 19070 20466 19122
rect 37214 19070 37266 19122
rect 39230 19070 39282 19122
rect 43486 19070 43538 19122
rect 44830 19070 44882 19122
rect 45950 19070 46002 19122
rect 7198 18958 7250 19010
rect 8542 18958 8594 19010
rect 9102 18958 9154 19010
rect 15598 18958 15650 19010
rect 20750 18958 20802 19010
rect 21422 18958 21474 19010
rect 29262 18958 29314 19010
rect 36878 18958 36930 19010
rect 37102 18958 37154 19010
rect 37886 18958 37938 19010
rect 38222 18958 38274 19010
rect 38670 18958 38722 19010
rect 38782 18958 38834 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 8654 18622 8706 18674
rect 11006 18622 11058 18674
rect 12014 18622 12066 18674
rect 17726 18622 17778 18674
rect 31726 18622 31778 18674
rect 31838 18622 31890 18674
rect 39790 18622 39842 18674
rect 17390 18510 17442 18562
rect 18286 18510 18338 18562
rect 19406 18510 19458 18562
rect 20190 18510 20242 18562
rect 25230 18510 25282 18562
rect 30046 18510 30098 18562
rect 32062 18510 32114 18562
rect 38894 18510 38946 18562
rect 39566 18510 39618 18562
rect 44158 18510 44210 18562
rect 44942 18510 44994 18562
rect 45166 18510 45218 18562
rect 45278 18510 45330 18562
rect 1822 18398 1874 18450
rect 2494 18398 2546 18450
rect 5294 18398 5346 18450
rect 6078 18398 6130 18450
rect 12238 18398 12290 18450
rect 15374 18398 15426 18450
rect 16606 18398 16658 18450
rect 18622 18398 18674 18450
rect 19070 18398 19122 18450
rect 19966 18398 20018 18450
rect 20414 18398 20466 18450
rect 20526 18398 20578 18450
rect 21310 18398 21362 18450
rect 21534 18398 21586 18450
rect 21758 18398 21810 18450
rect 22094 18398 22146 18450
rect 22430 18398 22482 18450
rect 23326 18398 23378 18450
rect 24334 18398 24386 18450
rect 25454 18398 25506 18450
rect 26350 18398 26402 18450
rect 29598 18398 29650 18450
rect 29822 18398 29874 18450
rect 30158 18398 30210 18450
rect 31502 18398 31554 18450
rect 31614 18398 31666 18450
rect 32510 18398 32562 18450
rect 33518 18398 33570 18450
rect 33854 18398 33906 18450
rect 40910 18398 40962 18450
rect 41694 18398 41746 18450
rect 44382 18398 44434 18450
rect 44830 18398 44882 18450
rect 4622 18286 4674 18338
rect 8206 18286 8258 18338
rect 8542 18286 8594 18338
rect 11118 18286 11170 18338
rect 11902 18286 11954 18338
rect 12574 18286 12626 18338
rect 14702 18286 14754 18338
rect 15934 18286 15986 18338
rect 16830 18286 16882 18338
rect 18734 18286 18786 18338
rect 20302 18286 20354 18338
rect 21646 18286 21698 18338
rect 22990 18286 23042 18338
rect 23886 18286 23938 18338
rect 27134 18286 27186 18338
rect 29262 18286 29314 18338
rect 29934 18286 29986 18338
rect 30718 18286 30770 18338
rect 39902 18286 39954 18338
rect 40238 18286 40290 18338
rect 43822 18286 43874 18338
rect 44606 18286 44658 18338
rect 45726 18286 45778 18338
rect 46174 18286 46226 18338
rect 11230 18174 11282 18226
rect 16270 18174 16322 18226
rect 40350 18174 40402 18226
rect 45614 18174 45666 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 20414 17838 20466 17890
rect 27806 17838 27858 17890
rect 29150 17838 29202 17890
rect 31726 17838 31778 17890
rect 42590 17838 42642 17890
rect 6526 17726 6578 17778
rect 10782 17726 10834 17778
rect 12910 17726 12962 17778
rect 19854 17726 19906 17778
rect 20750 17726 20802 17778
rect 22206 17726 22258 17778
rect 24558 17726 24610 17778
rect 26686 17726 26738 17778
rect 27918 17726 27970 17778
rect 29486 17726 29538 17778
rect 31390 17726 31442 17778
rect 32062 17726 32114 17778
rect 33406 17726 33458 17778
rect 42702 17726 42754 17778
rect 43374 17726 43426 17778
rect 44942 17726 44994 17778
rect 45390 17726 45442 17778
rect 2718 17614 2770 17666
rect 3054 17614 3106 17666
rect 3838 17614 3890 17666
rect 4174 17614 4226 17666
rect 6078 17614 6130 17666
rect 10110 17614 10162 17666
rect 13918 17614 13970 17666
rect 14254 17614 14306 17666
rect 14478 17614 14530 17666
rect 16046 17614 16098 17666
rect 22318 17614 22370 17666
rect 22766 17614 22818 17666
rect 23102 17614 23154 17666
rect 23774 17614 23826 17666
rect 29822 17614 29874 17666
rect 30830 17614 30882 17666
rect 32398 17614 32450 17666
rect 32846 17614 32898 17666
rect 33294 17614 33346 17666
rect 33742 17614 33794 17666
rect 33966 17614 34018 17666
rect 34526 17614 34578 17666
rect 36318 17614 36370 17666
rect 40798 17614 40850 17666
rect 43038 17614 43090 17666
rect 43262 17614 43314 17666
rect 2830 17502 2882 17554
rect 5742 17502 5794 17554
rect 23326 17502 23378 17554
rect 28590 17502 28642 17554
rect 31950 17502 32002 17554
rect 34302 17502 34354 17554
rect 34862 17502 34914 17554
rect 35534 17502 35586 17554
rect 36094 17502 36146 17554
rect 37438 17502 37490 17554
rect 43710 17502 43762 17554
rect 46174 17502 46226 17554
rect 3950 17390 4002 17442
rect 14366 17390 14418 17442
rect 20526 17390 20578 17442
rect 21758 17390 21810 17442
rect 22094 17390 22146 17442
rect 29374 17390 29426 17442
rect 30158 17390 30210 17442
rect 30494 17390 30546 17442
rect 33518 17390 33570 17442
rect 34750 17390 34802 17442
rect 35198 17390 35250 17442
rect 43486 17390 43538 17442
rect 44158 17390 44210 17442
rect 45838 17390 45890 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 13246 17054 13298 17106
rect 17502 17054 17554 17106
rect 20526 17054 20578 17106
rect 24670 17054 24722 17106
rect 27694 17054 27746 17106
rect 38334 17054 38386 17106
rect 38446 17054 38498 17106
rect 38670 17054 38722 17106
rect 39342 17054 39394 17106
rect 39454 17054 39506 17106
rect 41358 17054 41410 17106
rect 41582 17054 41634 17106
rect 42478 17054 42530 17106
rect 42702 17054 42754 17106
rect 10334 16942 10386 16994
rect 12798 16942 12850 16994
rect 19518 16942 19570 16994
rect 19742 16942 19794 16994
rect 22878 16942 22930 16994
rect 27134 16942 27186 16994
rect 28142 16942 28194 16994
rect 31726 16942 31778 16994
rect 33070 16942 33122 16994
rect 34302 16942 34354 16994
rect 35422 16942 35474 16994
rect 39230 16942 39282 16994
rect 39902 16942 39954 16994
rect 44046 16942 44098 16994
rect 1822 16830 1874 16882
rect 6190 16830 6242 16882
rect 9662 16830 9714 16882
rect 13022 16830 13074 16882
rect 14030 16830 14082 16882
rect 18286 16830 18338 16882
rect 19182 16830 19234 16882
rect 23662 16830 23714 16882
rect 25454 16830 25506 16882
rect 26126 16830 26178 16882
rect 26350 16830 26402 16882
rect 27246 16830 27298 16882
rect 31278 16830 31330 16882
rect 32286 16830 32338 16882
rect 33518 16830 33570 16882
rect 34078 16830 34130 16882
rect 34638 16830 34690 16882
rect 38558 16830 38610 16882
rect 38894 16830 38946 16882
rect 40014 16830 40066 16882
rect 41134 16830 41186 16882
rect 41806 16830 41858 16882
rect 42254 16830 42306 16882
rect 42926 16830 42978 16882
rect 43374 16830 43426 16882
rect 2494 16718 2546 16770
rect 4622 16718 4674 16770
rect 5518 16718 5570 16770
rect 6862 16718 6914 16770
rect 8990 16718 9042 16770
rect 12462 16718 12514 16770
rect 12910 16718 12962 16770
rect 14702 16718 14754 16770
rect 16830 16718 16882 16770
rect 17950 16718 18002 16770
rect 18174 16718 18226 16770
rect 19966 16718 20018 16770
rect 20750 16718 20802 16770
rect 24110 16718 24162 16770
rect 24334 16718 24386 16770
rect 28478 16718 28530 16770
rect 30606 16718 30658 16770
rect 37550 16718 37602 16770
rect 41470 16718 41522 16770
rect 42590 16718 42642 16770
rect 46174 16718 46226 16770
rect 4958 16606 5010 16658
rect 5294 16606 5346 16658
rect 18958 16606 19010 16658
rect 27134 16606 27186 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 4734 16270 4786 16322
rect 11230 16270 11282 16322
rect 11566 16270 11618 16322
rect 14926 16270 14978 16322
rect 15598 16270 15650 16322
rect 15934 16270 15986 16322
rect 17726 16270 17778 16322
rect 18398 16270 18450 16322
rect 21198 16270 21250 16322
rect 21422 16270 21474 16322
rect 30606 16270 30658 16322
rect 45726 16270 45778 16322
rect 46174 16270 46226 16322
rect 8654 16158 8706 16210
rect 10558 16158 10610 16210
rect 11790 16158 11842 16210
rect 17950 16158 18002 16210
rect 19406 16158 19458 16210
rect 20750 16158 20802 16210
rect 21422 16158 21474 16210
rect 22990 16158 23042 16210
rect 24670 16158 24722 16210
rect 26798 16158 26850 16210
rect 28590 16158 28642 16210
rect 30046 16158 30098 16210
rect 30494 16158 30546 16210
rect 31390 16158 31442 16210
rect 31838 16158 31890 16210
rect 32062 16158 32114 16210
rect 35198 16158 35250 16210
rect 35646 16158 35698 16210
rect 37214 16158 37266 16210
rect 38222 16158 38274 16210
rect 40350 16158 40402 16210
rect 41470 16158 41522 16210
rect 43598 16158 43650 16210
rect 44830 16158 44882 16210
rect 45278 16158 45330 16210
rect 45838 16158 45890 16210
rect 4062 16046 4114 16098
rect 4286 16046 4338 16098
rect 5854 16046 5906 16098
rect 8878 16046 8930 16098
rect 9550 16046 9602 16098
rect 9774 16046 9826 16098
rect 10110 16046 10162 16098
rect 16494 16046 16546 16098
rect 16942 16046 16994 16098
rect 17502 16046 17554 16098
rect 18958 16046 19010 16098
rect 19182 16046 19234 16098
rect 22430 16046 22482 16098
rect 23886 16046 23938 16098
rect 27582 16046 27634 16098
rect 27694 16046 27746 16098
rect 29486 16046 29538 16098
rect 29710 16046 29762 16098
rect 29934 16046 29986 16098
rect 32622 16046 32674 16098
rect 33182 16046 33234 16098
rect 33854 16046 33906 16098
rect 35086 16046 35138 16098
rect 36094 16046 36146 16098
rect 37438 16046 37490 16098
rect 40798 16046 40850 16098
rect 4846 15934 4898 15986
rect 5070 15934 5122 15986
rect 9662 15934 9714 15986
rect 10446 15934 10498 15986
rect 15038 15934 15090 15986
rect 15262 15934 15314 15986
rect 16382 15934 16434 15986
rect 20302 15934 20354 15986
rect 27806 15934 27858 15986
rect 30046 15934 30098 15986
rect 36430 15934 36482 15986
rect 44046 15934 44098 15986
rect 3502 15822 3554 15874
rect 3726 15822 3778 15874
rect 5630 15822 5682 15874
rect 5742 15822 5794 15874
rect 6078 15822 6130 15874
rect 9214 15822 9266 15874
rect 10670 15822 10722 15874
rect 15822 15822 15874 15874
rect 16270 15822 16322 15874
rect 18958 15822 19010 15874
rect 21870 15822 21922 15874
rect 27134 15822 27186 15874
rect 28478 15822 28530 15874
rect 32958 15822 33010 15874
rect 33630 15822 33682 15874
rect 43934 15822 43986 15874
rect 44942 15822 44994 15874
rect 45390 15822 45442 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 10110 15486 10162 15538
rect 14366 15486 14418 15538
rect 14702 15486 14754 15538
rect 15038 15486 15090 15538
rect 16830 15486 16882 15538
rect 17614 15486 17666 15538
rect 18062 15486 18114 15538
rect 18174 15486 18226 15538
rect 19182 15486 19234 15538
rect 19294 15486 19346 15538
rect 19406 15486 19458 15538
rect 21534 15486 21586 15538
rect 22542 15486 22594 15538
rect 26462 15486 26514 15538
rect 27806 15486 27858 15538
rect 28478 15486 28530 15538
rect 39790 15486 39842 15538
rect 17950 15374 18002 15426
rect 20862 15374 20914 15426
rect 27918 15374 27970 15426
rect 41134 15374 41186 15426
rect 1822 15262 1874 15314
rect 6078 15262 6130 15314
rect 10334 15262 10386 15314
rect 10782 15262 10834 15314
rect 11118 15262 11170 15314
rect 15262 15262 15314 15314
rect 18734 15262 18786 15314
rect 19742 15262 19794 15314
rect 19966 15262 20018 15314
rect 21086 15262 21138 15314
rect 25342 15262 25394 15314
rect 25790 15262 25842 15314
rect 26238 15262 26290 15314
rect 26462 15262 26514 15314
rect 26686 15262 26738 15314
rect 27358 15262 27410 15314
rect 27582 15262 27634 15314
rect 28030 15262 28082 15314
rect 28590 15262 28642 15314
rect 32174 15262 32226 15314
rect 37774 15262 37826 15314
rect 38670 15262 38722 15314
rect 45838 15262 45890 15314
rect 2494 15150 2546 15202
rect 4622 15150 4674 15202
rect 6750 15150 6802 15202
rect 8878 15150 8930 15202
rect 10222 15150 10274 15202
rect 11902 15150 11954 15202
rect 14030 15150 14082 15202
rect 17502 15150 17554 15202
rect 20302 15150 20354 15202
rect 22094 15150 22146 15202
rect 25230 15150 25282 15202
rect 25566 15150 25618 15202
rect 26910 15150 26962 15202
rect 27134 15150 27186 15202
rect 29262 15150 29314 15202
rect 31390 15150 31442 15202
rect 33630 15150 33682 15202
rect 40238 15150 40290 15202
rect 20190 15038 20242 15090
rect 38894 15038 38946 15090
rect 39230 15038 39282 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 3166 14702 3218 14754
rect 22542 14702 22594 14754
rect 26574 14702 26626 14754
rect 27134 14702 27186 14754
rect 4846 14590 4898 14642
rect 7758 14590 7810 14642
rect 9886 14590 9938 14642
rect 10222 14590 10274 14642
rect 12014 14590 12066 14642
rect 13022 14590 13074 14642
rect 15822 14590 15874 14642
rect 16270 14590 16322 14642
rect 18398 14590 18450 14642
rect 20526 14590 20578 14642
rect 23774 14590 23826 14642
rect 25902 14590 25954 14642
rect 30382 14590 30434 14642
rect 30830 14590 30882 14642
rect 30942 14590 30994 14642
rect 33182 14590 33234 14642
rect 36094 14590 36146 14642
rect 38334 14590 38386 14642
rect 42702 14590 42754 14642
rect 4062 14478 4114 14530
rect 4398 14478 4450 14530
rect 7086 14478 7138 14530
rect 10894 14478 10946 14530
rect 11118 14478 11170 14530
rect 11790 14478 11842 14530
rect 12238 14478 12290 14530
rect 13694 14478 13746 14530
rect 14142 14478 14194 14530
rect 14926 14478 14978 14530
rect 15486 14478 15538 14530
rect 19182 14478 19234 14530
rect 21422 14478 21474 14530
rect 23102 14478 23154 14530
rect 28030 14478 28082 14530
rect 28478 14478 28530 14530
rect 29374 14478 29426 14530
rect 29822 14478 29874 14530
rect 30046 14478 30098 14530
rect 32286 14478 32338 14530
rect 32734 14478 32786 14530
rect 34526 14478 34578 14530
rect 34862 14478 34914 14530
rect 35870 14478 35922 14530
rect 36206 14478 36258 14530
rect 37214 14478 37266 14530
rect 37998 14478 38050 14530
rect 41134 14478 41186 14530
rect 3278 14366 3330 14418
rect 3502 14366 3554 14418
rect 5630 14366 5682 14418
rect 5966 14366 6018 14418
rect 6638 14366 6690 14418
rect 10334 14366 10386 14418
rect 10558 14366 10610 14418
rect 12462 14366 12514 14418
rect 13582 14366 13634 14418
rect 19854 14366 19906 14418
rect 20078 14366 20130 14418
rect 21646 14366 21698 14418
rect 22430 14366 22482 14418
rect 27134 14366 27186 14418
rect 27246 14366 27298 14418
rect 27694 14366 27746 14418
rect 30382 14366 30434 14418
rect 31950 14366 32002 14418
rect 33518 14366 33570 14418
rect 33854 14366 33906 14418
rect 37550 14366 37602 14418
rect 37886 14366 37938 14418
rect 40462 14366 40514 14418
rect 41694 14366 41746 14418
rect 43150 14366 43202 14418
rect 43710 14366 43762 14418
rect 3838 14254 3890 14306
rect 3950 14254 4002 14306
rect 6302 14254 6354 14306
rect 11454 14254 11506 14306
rect 13470 14254 13522 14306
rect 14702 14254 14754 14306
rect 22206 14254 22258 14306
rect 22542 14254 22594 14306
rect 26350 14254 26402 14306
rect 26462 14254 26514 14306
rect 29038 14254 29090 14306
rect 29262 14254 29314 14306
rect 30270 14254 30322 14306
rect 31726 14254 31778 14306
rect 34190 14254 34242 14306
rect 34974 14254 35026 14306
rect 35086 14254 35138 14306
rect 35310 14254 35362 14306
rect 36430 14254 36482 14306
rect 36990 14254 37042 14306
rect 41806 14254 41858 14306
rect 42030 14254 42082 14306
rect 42590 14254 42642 14306
rect 43038 14254 43090 14306
rect 44046 14254 44098 14306
rect 44830 14254 44882 14306
rect 45278 14254 45330 14306
rect 45726 14254 45778 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 5854 13918 5906 13970
rect 6190 13918 6242 13970
rect 6974 13918 7026 13970
rect 7982 13918 8034 13970
rect 8878 13918 8930 13970
rect 9550 13918 9602 13970
rect 10446 13918 10498 13970
rect 10558 13918 10610 13970
rect 10670 13918 10722 13970
rect 11454 13918 11506 13970
rect 13470 13918 13522 13970
rect 15710 13918 15762 13970
rect 16158 13918 16210 13970
rect 23886 13918 23938 13970
rect 24558 13918 24610 13970
rect 29598 13918 29650 13970
rect 32174 13918 32226 13970
rect 33294 13918 33346 13970
rect 33742 13918 33794 13970
rect 39566 13918 39618 13970
rect 42926 13918 42978 13970
rect 8766 13806 8818 13858
rect 8990 13806 9042 13858
rect 11566 13806 11618 13858
rect 12126 13806 12178 13858
rect 13134 13806 13186 13858
rect 13806 13806 13858 13858
rect 14702 13806 14754 13858
rect 15374 13806 15426 13858
rect 22206 13806 22258 13858
rect 23550 13806 23602 13858
rect 23662 13806 23714 13858
rect 26798 13806 26850 13858
rect 26910 13806 26962 13858
rect 27694 13806 27746 13858
rect 28030 13806 28082 13858
rect 30270 13806 30322 13858
rect 34302 13806 34354 13858
rect 35422 13806 35474 13858
rect 38894 13806 38946 13858
rect 39230 13806 39282 13858
rect 40350 13806 40402 13858
rect 41246 13806 41298 13858
rect 42478 13806 42530 13858
rect 45390 13806 45442 13858
rect 1822 13694 1874 13746
rect 5182 13694 5234 13746
rect 7534 13694 7586 13746
rect 9886 13694 9938 13746
rect 10110 13694 10162 13746
rect 11118 13694 11170 13746
rect 12014 13694 12066 13746
rect 12238 13694 12290 13746
rect 12574 13694 12626 13746
rect 14030 13694 14082 13746
rect 14926 13694 14978 13746
rect 16718 13694 16770 13746
rect 22990 13694 23042 13746
rect 24222 13694 24274 13746
rect 24558 13694 24610 13746
rect 25566 13694 25618 13746
rect 26574 13694 26626 13746
rect 27470 13694 27522 13746
rect 28478 13694 28530 13746
rect 29038 13694 29090 13746
rect 29822 13694 29874 13746
rect 30046 13694 30098 13746
rect 30830 13694 30882 13746
rect 31278 13694 31330 13746
rect 34078 13694 34130 13746
rect 34638 13694 34690 13746
rect 38446 13694 38498 13746
rect 40014 13694 40066 13746
rect 41470 13694 41522 13746
rect 42142 13694 42194 13746
rect 42366 13694 42418 13746
rect 46062 13694 46114 13746
rect 2494 13582 2546 13634
rect 4622 13582 4674 13634
rect 4958 13582 5010 13634
rect 6750 13582 6802 13634
rect 18398 13582 18450 13634
rect 20078 13582 20130 13634
rect 25790 13582 25842 13634
rect 32510 13582 32562 13634
rect 37550 13582 37602 13634
rect 37998 13582 38050 13634
rect 41806 13582 41858 13634
rect 43262 13582 43314 13634
rect 5518 13470 5570 13522
rect 7310 13470 7362 13522
rect 11454 13470 11506 13522
rect 12910 13470 12962 13522
rect 18286 13470 18338 13522
rect 24446 13470 24498 13522
rect 25230 13470 25282 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 2942 13134 2994 13186
rect 4734 13134 4786 13186
rect 27022 13134 27074 13186
rect 38446 13134 38498 13186
rect 8430 13022 8482 13074
rect 19182 13022 19234 13074
rect 23550 13022 23602 13074
rect 27918 13022 27970 13074
rect 29710 13022 29762 13074
rect 34302 13022 34354 13074
rect 36430 13022 36482 13074
rect 38334 13022 38386 13074
rect 38782 13022 38834 13074
rect 42366 13022 42418 13074
rect 3838 12910 3890 12962
rect 4510 12910 4562 12962
rect 5630 12910 5682 12962
rect 5854 12910 5906 12962
rect 12910 12910 12962 12962
rect 13694 12910 13746 12962
rect 14254 12910 14306 12962
rect 16382 12910 16434 12962
rect 21310 12910 21362 12962
rect 27358 12910 27410 12962
rect 27694 12910 27746 12962
rect 27806 12910 27858 12962
rect 28030 12910 28082 12962
rect 32622 12910 32674 12962
rect 33630 12910 33682 12962
rect 36878 12910 36930 12962
rect 37214 12910 37266 12962
rect 37998 12910 38050 12962
rect 40686 12910 40738 12962
rect 41134 12910 41186 12962
rect 41358 12910 41410 12962
rect 42478 12910 42530 12962
rect 43150 12910 43202 12962
rect 43486 12910 43538 12962
rect 43710 12910 43762 12962
rect 46062 12910 46114 12962
rect 3054 12798 3106 12850
rect 3278 12798 3330 12850
rect 3726 12798 3778 12850
rect 6078 12798 6130 12850
rect 17054 12798 17106 12850
rect 19518 12798 19570 12850
rect 26910 12798 26962 12850
rect 28590 12798 28642 12850
rect 29262 12798 29314 12850
rect 29374 12798 29426 12850
rect 31838 12798 31890 12850
rect 37550 12798 37602 12850
rect 39342 12798 39394 12850
rect 39902 12798 39954 12850
rect 40350 12798 40402 12850
rect 40798 12798 40850 12850
rect 45502 12798 45554 12850
rect 45838 12798 45890 12850
rect 3614 12686 3666 12738
rect 4062 12686 4114 12738
rect 5070 12686 5122 12738
rect 5742 12686 5794 12738
rect 13470 12686 13522 12738
rect 19630 12686 19682 12738
rect 19854 12686 19906 12738
rect 20750 12686 20802 12738
rect 33182 12686 33234 12738
rect 37214 12686 37266 12738
rect 37886 12686 37938 12738
rect 38894 12686 38946 12738
rect 39230 12686 39282 12738
rect 39790 12686 39842 12738
rect 40238 12686 40290 12738
rect 41582 12686 41634 12738
rect 41694 12686 41746 12738
rect 44046 12686 44098 12738
rect 45166 12686 45218 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 5630 12350 5682 12402
rect 9662 12350 9714 12402
rect 10110 12350 10162 12402
rect 15934 12350 15986 12402
rect 16718 12350 16770 12402
rect 17838 12350 17890 12402
rect 18174 12350 18226 12402
rect 21086 12350 21138 12402
rect 21646 12350 21698 12402
rect 30158 12350 30210 12402
rect 30270 12350 30322 12402
rect 30494 12350 30546 12402
rect 33518 12350 33570 12402
rect 34414 12350 34466 12402
rect 39118 12350 39170 12402
rect 5518 12238 5570 12290
rect 7310 12238 7362 12290
rect 13470 12238 13522 12290
rect 16270 12238 16322 12290
rect 16606 12238 16658 12290
rect 18398 12238 18450 12290
rect 18846 12238 18898 12290
rect 19294 12238 19346 12290
rect 20414 12238 20466 12290
rect 21982 12238 22034 12290
rect 23998 12238 24050 12290
rect 27134 12238 27186 12290
rect 27246 12238 27298 12290
rect 27694 12238 27746 12290
rect 27806 12238 27858 12290
rect 28926 12238 28978 12290
rect 29150 12238 29202 12290
rect 29934 12238 29986 12290
rect 34862 12238 34914 12290
rect 34974 12238 35026 12290
rect 35086 12238 35138 12290
rect 35758 12238 35810 12290
rect 36654 12238 36706 12290
rect 40126 12238 40178 12290
rect 41358 12238 41410 12290
rect 42366 12238 42418 12290
rect 42814 12238 42866 12290
rect 45390 12238 45442 12290
rect 1822 12126 1874 12178
rect 5742 12126 5794 12178
rect 6190 12126 6242 12178
rect 6414 12126 6466 12178
rect 6638 12126 6690 12178
rect 7086 12126 7138 12178
rect 7534 12126 7586 12178
rect 11342 12126 11394 12178
rect 12686 12126 12738 12178
rect 16942 12126 16994 12178
rect 17390 12126 17442 12178
rect 17726 12126 17778 12178
rect 18062 12126 18114 12178
rect 18510 12126 18562 12178
rect 19070 12126 19122 12178
rect 20078 12126 20130 12178
rect 21422 12126 21474 12178
rect 22430 12126 22482 12178
rect 22878 12126 22930 12178
rect 23662 12126 23714 12178
rect 23886 12126 23938 12178
rect 24110 12126 24162 12178
rect 25342 12126 25394 12178
rect 25566 12126 25618 12178
rect 25790 12126 25842 12178
rect 26462 12126 26514 12178
rect 26910 12126 26962 12178
rect 28030 12126 28082 12178
rect 29374 12126 29426 12178
rect 29598 12126 29650 12178
rect 30382 12126 30434 12178
rect 33070 12126 33122 12178
rect 33294 12126 33346 12178
rect 33742 12126 33794 12178
rect 35982 12126 36034 12178
rect 36430 12126 36482 12178
rect 37326 12126 37378 12178
rect 39454 12126 39506 12178
rect 40014 12126 40066 12178
rect 41134 12126 41186 12178
rect 41246 12126 41298 12178
rect 41806 12126 41858 12178
rect 46062 12126 46114 12178
rect 2494 12014 2546 12066
rect 4622 12014 4674 12066
rect 6862 12014 6914 12066
rect 10110 12014 10162 12066
rect 10334 12014 10386 12066
rect 10670 12014 10722 12066
rect 11454 12014 11506 12066
rect 15598 12014 15650 12066
rect 25678 12014 25730 12066
rect 26126 12014 26178 12066
rect 26686 12014 26738 12066
rect 28478 12014 28530 12066
rect 29262 12014 29314 12066
rect 31054 12014 31106 12066
rect 31502 12014 31554 12066
rect 32174 12014 32226 12066
rect 32398 12014 32450 12066
rect 33182 12014 33234 12066
rect 35646 12014 35698 12066
rect 38110 12014 38162 12066
rect 39678 12014 39730 12066
rect 43262 12014 43314 12066
rect 23214 11902 23266 11954
rect 28590 11902 28642 11954
rect 30830 11902 30882 11954
rect 31278 11902 31330 11954
rect 31502 11902 31554 11954
rect 31726 11902 31778 11954
rect 32510 11902 32562 11954
rect 38222 11902 38274 11954
rect 42030 11902 42082 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 18734 11566 18786 11618
rect 27582 11566 27634 11618
rect 41582 11566 41634 11618
rect 42926 11566 42978 11618
rect 6078 11454 6130 11506
rect 10110 11454 10162 11506
rect 12238 11454 12290 11506
rect 12574 11454 12626 11506
rect 17166 11454 17218 11506
rect 19070 11454 19122 11506
rect 20190 11454 20242 11506
rect 24558 11454 24610 11506
rect 26686 11454 26738 11506
rect 34526 11454 34578 11506
rect 34862 11454 34914 11506
rect 35086 11454 35138 11506
rect 37102 11454 37154 11506
rect 37774 11454 37826 11506
rect 38782 11454 38834 11506
rect 40686 11454 40738 11506
rect 41358 11454 41410 11506
rect 4846 11342 4898 11394
rect 5070 11342 5122 11394
rect 8878 11342 8930 11394
rect 9326 11342 9378 11394
rect 15598 11342 15650 11394
rect 16270 11342 16322 11394
rect 18398 11342 18450 11394
rect 19294 11342 19346 11394
rect 20302 11342 20354 11394
rect 21646 11342 21698 11394
rect 23774 11342 23826 11394
rect 28366 11342 28418 11394
rect 28590 11342 28642 11394
rect 34414 11342 34466 11394
rect 35870 11342 35922 11394
rect 36206 11342 36258 11394
rect 38222 11342 38274 11394
rect 38558 11342 38610 11394
rect 39006 11342 39058 11394
rect 39118 11342 39170 11394
rect 39454 11342 39506 11394
rect 41918 11342 41970 11394
rect 42366 11342 42418 11394
rect 42478 11342 42530 11394
rect 42702 11342 42754 11394
rect 43038 11342 43090 11394
rect 43822 11342 43874 11394
rect 44830 11342 44882 11394
rect 4510 11230 4562 11282
rect 8206 11230 8258 11282
rect 12910 11230 12962 11282
rect 13358 11230 13410 11282
rect 13582 11230 13634 11282
rect 13694 11230 13746 11282
rect 15262 11230 15314 11282
rect 15374 11230 15426 11282
rect 19966 11230 20018 11282
rect 27694 11230 27746 11282
rect 31278 11230 31330 11282
rect 35982 11230 36034 11282
rect 40126 11230 40178 11282
rect 41022 11230 41074 11282
rect 4622 11118 4674 11170
rect 12686 11118 12738 11170
rect 14926 11118 14978 11170
rect 15150 11118 15202 11170
rect 16046 11118 16098 11170
rect 16158 11118 16210 11170
rect 18622 11118 18674 11170
rect 19630 11118 19682 11170
rect 21310 11118 21362 11170
rect 22430 11118 22482 11170
rect 27246 11118 27298 11170
rect 28030 11118 28082 11170
rect 35198 11118 35250 11170
rect 37214 11118 37266 11170
rect 37662 11118 37714 11170
rect 37774 11118 37826 11170
rect 37998 11118 38050 11170
rect 38782 11118 38834 11170
rect 39902 11118 39954 11170
rect 40014 11118 40066 11170
rect 40798 11118 40850 11170
rect 43598 11118 43650 11170
rect 45166 11118 45218 11170
rect 45838 11118 45890 11170
rect 46174 11118 46226 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 5406 10782 5458 10834
rect 17390 10782 17442 10834
rect 31950 10782 32002 10834
rect 32062 10782 32114 10834
rect 32286 10782 32338 10834
rect 36430 10782 36482 10834
rect 36542 10782 36594 10834
rect 38334 10782 38386 10834
rect 39454 10782 39506 10834
rect 41470 10782 41522 10834
rect 2830 10670 2882 10722
rect 5630 10670 5682 10722
rect 6414 10670 6466 10722
rect 6526 10670 6578 10722
rect 8094 10670 8146 10722
rect 8542 10670 8594 10722
rect 11230 10670 11282 10722
rect 12574 10670 12626 10722
rect 15486 10670 15538 10722
rect 16046 10670 16098 10722
rect 19070 10670 19122 10722
rect 26014 10670 26066 10722
rect 30606 10670 30658 10722
rect 32510 10670 32562 10722
rect 33854 10670 33906 10722
rect 36654 10670 36706 10722
rect 37438 10670 37490 10722
rect 38222 10670 38274 10722
rect 39230 10670 39282 10722
rect 40014 10670 40066 10722
rect 42366 10670 42418 10722
rect 45390 10670 45442 10722
rect 2046 10558 2098 10610
rect 6190 10558 6242 10610
rect 7758 10558 7810 10610
rect 7982 10558 8034 10610
rect 10894 10558 10946 10610
rect 11454 10558 11506 10610
rect 11902 10558 11954 10610
rect 15822 10558 15874 10610
rect 17502 10558 17554 10610
rect 18398 10558 18450 10610
rect 21646 10558 21698 10610
rect 25342 10558 25394 10610
rect 31278 10558 31330 10610
rect 33070 10558 33122 10610
rect 36766 10558 36818 10610
rect 37102 10558 37154 10610
rect 37774 10558 37826 10610
rect 39566 10558 39618 10610
rect 41246 10558 41298 10610
rect 42590 10558 42642 10610
rect 46062 10558 46114 10610
rect 4958 10446 5010 10498
rect 5294 10446 5346 10498
rect 11006 10446 11058 10498
rect 14702 10446 14754 10498
rect 15038 10446 15090 10498
rect 15598 10446 15650 10498
rect 21198 10446 21250 10498
rect 22318 10446 22370 10498
rect 24446 10446 24498 10498
rect 28142 10446 28194 10498
rect 28478 10446 28530 10498
rect 32174 10446 32226 10498
rect 35982 10446 36034 10498
rect 37662 10446 37714 10498
rect 38894 10446 38946 10498
rect 42030 10446 42082 10498
rect 43262 10446 43314 10498
rect 6974 10334 7026 10386
rect 7646 10334 7698 10386
rect 15150 10334 15202 10386
rect 38334 10334 38386 10386
rect 39006 10334 39058 10386
rect 39902 10334 39954 10386
rect 40238 10334 40290 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 42926 9998 42978 10050
rect 4622 9886 4674 9938
rect 9438 9886 9490 9938
rect 11566 9886 11618 9938
rect 12014 9886 12066 9938
rect 14478 9886 14530 9938
rect 15598 9886 15650 9938
rect 17726 9886 17778 9938
rect 23326 9886 23378 9938
rect 24222 9886 24274 9938
rect 27694 9886 27746 9938
rect 28590 9886 28642 9938
rect 32062 9886 32114 9938
rect 32510 9886 32562 9938
rect 32958 9886 33010 9938
rect 33294 9886 33346 9938
rect 35422 9886 35474 9938
rect 42142 9886 42194 9938
rect 1822 9774 1874 9826
rect 7086 9774 7138 9826
rect 8766 9774 8818 9826
rect 11902 9774 11954 9826
rect 14814 9774 14866 9826
rect 21646 9774 21698 9826
rect 22990 9774 23042 9826
rect 27134 9774 27186 9826
rect 29262 9774 29314 9826
rect 36094 9774 36146 9826
rect 38894 9774 38946 9826
rect 39454 9774 39506 9826
rect 40014 9774 40066 9826
rect 40462 9774 40514 9826
rect 40798 9774 40850 9826
rect 41022 9774 41074 9826
rect 41694 9774 41746 9826
rect 42366 9774 42418 9826
rect 42702 9774 42754 9826
rect 2494 9662 2546 9714
rect 12350 9662 12402 9714
rect 13470 9662 13522 9714
rect 13806 9662 13858 9714
rect 18398 9662 18450 9714
rect 20638 9662 20690 9714
rect 22654 9662 22706 9714
rect 23662 9662 23714 9714
rect 26350 9662 26402 9714
rect 29934 9662 29986 9714
rect 38334 9662 38386 9714
rect 38670 9662 38722 9714
rect 39006 9662 39058 9714
rect 43262 9662 43314 9714
rect 45166 9662 45218 9714
rect 46174 9662 46226 9714
rect 7534 9550 7586 9602
rect 7646 9550 7698 9602
rect 7758 9550 7810 9602
rect 12126 9550 12178 9602
rect 18174 9550 18226 9602
rect 18286 9550 18338 9602
rect 20750 9550 20802 9602
rect 22206 9550 22258 9602
rect 23438 9550 23490 9602
rect 28142 9550 28194 9602
rect 37102 9550 37154 9602
rect 37886 9550 37938 9602
rect 38222 9550 38274 9602
rect 40686 9550 40738 9602
rect 41806 9550 41858 9602
rect 41918 9550 41970 9602
rect 43598 9550 43650 9602
rect 43934 9550 43986 9602
rect 44830 9550 44882 9602
rect 45838 9550 45890 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2270 9214 2322 9266
rect 11230 9214 11282 9266
rect 13022 9214 13074 9266
rect 14702 9214 14754 9266
rect 16046 9214 16098 9266
rect 16606 9214 16658 9266
rect 2718 9102 2770 9154
rect 10110 9102 10162 9154
rect 11342 9102 11394 9154
rect 11902 9102 11954 9154
rect 12126 9102 12178 9154
rect 14030 9102 14082 9154
rect 14366 9102 14418 9154
rect 15150 9102 15202 9154
rect 15710 9102 15762 9154
rect 24782 9214 24834 9266
rect 26574 9214 26626 9266
rect 27134 9214 27186 9266
rect 27470 9214 27522 9266
rect 27918 9214 27970 9266
rect 28814 9214 28866 9266
rect 30494 9214 30546 9266
rect 33630 9214 33682 9266
rect 39342 9214 39394 9266
rect 39566 9214 39618 9266
rect 39902 9214 39954 9266
rect 41134 9214 41186 9266
rect 41358 9214 41410 9266
rect 41470 9214 41522 9266
rect 25790 9102 25842 9154
rect 26014 9102 26066 9154
rect 30158 9102 30210 9154
rect 30606 9102 30658 9154
rect 39118 9102 39170 9154
rect 40910 9102 40962 9154
rect 45390 9102 45442 9154
rect 8542 8990 8594 9042
rect 9438 8990 9490 9042
rect 9774 8990 9826 9042
rect 11790 8990 11842 9042
rect 12238 8990 12290 9042
rect 12686 8990 12738 9042
rect 13694 8990 13746 9042
rect 15486 8990 15538 9042
rect 15710 8990 15762 9042
rect 17390 8990 17442 9042
rect 23550 8990 23602 9042
rect 25230 8990 25282 9042
rect 25566 8990 25618 9042
rect 31390 8990 31442 9042
rect 33182 8990 33234 9042
rect 33406 8990 33458 9042
rect 33854 8990 33906 9042
rect 34302 8990 34354 9042
rect 37550 8990 37602 9042
rect 37998 8990 38050 9042
rect 40126 8990 40178 9042
rect 40350 8990 40402 9042
rect 42254 8990 42306 9042
rect 42814 8990 42866 9042
rect 46062 8990 46114 9042
rect 2606 8878 2658 8930
rect 3614 8878 3666 8930
rect 8990 8878 9042 8930
rect 9662 8878 9714 8930
rect 10670 8878 10722 8930
rect 16158 8878 16210 8930
rect 16718 8878 16770 8930
rect 18174 8878 18226 8930
rect 20302 8878 20354 8930
rect 20638 8878 20690 8930
rect 22766 8878 22818 8930
rect 23998 8878 24050 8930
rect 25678 8878 25730 8930
rect 28478 8878 28530 8930
rect 29262 8878 29314 8930
rect 29710 8878 29762 8930
rect 31502 8878 31554 8930
rect 32398 8878 32450 8930
rect 33518 8878 33570 8930
rect 34974 8878 35026 8930
rect 37102 8878 37154 8930
rect 39454 8878 39506 8930
rect 39790 8878 39842 8930
rect 41358 8878 41410 8930
rect 42926 8878 42978 8930
rect 43262 8878 43314 8930
rect 2942 8766 2994 8818
rect 11230 8766 11282 8818
rect 15262 8766 15314 8818
rect 16830 8766 16882 8818
rect 31838 8766 31890 8818
rect 32286 8766 32338 8818
rect 37774 8766 37826 8818
rect 38446 8766 38498 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 22318 8430 22370 8482
rect 22654 8430 22706 8482
rect 23326 8430 23378 8482
rect 38894 8430 38946 8482
rect 41022 8430 41074 8482
rect 3502 8318 3554 8370
rect 4846 8318 4898 8370
rect 6414 8318 6466 8370
rect 8542 8318 8594 8370
rect 11118 8318 11170 8370
rect 14814 8318 14866 8370
rect 23662 8318 23714 8370
rect 25118 8318 25170 8370
rect 27358 8318 27410 8370
rect 28142 8318 28194 8370
rect 31614 8318 31666 8370
rect 33742 8318 33794 8370
rect 34414 8318 34466 8370
rect 38670 8318 38722 8370
rect 40126 8318 40178 8370
rect 40910 8318 40962 8370
rect 41358 8318 41410 8370
rect 43486 8318 43538 8370
rect 44830 8318 44882 8370
rect 3054 8206 3106 8258
rect 4062 8206 4114 8258
rect 4622 8206 4674 8258
rect 5630 8206 5682 8258
rect 9326 8206 9378 8258
rect 9438 8206 9490 8258
rect 9662 8206 9714 8258
rect 11454 8206 11506 8258
rect 19742 8206 19794 8258
rect 20302 8206 20354 8258
rect 20638 8206 20690 8258
rect 21982 8206 22034 8258
rect 22430 8206 22482 8258
rect 24110 8206 24162 8258
rect 24334 8206 24386 8258
rect 25006 8206 25058 8258
rect 25566 8206 25618 8258
rect 26126 8206 26178 8258
rect 26350 8206 26402 8258
rect 27470 8206 27522 8258
rect 27806 8206 27858 8258
rect 29038 8206 29090 8258
rect 29374 8206 29426 8258
rect 29598 8206 29650 8258
rect 30494 8206 30546 8258
rect 30942 8206 30994 8258
rect 34078 8206 34130 8258
rect 34526 8206 34578 8258
rect 34750 8206 34802 8258
rect 35310 8206 35362 8258
rect 36990 8206 37042 8258
rect 37214 8206 37266 8258
rect 37438 8206 37490 8258
rect 37662 8206 37714 8258
rect 37998 8206 38050 8258
rect 38558 8206 38610 8258
rect 38782 8206 38834 8258
rect 40014 8206 40066 8258
rect 44270 8206 44322 8258
rect 45054 8206 45106 8258
rect 45390 8206 45442 8258
rect 45950 8206 46002 8258
rect 4286 8094 4338 8146
rect 10222 8094 10274 8146
rect 10446 8094 10498 8146
rect 10782 8094 10834 8146
rect 12910 8094 12962 8146
rect 14142 8094 14194 8146
rect 21758 8094 21810 8146
rect 25342 8094 25394 8146
rect 25902 8094 25954 8146
rect 28478 8094 28530 8146
rect 29262 8094 29314 8146
rect 35086 8094 35138 8146
rect 36094 8094 36146 8146
rect 2270 7982 2322 8034
rect 2606 7982 2658 8034
rect 2830 7982 2882 8034
rect 2942 7982 2994 8034
rect 3390 7982 3442 8034
rect 3614 7982 3666 8034
rect 8878 7982 8930 8034
rect 10334 7982 10386 8034
rect 13806 7982 13858 8034
rect 20190 7982 20242 8034
rect 20414 7982 20466 8034
rect 20526 7982 20578 8034
rect 21422 7982 21474 8034
rect 22542 7982 22594 8034
rect 23214 7982 23266 8034
rect 24446 7982 24498 8034
rect 24670 7982 24722 8034
rect 26014 7982 26066 8034
rect 27694 7982 27746 8034
rect 28254 7982 28306 8034
rect 30158 7982 30210 8034
rect 34302 7982 34354 8034
rect 36206 7982 36258 8034
rect 37102 7982 37154 8034
rect 45726 7982 45778 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 16606 7646 16658 7698
rect 20638 7646 20690 7698
rect 22990 7646 23042 7698
rect 23662 7646 23714 7698
rect 30830 7646 30882 7698
rect 32062 7646 32114 7698
rect 32174 7646 32226 7698
rect 33182 7646 33234 7698
rect 34078 7646 34130 7698
rect 34526 7646 34578 7698
rect 38558 7646 38610 7698
rect 40014 7646 40066 7698
rect 4958 7534 5010 7586
rect 5182 7534 5234 7586
rect 10334 7534 10386 7586
rect 13918 7534 13970 7586
rect 16830 7534 16882 7586
rect 20302 7534 20354 7586
rect 22206 7534 22258 7586
rect 22878 7534 22930 7586
rect 25230 7534 25282 7586
rect 25566 7534 25618 7586
rect 26238 7534 26290 7586
rect 26350 7534 26402 7586
rect 28030 7534 28082 7586
rect 31502 7534 31554 7586
rect 32510 7534 32562 7586
rect 33630 7534 33682 7586
rect 33966 7534 34018 7586
rect 36990 7534 37042 7586
rect 39678 7534 39730 7586
rect 39902 7534 39954 7586
rect 40238 7534 40290 7586
rect 44158 7534 44210 7586
rect 4510 7422 4562 7474
rect 5630 7422 5682 7474
rect 9550 7422 9602 7474
rect 13134 7422 13186 7474
rect 17390 7422 17442 7474
rect 20526 7422 20578 7474
rect 20750 7422 20802 7474
rect 20974 7422 21026 7474
rect 21870 7422 21922 7474
rect 22654 7422 22706 7474
rect 22766 7422 22818 7474
rect 23214 7422 23266 7474
rect 24334 7422 24386 7474
rect 24558 7422 24610 7474
rect 26126 7422 26178 7474
rect 27358 7422 27410 7474
rect 31278 7422 31330 7474
rect 31838 7422 31890 7474
rect 32286 7422 32338 7474
rect 34414 7422 34466 7474
rect 37662 7422 37714 7474
rect 38334 7422 38386 7474
rect 38446 7422 38498 7474
rect 38670 7422 38722 7474
rect 38894 7422 38946 7474
rect 44718 7422 44770 7474
rect 1710 7310 1762 7362
rect 3838 7310 3890 7362
rect 5070 7310 5122 7362
rect 6414 7310 6466 7362
rect 8542 7310 8594 7362
rect 8990 7310 9042 7362
rect 12462 7310 12514 7362
rect 16046 7310 16098 7362
rect 16494 7310 16546 7362
rect 18510 7310 18562 7362
rect 21646 7310 21698 7362
rect 22094 7310 22146 7362
rect 24222 7310 24274 7362
rect 26798 7310 26850 7362
rect 30158 7310 30210 7362
rect 34862 7310 34914 7362
rect 39342 7310 39394 7362
rect 24670 7198 24722 7250
rect 39230 7198 39282 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 3838 6862 3890 6914
rect 12238 6862 12290 6914
rect 12910 6862 12962 6914
rect 21870 6862 21922 6914
rect 22654 6862 22706 6914
rect 23438 6862 23490 6914
rect 43598 6862 43650 6914
rect 43710 6862 43762 6914
rect 43934 6862 43986 6914
rect 44158 6862 44210 6914
rect 45278 6862 45330 6914
rect 45502 6862 45554 6914
rect 3278 6750 3330 6802
rect 4958 6750 5010 6802
rect 5630 6750 5682 6802
rect 5742 6750 5794 6802
rect 6414 6750 6466 6802
rect 11006 6750 11058 6802
rect 12574 6750 12626 6802
rect 15598 6750 15650 6802
rect 19182 6750 19234 6802
rect 19854 6750 19906 6802
rect 23214 6750 23266 6802
rect 24670 6750 24722 6802
rect 26798 6750 26850 6802
rect 29150 6750 29202 6802
rect 44942 6750 44994 6802
rect 45054 6750 45106 6802
rect 3614 6638 3666 6690
rect 4174 6638 4226 6690
rect 4398 6638 4450 6690
rect 5070 6638 5122 6690
rect 5966 6638 6018 6690
rect 6190 6638 6242 6690
rect 6862 6638 6914 6690
rect 7310 6638 7362 6690
rect 7870 6638 7922 6690
rect 8206 6638 8258 6690
rect 15374 6638 15426 6690
rect 16382 6638 16434 6690
rect 17054 6638 17106 6690
rect 19630 6638 19682 6690
rect 20190 6638 20242 6690
rect 21870 6638 21922 6690
rect 23998 6638 24050 6690
rect 28142 6638 28194 6690
rect 28366 6638 28418 6690
rect 31950 6638 32002 6690
rect 32734 6638 32786 6690
rect 36206 6638 36258 6690
rect 39454 6638 39506 6690
rect 40462 6638 40514 6690
rect 40686 6638 40738 6690
rect 40910 6638 40962 6690
rect 41918 6638 41970 6690
rect 42814 6638 42866 6690
rect 45614 6638 45666 6690
rect 6638 6526 6690 6578
rect 8878 6526 8930 6578
rect 12014 6526 12066 6578
rect 12686 6526 12738 6578
rect 14254 6526 14306 6578
rect 15710 6526 15762 6578
rect 21310 6526 21362 6578
rect 21534 6526 21586 6578
rect 22878 6526 22930 6578
rect 28590 6526 28642 6578
rect 31278 6526 31330 6578
rect 35646 6526 35698 6578
rect 36430 6526 36482 6578
rect 37774 6526 37826 6578
rect 40014 6526 40066 6578
rect 40238 6526 40290 6578
rect 42142 6526 42194 6578
rect 42926 6526 42978 6578
rect 4846 6414 4898 6466
rect 7198 6414 7250 6466
rect 7422 6414 7474 6466
rect 11566 6414 11618 6466
rect 12126 6414 12178 6466
rect 13582 6414 13634 6466
rect 13918 6414 13970 6466
rect 14478 6414 14530 6466
rect 14590 6414 14642 6466
rect 14702 6414 14754 6466
rect 14814 6414 14866 6466
rect 15486 6414 15538 6466
rect 15822 6414 15874 6466
rect 19742 6414 19794 6466
rect 19966 6414 20018 6466
rect 20750 6414 20802 6466
rect 21758 6414 21810 6466
rect 23550 6414 23602 6466
rect 33742 6414 33794 6466
rect 35758 6414 35810 6466
rect 40798 6414 40850 6466
rect 44046 6414 44098 6466
rect 46062 6414 46114 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 6190 6078 6242 6130
rect 8542 6078 8594 6130
rect 15262 6078 15314 6130
rect 15374 6078 15426 6130
rect 15598 6078 15650 6130
rect 16382 6078 16434 6130
rect 17726 6078 17778 6130
rect 18062 6078 18114 6130
rect 18622 6078 18674 6130
rect 26238 6078 26290 6130
rect 33294 6078 33346 6130
rect 33518 6078 33570 6130
rect 40238 6078 40290 6130
rect 41022 6078 41074 6130
rect 41134 6078 41186 6130
rect 41246 6078 41298 6130
rect 2494 5966 2546 6018
rect 9102 5966 9154 6018
rect 15822 5966 15874 6018
rect 21646 5966 21698 6018
rect 25566 5966 25618 6018
rect 27358 5966 27410 6018
rect 33742 5966 33794 6018
rect 40350 5966 40402 6018
rect 42254 5966 42306 6018
rect 42366 5966 42418 6018
rect 45390 5966 45442 6018
rect 1822 5854 1874 5906
rect 4958 5854 5010 5906
rect 5182 5854 5234 5906
rect 5966 5854 6018 5906
rect 7086 5854 7138 5906
rect 7198 5854 7250 5906
rect 7310 5854 7362 5906
rect 7534 5854 7586 5906
rect 7982 5854 8034 5906
rect 8206 5854 8258 5906
rect 10110 5854 10162 5906
rect 16158 5854 16210 5906
rect 16606 5854 16658 5906
rect 16718 5854 16770 5906
rect 18398 5854 18450 5906
rect 18846 5854 18898 5906
rect 18958 5854 19010 5906
rect 23662 5854 23714 5906
rect 25230 5854 25282 5906
rect 26574 5854 26626 5906
rect 31166 5854 31218 5906
rect 33182 5854 33234 5906
rect 39566 5854 39618 5906
rect 40014 5854 40066 5906
rect 41470 5854 41522 5906
rect 41694 5854 41746 5906
rect 42142 5854 42194 5906
rect 46174 5854 46226 5906
rect 4622 5742 4674 5794
rect 13134 5742 13186 5794
rect 15374 5742 15426 5794
rect 16494 5742 16546 5794
rect 18734 5742 18786 5794
rect 33406 5742 33458 5794
rect 34638 5742 34690 5794
rect 42814 5742 42866 5794
rect 43262 5742 43314 5794
rect 5518 5630 5570 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 9662 5294 9714 5346
rect 25678 5294 25730 5346
rect 26350 5294 26402 5346
rect 26798 5294 26850 5346
rect 29150 5294 29202 5346
rect 29486 5294 29538 5346
rect 30046 5294 30098 5346
rect 30382 5294 30434 5346
rect 40798 5294 40850 5346
rect 45390 5294 45442 5346
rect 8206 5182 8258 5234
rect 8542 5182 8594 5234
rect 9550 5182 9602 5234
rect 10782 5182 10834 5234
rect 12910 5182 12962 5234
rect 16942 5182 16994 5234
rect 19070 5182 19122 5234
rect 22094 5182 22146 5234
rect 24222 5182 24274 5234
rect 24558 5182 24610 5234
rect 24782 5182 24834 5234
rect 26014 5182 26066 5234
rect 26462 5182 26514 5234
rect 27470 5182 27522 5234
rect 33854 5182 33906 5234
rect 34526 5182 34578 5234
rect 35422 5182 35474 5234
rect 36318 5182 36370 5234
rect 37774 5182 37826 5234
rect 39902 5182 39954 5234
rect 41022 5182 41074 5234
rect 41358 5182 41410 5234
rect 43486 5182 43538 5234
rect 44830 5182 44882 5234
rect 4846 5070 4898 5122
rect 5182 5070 5234 5122
rect 6078 5070 6130 5122
rect 6302 5070 6354 5122
rect 10110 5070 10162 5122
rect 15934 5070 15986 5122
rect 19854 5070 19906 5122
rect 20638 5070 20690 5122
rect 21422 5070 21474 5122
rect 25118 5070 25170 5122
rect 27582 5070 27634 5122
rect 27806 5070 27858 5122
rect 29710 5070 29762 5122
rect 30382 5070 30434 5122
rect 30942 5070 30994 5122
rect 34302 5070 34354 5122
rect 34414 5070 34466 5122
rect 34750 5070 34802 5122
rect 35198 5070 35250 5122
rect 36990 5070 37042 5122
rect 44270 5070 44322 5122
rect 45054 5070 45106 5122
rect 45950 5070 46002 5122
rect 4958 4958 5010 5010
rect 6974 4958 7026 5010
rect 9438 4958 9490 5010
rect 20414 4958 20466 5010
rect 25902 4958 25954 5010
rect 27022 4958 27074 5010
rect 31726 4958 31778 5010
rect 35646 4958 35698 5010
rect 35870 4958 35922 5010
rect 8990 4846 9042 4898
rect 15374 4846 15426 4898
rect 26910 4846 26962 4898
rect 34638 4846 34690 4898
rect 35422 4846 35474 4898
rect 36430 4846 36482 4898
rect 40462 4846 40514 4898
rect 45726 4846 45778 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 8654 4510 8706 4562
rect 17726 4510 17778 4562
rect 31838 4510 31890 4562
rect 32286 4510 32338 4562
rect 41022 4510 41074 4562
rect 7422 4398 7474 4450
rect 9662 4398 9714 4450
rect 10782 4398 10834 4450
rect 13582 4398 13634 4450
rect 14702 4398 14754 4450
rect 21982 4398 22034 4450
rect 24446 4398 24498 4450
rect 26014 4398 26066 4450
rect 31950 4398 32002 4450
rect 32398 4398 32450 4450
rect 33854 4398 33906 4450
rect 37102 4398 37154 4450
rect 40126 4398 40178 4450
rect 42478 4398 42530 4450
rect 45390 4398 45442 4450
rect 7086 4286 7138 4338
rect 7758 4286 7810 4338
rect 8430 4286 8482 4338
rect 10110 4286 10162 4338
rect 13246 4286 13298 4338
rect 14030 4286 14082 4338
rect 18062 4286 18114 4338
rect 21310 4286 21362 4338
rect 25230 4286 25282 4338
rect 28590 4286 28642 4338
rect 31614 4286 31666 4338
rect 33070 4286 33122 4338
rect 36318 4286 36370 4338
rect 40014 4286 40066 4338
rect 40350 4286 40402 4338
rect 40798 4286 40850 4338
rect 41134 4286 41186 4338
rect 42030 4286 42082 4338
rect 46174 4286 46226 4338
rect 4174 4174 4226 4226
rect 6302 4174 6354 4226
rect 7534 4174 7586 4226
rect 12910 4174 12962 4226
rect 13358 4174 13410 4226
rect 16830 4174 16882 4226
rect 18734 4174 18786 4226
rect 20862 4174 20914 4226
rect 24110 4174 24162 4226
rect 28142 4174 28194 4226
rect 29262 4174 29314 4226
rect 31390 4174 31442 4226
rect 35982 4174 36034 4226
rect 39230 4174 39282 4226
rect 41582 4174 41634 4226
rect 42814 4174 42866 4226
rect 43262 4174 43314 4226
rect 39566 4062 39618 4114
rect 42926 4062 42978 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 8766 3726 8818 3778
rect 23662 3726 23714 3778
rect 27470 3726 27522 3778
rect 38894 3726 38946 3778
rect 39230 3726 39282 3778
rect 44606 3726 44658 3778
rect 12574 3614 12626 3666
rect 13918 3614 13970 3666
rect 16046 3614 16098 3666
rect 18622 3614 18674 3666
rect 21870 3614 21922 3666
rect 23774 3614 23826 3666
rect 27582 3614 27634 3666
rect 29486 3614 29538 3666
rect 31614 3614 31666 3666
rect 36990 3614 37042 3666
rect 40126 3614 40178 3666
rect 42254 3614 42306 3666
rect 9774 3502 9826 3554
rect 13134 3502 13186 3554
rect 17278 3502 17330 3554
rect 17614 3502 17666 3554
rect 20974 3502 21026 3554
rect 23998 3502 24050 3554
rect 26686 3502 26738 3554
rect 28702 3502 28754 3554
rect 32174 3502 32226 3554
rect 35198 3502 35250 3554
rect 35982 3502 36034 3554
rect 43038 3502 43090 3554
rect 43710 3502 43762 3554
rect 8542 3390 8594 3442
rect 8654 3390 8706 3442
rect 10446 3390 10498 3442
rect 16942 3390 16994 3442
rect 26350 3390 26402 3442
rect 33742 3390 33794 3442
rect 35422 3390 35474 3442
rect 39118 3390 39170 3442
rect 2942 3278 2994 3330
rect 4510 3278 4562 3330
rect 6078 3278 6130 3330
rect 7534 3278 7586 3330
rect 8094 3278 8146 3330
rect 24894 3278 24946 3330
rect 25342 3278 25394 3330
rect 26014 3278 26066 3330
rect 27022 3278 27074 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 6048 47200 6160 48000
rect 17920 47200 18032 48000
rect 29792 47200 29904 48000
rect 41664 47200 41776 48000
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 6076 43708 6132 47200
rect 17948 45220 18004 47200
rect 17948 45164 18228 45220
rect 13580 44882 13636 44894
rect 13580 44830 13582 44882
rect 13634 44830 13636 44882
rect 10108 44436 10164 44446
rect 13580 44436 13636 44830
rect 14476 44882 14532 44894
rect 14476 44830 14478 44882
rect 14530 44830 14532 44882
rect 10108 44434 10724 44436
rect 10108 44382 10110 44434
rect 10162 44382 10724 44434
rect 10108 44380 10724 44382
rect 10108 44370 10164 44380
rect 9772 44210 9828 44222
rect 9772 44158 9774 44210
rect 9826 44158 9828 44210
rect 9548 44098 9604 44110
rect 9548 44046 9550 44098
rect 9602 44046 9604 44098
rect 9548 43876 9604 44046
rect 9212 43820 9548 43876
rect 8876 43764 8932 43774
rect 9212 43764 9268 43820
rect 9548 43810 9604 43820
rect 8876 43762 9268 43764
rect 8876 43710 8878 43762
rect 8930 43710 9268 43762
rect 8876 43708 9268 43710
rect 6076 43652 6244 43708
rect 8876 43698 8932 43708
rect 5964 43538 6020 43550
rect 5964 43486 5966 43538
rect 6018 43486 6020 43538
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5964 41972 6020 43486
rect 5964 41970 6132 41972
rect 5964 41918 5966 41970
rect 6018 41918 6132 41970
rect 5964 41916 6132 41918
rect 5964 41906 6020 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 6076 41188 6132 41916
rect 6076 40402 6132 41132
rect 6076 40350 6078 40402
rect 6130 40350 6132 40402
rect 6076 40338 6132 40350
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4620 39730 4676 39742
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 1820 39618 1876 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 37268 1876 39566
rect 2492 39508 2548 39518
rect 2492 39506 2772 39508
rect 2492 39454 2494 39506
rect 2546 39454 2772 39506
rect 2492 39452 2772 39454
rect 2492 39442 2548 39452
rect 2716 38722 2772 39452
rect 4620 39172 4676 39678
rect 4060 39116 4676 39172
rect 6076 39284 6132 39294
rect 2828 38948 2884 38958
rect 2828 38854 2884 38892
rect 3500 38948 3556 38958
rect 3500 38854 3556 38892
rect 3724 38834 3780 38846
rect 3724 38782 3726 38834
rect 3778 38782 3780 38834
rect 2716 38670 2718 38722
rect 2770 38670 2772 38722
rect 2716 38658 2772 38670
rect 3052 38724 3108 38734
rect 3052 38630 3108 38668
rect 3388 38612 3444 38622
rect 3388 38610 3556 38612
rect 3388 38558 3390 38610
rect 3442 38558 3556 38610
rect 3388 38556 3556 38558
rect 3388 38546 3444 38556
rect 1708 37156 1764 37166
rect 1708 37062 1764 37100
rect 1820 35698 1876 37212
rect 3388 38050 3444 38062
rect 3388 37998 3390 38050
rect 3442 37998 3444 38050
rect 3388 37156 3444 37998
rect 3388 37090 3444 37100
rect 3500 37940 3556 38556
rect 3724 38500 3780 38782
rect 3948 38834 4004 38846
rect 3948 38782 3950 38834
rect 4002 38782 4004 38834
rect 3948 38724 4004 38782
rect 3948 38658 4004 38668
rect 4060 38500 4116 39116
rect 4172 39004 4900 39060
rect 4172 38946 4228 39004
rect 4172 38894 4174 38946
rect 4226 38894 4228 38946
rect 4172 38882 4228 38894
rect 3724 38444 4116 38500
rect 3612 38276 3668 38286
rect 3612 38162 3668 38220
rect 3612 38110 3614 38162
rect 3666 38110 3668 38162
rect 3612 38098 3668 38110
rect 3948 37940 4004 37950
rect 2828 36484 2884 36494
rect 2828 36390 2884 36428
rect 3052 36482 3108 36494
rect 3276 36484 3332 36494
rect 3052 36430 3054 36482
rect 3106 36430 3108 36482
rect 2716 36372 2772 36382
rect 2492 36370 2772 36372
rect 2492 36318 2718 36370
rect 2770 36318 2772 36370
rect 2492 36316 2772 36318
rect 2492 35810 2548 36316
rect 2716 36306 2772 36316
rect 2492 35758 2494 35810
rect 2546 35758 2548 35810
rect 2492 35746 2548 35758
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35634 1876 35646
rect 3052 35026 3108 36430
rect 3052 34974 3054 35026
rect 3106 34974 3108 35026
rect 3052 34962 3108 34974
rect 3164 36428 3276 36484
rect 2828 34916 2884 34926
rect 2828 34580 2884 34860
rect 2940 34804 2996 34814
rect 2940 34802 3108 34804
rect 2940 34750 2942 34802
rect 2994 34750 3108 34802
rect 2940 34748 3108 34750
rect 2940 34738 2996 34748
rect 2828 34524 2996 34580
rect 2828 34356 2884 34366
rect 1932 34354 2884 34356
rect 1932 34302 2830 34354
rect 2882 34302 2884 34354
rect 1932 34300 2884 34302
rect 1932 34130 1988 34300
rect 2828 34290 2884 34300
rect 2940 34354 2996 34524
rect 2940 34302 2942 34354
rect 2994 34302 2996 34354
rect 1932 34078 1934 34130
rect 1986 34078 1988 34130
rect 1932 34066 1988 34078
rect 2156 34130 2212 34142
rect 2156 34078 2158 34130
rect 2210 34078 2212 34130
rect 2156 34020 2212 34078
rect 2492 34132 2548 34142
rect 2716 34132 2772 34142
rect 2492 34130 2716 34132
rect 2492 34078 2494 34130
rect 2546 34078 2716 34130
rect 2492 34076 2716 34078
rect 2492 34066 2548 34076
rect 2716 34038 2772 34076
rect 2156 33954 2212 33964
rect 2268 34018 2324 34030
rect 2268 33966 2270 34018
rect 2322 33966 2324 34018
rect 2268 33572 2324 33966
rect 2940 34020 2996 34302
rect 3052 34132 3108 34748
rect 3164 34580 3220 36428
rect 3276 36390 3332 36428
rect 3388 36484 3444 36494
rect 3500 36484 3556 37884
rect 3836 37938 4004 37940
rect 3836 37886 3950 37938
rect 4002 37886 4004 37938
rect 3836 37884 4004 37886
rect 3836 37380 3892 37884
rect 3948 37874 4004 37884
rect 4060 37492 4116 38444
rect 4284 38834 4340 38846
rect 4284 38782 4286 38834
rect 4338 38782 4340 38834
rect 4284 38276 4340 38782
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4396 38276 4452 38286
rect 4340 38274 4452 38276
rect 4340 38222 4398 38274
rect 4450 38222 4452 38274
rect 4340 38220 4452 38222
rect 4284 38210 4340 38220
rect 4396 38210 4452 38220
rect 4284 38050 4340 38062
rect 4284 37998 4286 38050
rect 4338 37998 4340 38050
rect 4172 37940 4228 37950
rect 4284 37940 4340 37998
rect 4228 37884 4340 37940
rect 4172 37874 4228 37884
rect 4396 37826 4452 37838
rect 4396 37774 4398 37826
rect 4450 37774 4452 37826
rect 4396 37492 4452 37774
rect 4060 37436 4452 37492
rect 3612 37324 3892 37380
rect 3612 36706 3668 37324
rect 3612 36654 3614 36706
rect 3666 36654 3668 36706
rect 3612 36642 3668 36654
rect 3836 37154 3892 37166
rect 3836 37102 3838 37154
rect 3890 37102 3892 37154
rect 3836 36594 3892 37102
rect 3836 36542 3838 36594
rect 3890 36542 3892 36594
rect 3836 36530 3892 36542
rect 3948 37156 4004 37166
rect 3444 36428 3556 36484
rect 3388 36418 3444 36428
rect 3836 36260 3892 36270
rect 3836 35812 3892 36204
rect 3836 35746 3892 35756
rect 3276 34916 3332 34926
rect 3276 34822 3332 34860
rect 3948 34914 4004 37100
rect 3948 34862 3950 34914
rect 4002 34862 4004 34914
rect 3948 34850 4004 34862
rect 4060 34916 4116 34926
rect 4172 34916 4228 37436
rect 4620 37268 4676 37278
rect 4620 37174 4676 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4732 36258 4788 36270
rect 4732 36206 4734 36258
rect 4786 36206 4788 36258
rect 4732 35812 4788 36206
rect 4844 36260 4900 39004
rect 6076 38946 6132 39228
rect 6076 38894 6078 38946
rect 6130 38894 6132 38946
rect 6076 38882 6132 38894
rect 5068 38836 5124 38846
rect 5068 37490 5124 38780
rect 5292 38834 5348 38846
rect 5292 38782 5294 38834
rect 5346 38782 5348 38834
rect 5292 38668 5348 38782
rect 6188 38668 6244 43652
rect 6636 43426 6692 43438
rect 6636 43374 6638 43426
rect 6690 43374 6692 43426
rect 6636 42980 6692 43374
rect 6636 42914 6692 42924
rect 9212 42866 9268 43708
rect 9772 43708 9828 44158
rect 9996 44100 10052 44110
rect 9996 44098 10164 44100
rect 9996 44046 9998 44098
rect 10050 44046 10164 44098
rect 9996 44044 10164 44046
rect 9996 44034 10052 44044
rect 10108 43876 10164 44044
rect 9772 43652 9940 43708
rect 9548 43316 9604 43326
rect 9212 42814 9214 42866
rect 9266 42814 9268 42866
rect 9212 42802 9268 42814
rect 9436 43314 9604 43316
rect 9436 43262 9550 43314
rect 9602 43262 9604 43314
rect 9436 43260 9604 43262
rect 6636 42644 6692 42654
rect 6636 41970 6692 42588
rect 6636 41918 6638 41970
rect 6690 41918 6692 41970
rect 6636 41906 6692 41918
rect 9324 42084 9380 42094
rect 9436 42084 9492 43260
rect 9548 43250 9604 43260
rect 9884 43316 9940 43652
rect 10108 43538 10164 43820
rect 10108 43486 10110 43538
rect 10162 43486 10164 43538
rect 10108 43474 10164 43486
rect 9884 43314 10164 43316
rect 9884 43262 9886 43314
rect 9938 43262 10164 43314
rect 9884 43260 10164 43262
rect 9884 43250 9940 43260
rect 10108 43092 10164 43260
rect 10108 43026 10164 43036
rect 9996 42980 10052 42990
rect 9772 42978 10052 42980
rect 9772 42926 9998 42978
rect 10050 42926 10052 42978
rect 9772 42924 10052 42926
rect 9660 42756 9716 42766
rect 9660 42662 9716 42700
rect 9548 42644 9604 42654
rect 9548 42550 9604 42588
rect 9380 42028 9492 42084
rect 8764 41858 8820 41870
rect 8764 41806 8766 41858
rect 8818 41806 8820 41858
rect 8764 41188 8820 41806
rect 9324 41410 9380 42028
rect 9324 41358 9326 41410
rect 9378 41358 9380 41410
rect 9324 41346 9380 41358
rect 9660 41412 9716 41422
rect 9772 41412 9828 42924
rect 9996 42914 10052 42924
rect 10668 42978 10724 44380
rect 13580 44380 13972 44436
rect 13580 44322 13636 44380
rect 13580 44270 13582 44322
rect 13634 44270 13636 44322
rect 11900 44100 11956 44110
rect 10668 42926 10670 42978
rect 10722 42926 10724 42978
rect 10668 42914 10724 42926
rect 10780 43538 10836 43550
rect 10780 43486 10782 43538
rect 10834 43486 10836 43538
rect 9884 42754 9940 42766
rect 9884 42702 9886 42754
rect 9938 42702 9940 42754
rect 9884 42084 9940 42702
rect 10556 42754 10612 42766
rect 10556 42702 10558 42754
rect 10610 42702 10612 42754
rect 10556 42084 10612 42702
rect 9884 42028 10276 42084
rect 9660 41410 9828 41412
rect 9660 41358 9662 41410
rect 9714 41358 9828 41410
rect 9660 41356 9828 41358
rect 9660 41346 9716 41356
rect 9100 41188 9156 41198
rect 8764 41186 9156 41188
rect 8764 41134 9102 41186
rect 9154 41134 9156 41186
rect 8764 41132 9156 41134
rect 9100 40404 9156 41132
rect 9100 40338 9156 40348
rect 9772 40402 9828 41356
rect 10108 41858 10164 41870
rect 10108 41806 10110 41858
rect 10162 41806 10164 41858
rect 10108 41188 10164 41806
rect 9772 40350 9774 40402
rect 9826 40350 9828 40402
rect 6860 40290 6916 40302
rect 6860 40238 6862 40290
rect 6914 40238 6916 40290
rect 6860 39844 6916 40238
rect 6860 39778 6916 39788
rect 8988 40290 9044 40302
rect 8988 40238 8990 40290
rect 9042 40238 9044 40290
rect 8092 39620 8148 39630
rect 8316 39620 8372 39630
rect 8092 39618 8372 39620
rect 8092 39566 8094 39618
rect 8146 39566 8318 39618
rect 8370 39566 8372 39618
rect 8092 39564 8372 39566
rect 8092 39554 8148 39564
rect 8316 39554 8372 39564
rect 7756 39506 7812 39518
rect 7756 39454 7758 39506
rect 7810 39454 7812 39506
rect 7084 39396 7140 39406
rect 7084 39302 7140 39340
rect 7420 39394 7476 39406
rect 7420 39342 7422 39394
rect 7474 39342 7476 39394
rect 5292 38612 5908 38668
rect 5852 37938 5908 38612
rect 5852 37886 5854 37938
rect 5906 37886 5908 37938
rect 5068 37438 5070 37490
rect 5122 37438 5124 37490
rect 5068 37426 5124 37438
rect 5180 37492 5236 37502
rect 5180 37398 5236 37436
rect 5740 37268 5796 37278
rect 5852 37268 5908 37886
rect 5796 37212 5908 37268
rect 6076 38612 6244 38668
rect 6412 38948 6468 38958
rect 5740 37174 5796 37212
rect 4956 37044 5012 37054
rect 4956 36482 5012 36988
rect 4956 36430 4958 36482
rect 5010 36430 5012 36482
rect 4956 36418 5012 36430
rect 5628 36594 5684 36606
rect 5628 36542 5630 36594
rect 5682 36542 5684 36594
rect 4844 36204 5012 36260
rect 4732 35746 4788 35756
rect 4620 35588 4676 35598
rect 4060 34914 4228 34916
rect 4060 34862 4062 34914
rect 4114 34862 4228 34914
rect 4060 34860 4228 34862
rect 4284 35586 4676 35588
rect 4284 35534 4622 35586
rect 4674 35534 4676 35586
rect 4284 35532 4676 35534
rect 4060 34850 4116 34860
rect 3500 34802 3556 34814
rect 3500 34750 3502 34802
rect 3554 34750 3556 34802
rect 3500 34692 3556 34750
rect 4284 34802 4340 35532
rect 4620 35522 4676 35532
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4844 35028 4900 35038
rect 4844 34934 4900 34972
rect 4396 34916 4452 34926
rect 4396 34822 4452 34860
rect 4284 34750 4286 34802
rect 4338 34750 4340 34802
rect 4284 34692 4340 34750
rect 3500 34636 4676 34692
rect 3164 34524 4004 34580
rect 3948 34354 4004 34524
rect 3948 34302 3950 34354
rect 4002 34302 4004 34354
rect 3948 34290 4004 34302
rect 4396 34244 4452 34254
rect 4396 34150 4452 34188
rect 4620 34242 4676 34636
rect 4620 34190 4622 34242
rect 4674 34190 4676 34242
rect 4620 34178 4676 34190
rect 3052 34066 3108 34076
rect 3276 34130 3332 34142
rect 3276 34078 3278 34130
rect 3330 34078 3332 34130
rect 3276 34020 3332 34078
rect 4508 34132 4564 34142
rect 4508 34038 4564 34076
rect 3388 34020 3444 34030
rect 3276 33964 3388 34020
rect 2940 33954 2996 33964
rect 3388 33954 3444 33964
rect 4844 34020 4900 34030
rect 4956 34020 5012 36204
rect 5628 35700 5684 36542
rect 5852 36372 5908 36382
rect 5852 35922 5908 36316
rect 5852 35870 5854 35922
rect 5906 35870 5908 35922
rect 5852 35858 5908 35870
rect 5628 35634 5684 35644
rect 5740 35812 5796 35822
rect 5292 35586 5348 35598
rect 5292 35534 5294 35586
rect 5346 35534 5348 35586
rect 5180 35474 5236 35486
rect 5180 35422 5182 35474
rect 5234 35422 5236 35474
rect 5068 34916 5124 34926
rect 5068 34354 5124 34860
rect 5068 34302 5070 34354
rect 5122 34302 5124 34354
rect 5068 34290 5124 34302
rect 5180 34244 5236 35422
rect 5292 35252 5348 35534
rect 5292 35186 5348 35196
rect 5180 34178 5236 34188
rect 4900 33964 5012 34020
rect 5292 34132 5348 34142
rect 5740 34132 5796 35756
rect 5964 35588 6020 35598
rect 5964 35494 6020 35532
rect 6076 34244 6132 38612
rect 6412 37378 6468 38892
rect 7420 38052 7476 39342
rect 7756 39396 7812 39454
rect 7756 38724 7812 39340
rect 7868 39394 7924 39406
rect 7868 39342 7870 39394
rect 7922 39342 7924 39394
rect 7868 38724 7924 39342
rect 8652 39394 8708 39406
rect 8652 39342 8654 39394
rect 8706 39342 8708 39394
rect 8652 39060 8708 39342
rect 8764 39396 8820 39406
rect 8764 39302 8820 39340
rect 8876 39394 8932 39406
rect 8876 39342 8878 39394
rect 8930 39342 8932 39394
rect 8652 39004 8820 39060
rect 8652 38836 8708 38846
rect 8652 38742 8708 38780
rect 8204 38724 8260 38734
rect 7868 38722 8260 38724
rect 7868 38670 8206 38722
rect 8258 38670 8260 38722
rect 7868 38668 8260 38670
rect 7756 38658 7812 38668
rect 7420 37986 7476 37996
rect 6412 37326 6414 37378
rect 6466 37326 6468 37378
rect 6412 37314 6468 37326
rect 8204 37380 8260 38668
rect 8764 37604 8820 39004
rect 8876 38948 8932 39342
rect 8988 39396 9044 40238
rect 9660 39620 9716 39630
rect 9772 39620 9828 40350
rect 9660 39618 9828 39620
rect 9660 39566 9662 39618
rect 9714 39566 9828 39618
rect 9660 39564 9828 39566
rect 9884 41132 10108 41188
rect 9660 39554 9716 39564
rect 8988 39330 9044 39340
rect 9436 39394 9492 39406
rect 9436 39342 9438 39394
rect 9490 39342 9492 39394
rect 8988 38948 9044 38958
rect 8876 38892 8988 38948
rect 8988 38854 9044 38892
rect 9436 38724 9492 39342
rect 9772 39396 9828 39406
rect 9772 39302 9828 39340
rect 9884 38834 9940 41132
rect 10108 41094 10164 41132
rect 10108 40402 10164 40414
rect 10108 40350 10110 40402
rect 10162 40350 10164 40402
rect 10108 39844 10164 40350
rect 10108 39778 10164 39788
rect 10220 39842 10276 42028
rect 10220 39790 10222 39842
rect 10274 39790 10276 39842
rect 10220 39778 10276 39790
rect 10332 40404 10388 40414
rect 10332 39506 10388 40348
rect 10556 39842 10612 42028
rect 10780 41300 10836 43486
rect 11452 43426 11508 43438
rect 11452 43374 11454 43426
rect 11506 43374 11508 43426
rect 11004 42980 11060 42990
rect 11004 42886 11060 42924
rect 11340 42980 11396 42990
rect 11452 42980 11508 43374
rect 11340 42978 11508 42980
rect 11340 42926 11342 42978
rect 11394 42926 11508 42978
rect 11340 42924 11508 42926
rect 11676 42980 11732 42990
rect 11340 42914 11396 42924
rect 11676 42886 11732 42924
rect 10892 42756 10948 42766
rect 10892 42662 10948 42700
rect 11452 42756 11508 42766
rect 11452 42662 11508 42700
rect 11900 42754 11956 44044
rect 13580 43426 13636 44270
rect 13580 43374 13582 43426
rect 13634 43374 13636 43426
rect 13580 43362 13636 43374
rect 13692 44210 13748 44222
rect 13692 44158 13694 44210
rect 13746 44158 13748 44210
rect 13468 42980 13524 42990
rect 13468 42886 13524 42924
rect 11900 42702 11902 42754
rect 11954 42702 11956 42754
rect 11900 42690 11956 42702
rect 12460 42756 12516 42766
rect 10668 41244 10836 41300
rect 10668 41188 10724 41244
rect 10668 41122 10724 41132
rect 11788 41188 11844 41198
rect 10780 41076 10836 41086
rect 11452 41076 11508 41086
rect 10780 41074 11172 41076
rect 10780 41022 10782 41074
rect 10834 41022 11172 41074
rect 10780 41020 11172 41022
rect 10780 41010 10836 41020
rect 10668 40292 10724 40302
rect 10668 40290 11060 40292
rect 10668 40238 10670 40290
rect 10722 40238 11060 40290
rect 10668 40236 11060 40238
rect 10668 40226 10724 40236
rect 10556 39790 10558 39842
rect 10610 39790 10612 39842
rect 10556 39778 10612 39790
rect 11004 39842 11060 40236
rect 11116 40290 11172 41020
rect 11116 40238 11118 40290
rect 11170 40238 11172 40290
rect 11116 40226 11172 40238
rect 11228 40514 11284 40526
rect 11228 40462 11230 40514
rect 11282 40462 11284 40514
rect 11004 39790 11006 39842
rect 11058 39790 11060 39842
rect 11004 39778 11060 39790
rect 11116 39732 11172 39742
rect 11116 39638 11172 39676
rect 10332 39454 10334 39506
rect 10386 39454 10388 39506
rect 10332 39442 10388 39454
rect 11228 39508 11284 40462
rect 11452 40290 11508 41020
rect 11788 40402 11844 41132
rect 11788 40350 11790 40402
rect 11842 40350 11844 40402
rect 11788 40338 11844 40350
rect 11452 40238 11454 40290
rect 11506 40238 11508 40290
rect 11452 40226 11508 40238
rect 11788 39844 11844 39854
rect 11788 39750 11844 39788
rect 11900 39618 11956 39630
rect 11900 39566 11902 39618
rect 11954 39566 11956 39618
rect 11676 39508 11732 39518
rect 11228 39506 11676 39508
rect 11228 39454 11230 39506
rect 11282 39454 11676 39506
rect 11228 39452 11676 39454
rect 11228 39442 11284 39452
rect 9884 38782 9886 38834
rect 9938 38782 9940 38834
rect 9884 38770 9940 38782
rect 9996 39394 10052 39406
rect 9996 39342 9998 39394
rect 10050 39342 10052 39394
rect 9436 38658 9492 38668
rect 8764 37538 8820 37548
rect 9884 38500 9940 38510
rect 9884 38164 9940 38444
rect 9996 38276 10052 39342
rect 11676 39172 11732 39452
rect 11900 39396 11956 39566
rect 12460 39396 12516 42700
rect 12908 42644 12964 42654
rect 12796 42530 12852 42542
rect 12796 42478 12798 42530
rect 12850 42478 12852 42530
rect 12796 41300 12852 42478
rect 12796 41234 12852 41244
rect 12908 41298 12964 42588
rect 13692 42644 13748 44158
rect 13804 44100 13860 44110
rect 13804 44006 13860 44044
rect 13916 43204 13972 44380
rect 14476 44434 14532 44830
rect 14476 44382 14478 44434
rect 14530 44382 14532 44434
rect 14476 44370 14532 44382
rect 14588 44436 14644 44446
rect 14588 44342 14644 44380
rect 15596 44436 15652 44446
rect 15596 44342 15652 44380
rect 15820 44434 15876 44446
rect 15820 44382 15822 44434
rect 15874 44382 15876 44434
rect 14140 44324 14196 44334
rect 14140 44322 14420 44324
rect 14140 44270 14142 44322
rect 14194 44270 14420 44322
rect 14140 44268 14420 44270
rect 14140 44258 14196 44268
rect 14028 43540 14084 43550
rect 14028 43538 14308 43540
rect 14028 43486 14030 43538
rect 14082 43486 14308 43538
rect 14028 43484 14308 43486
rect 14028 43474 14084 43484
rect 13916 43148 14196 43204
rect 13916 42756 13972 42766
rect 13916 42662 13972 42700
rect 14140 42754 14196 43148
rect 14140 42702 14142 42754
rect 14194 42702 14196 42754
rect 14140 42690 14196 42702
rect 13692 42578 13748 42588
rect 14028 42644 14084 42654
rect 14028 42550 14084 42588
rect 12908 41246 12910 41298
rect 12962 41246 12964 41298
rect 12908 41234 12964 41246
rect 13692 41970 13748 41982
rect 13692 41918 13694 41970
rect 13746 41918 13748 41970
rect 13692 41860 13748 41918
rect 13692 40964 13748 41804
rect 14028 41076 14084 41086
rect 14028 40982 14084 41020
rect 13692 40962 13972 40964
rect 13692 40910 13694 40962
rect 13746 40910 13972 40962
rect 13692 40908 13972 40910
rect 13692 40898 13748 40908
rect 12572 40292 12628 40302
rect 12572 40198 12628 40236
rect 13468 40292 13524 40302
rect 13468 39842 13524 40236
rect 13468 39790 13470 39842
rect 13522 39790 13524 39842
rect 13468 39778 13524 39790
rect 12908 39620 12964 39630
rect 12908 39526 12964 39564
rect 13468 39618 13524 39630
rect 13468 39566 13470 39618
rect 13522 39566 13524 39618
rect 13468 39508 13524 39566
rect 13468 39442 13524 39452
rect 13804 39508 13860 39518
rect 13804 39414 13860 39452
rect 12572 39396 12628 39406
rect 12460 39394 12628 39396
rect 12460 39342 12574 39394
rect 12626 39342 12628 39394
rect 12460 39340 12628 39342
rect 11900 39330 11956 39340
rect 11676 39116 11844 39172
rect 10556 38724 10612 38734
rect 10556 38722 11396 38724
rect 10556 38670 10558 38722
rect 10610 38670 11396 38722
rect 10556 38668 11396 38670
rect 10556 38658 10612 38668
rect 9996 38210 10052 38220
rect 11116 38276 11172 38286
rect 8988 37492 9044 37502
rect 9044 37436 9156 37492
rect 8988 37398 9044 37436
rect 8204 37314 8260 37324
rect 8876 37380 8932 37390
rect 8876 37286 8932 37324
rect 8540 37154 8596 37166
rect 8540 37102 8542 37154
rect 8594 37102 8596 37154
rect 8540 36708 8596 37102
rect 8876 36708 8932 36718
rect 8428 36706 8932 36708
rect 8428 36654 8878 36706
rect 8930 36654 8932 36706
rect 8428 36652 8932 36654
rect 7756 36372 7812 36382
rect 7756 36278 7812 36316
rect 6972 36260 7028 36270
rect 6972 35924 7028 36204
rect 6972 35922 7140 35924
rect 6972 35870 6974 35922
rect 7026 35870 7140 35922
rect 6972 35868 7140 35870
rect 6972 35858 7028 35868
rect 6748 35700 6804 35710
rect 6748 35606 6804 35644
rect 6524 35586 6580 35598
rect 6524 35534 6526 35586
rect 6578 35534 6580 35586
rect 6300 35474 6356 35486
rect 6300 35422 6302 35474
rect 6354 35422 6356 35474
rect 6300 34916 6356 35422
rect 6524 35252 6580 35534
rect 6860 35588 6916 35598
rect 6860 35494 6916 35532
rect 6524 35186 6580 35196
rect 6524 35028 6580 35038
rect 6300 34850 6356 34860
rect 6412 34972 6524 35028
rect 6412 34692 6468 34972
rect 6524 34962 6580 34972
rect 7084 34804 7140 35868
rect 7868 35810 7924 35822
rect 7868 35758 7870 35810
rect 7922 35758 7924 35810
rect 7756 35698 7812 35710
rect 7756 35646 7758 35698
rect 7810 35646 7812 35698
rect 7644 35586 7700 35598
rect 7644 35534 7646 35586
rect 7698 35534 7700 35586
rect 7196 35252 7252 35262
rect 7196 35138 7252 35196
rect 7196 35086 7198 35138
rect 7250 35086 7252 35138
rect 7196 35074 7252 35086
rect 7644 34914 7700 35534
rect 7756 35028 7812 35646
rect 7868 35140 7924 35758
rect 8428 35698 8484 36652
rect 8876 36642 8932 36652
rect 8428 35646 8430 35698
rect 8482 35646 8484 35698
rect 8428 35634 8484 35646
rect 8540 36482 8596 36494
rect 8540 36430 8542 36482
rect 8594 36430 8596 36482
rect 8540 35588 8596 36430
rect 9100 36370 9156 37436
rect 9548 37380 9604 37390
rect 9548 37286 9604 37324
rect 9324 37268 9380 37278
rect 9100 36318 9102 36370
rect 9154 36318 9156 36370
rect 8988 36260 9044 36270
rect 8988 36166 9044 36204
rect 8988 35700 9044 35710
rect 9100 35700 9156 36318
rect 8988 35698 9156 35700
rect 8988 35646 8990 35698
rect 9042 35646 9156 35698
rect 8988 35644 9156 35646
rect 9212 37212 9324 37268
rect 8988 35634 9044 35644
rect 8876 35588 8932 35598
rect 8540 35532 8876 35588
rect 7868 35074 7924 35084
rect 8204 35252 8260 35262
rect 7756 34962 7812 34972
rect 8092 35026 8148 35038
rect 8092 34974 8094 35026
rect 8146 34974 8148 35026
rect 7644 34862 7646 34914
rect 7698 34862 7700 34914
rect 7644 34850 7700 34862
rect 7868 34916 7924 34926
rect 7868 34822 7924 34860
rect 7196 34804 7252 34814
rect 7084 34802 7252 34804
rect 7084 34750 7198 34802
rect 7250 34750 7252 34802
rect 7084 34748 7252 34750
rect 7196 34738 7252 34748
rect 7308 34804 7364 34814
rect 7308 34710 7364 34748
rect 5964 34188 6132 34244
rect 6300 34636 6468 34692
rect 6300 34242 6356 34636
rect 7868 34356 7924 34366
rect 7420 34354 7924 34356
rect 7420 34302 7870 34354
rect 7922 34302 7924 34354
rect 7420 34300 7924 34302
rect 6300 34190 6302 34242
rect 6354 34190 6356 34242
rect 5852 34132 5908 34142
rect 5740 34130 5908 34132
rect 5740 34078 5854 34130
rect 5906 34078 5908 34130
rect 5740 34076 5908 34078
rect 4844 33954 4900 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5292 33684 5348 34076
rect 5852 34066 5908 34076
rect 5292 33618 5348 33628
rect 4620 33572 4676 33582
rect 2268 33516 2548 33572
rect 2492 33458 2548 33516
rect 2492 33406 2494 33458
rect 2546 33406 2548 33458
rect 2492 33394 2548 33406
rect 4620 33458 4676 33516
rect 4620 33406 4622 33458
rect 4674 33406 4676 33458
rect 4620 33394 4676 33406
rect 1820 33346 1876 33358
rect 1820 33294 1822 33346
rect 1874 33294 1876 33346
rect 1820 31778 1876 33294
rect 5628 33346 5684 33358
rect 5628 33294 5630 33346
rect 5682 33294 5684 33346
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4620 31892 4676 31902
rect 4620 31798 4676 31836
rect 1820 31726 1822 31778
rect 1874 31726 1876 31778
rect 1708 30322 1764 30334
rect 1708 30270 1710 30322
rect 1762 30270 1764 30322
rect 1708 29540 1764 30270
rect 1820 29764 1876 31726
rect 2492 31666 2548 31678
rect 2492 31614 2494 31666
rect 2546 31614 2548 31666
rect 2492 29988 2548 31614
rect 5516 31556 5572 31566
rect 5516 31462 5572 31500
rect 5628 31106 5684 33294
rect 5964 32788 6020 34188
rect 6300 34178 6356 34190
rect 6860 34244 6916 34254
rect 6860 34150 6916 34188
rect 7420 34242 7476 34300
rect 7868 34290 7924 34300
rect 7420 34190 7422 34242
rect 7474 34190 7476 34242
rect 7420 34178 7476 34190
rect 6412 34132 6468 34142
rect 6412 34038 6468 34076
rect 6972 34132 7028 34142
rect 6972 34038 7028 34076
rect 7196 34130 7252 34142
rect 7196 34078 7198 34130
rect 7250 34078 7252 34130
rect 6076 34018 6132 34030
rect 6076 33966 6078 34018
rect 6130 33966 6132 34018
rect 6076 33572 6132 33966
rect 7196 33908 7252 34078
rect 7756 34132 7812 34142
rect 7756 34038 7812 34076
rect 7980 34130 8036 34142
rect 7980 34078 7982 34130
rect 8034 34078 8036 34130
rect 7980 33908 8036 34078
rect 8092 34132 8148 34974
rect 8092 34066 8148 34076
rect 8204 34242 8260 35196
rect 8764 35140 8820 35150
rect 8764 34914 8820 35084
rect 8764 34862 8766 34914
rect 8818 34862 8820 34914
rect 8764 34850 8820 34862
rect 8204 34190 8206 34242
rect 8258 34190 8260 34242
rect 8204 34020 8260 34190
rect 8204 33954 8260 33964
rect 7196 33852 8036 33908
rect 7532 33572 7588 33582
rect 6076 33516 6468 33572
rect 6412 33458 6468 33516
rect 6412 33406 6414 33458
rect 6466 33406 6468 33458
rect 6412 33394 6468 33406
rect 5964 32732 6132 32788
rect 5628 31054 5630 31106
rect 5682 31054 5684 31106
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5180 30548 5236 30558
rect 4396 30436 4452 30446
rect 2492 29922 2548 29932
rect 3164 30324 3220 30334
rect 1820 29698 1876 29708
rect 3164 29650 3220 30268
rect 3164 29598 3166 29650
rect 3218 29598 3220 29650
rect 3164 29586 3220 29598
rect 3276 30212 3332 30222
rect 2044 29540 2100 29550
rect 1708 29538 2100 29540
rect 1708 29486 2046 29538
rect 2098 29486 2100 29538
rect 1708 29484 2100 29486
rect 1820 29316 1876 29326
rect 1708 28754 1764 28766
rect 1708 28702 1710 28754
rect 1762 28702 1764 28754
rect 1708 28532 1764 28702
rect 1708 28466 1764 28476
rect 1820 27074 1876 29260
rect 1932 28420 1988 29484
rect 2044 29474 2100 29484
rect 2604 29538 2660 29550
rect 2604 29486 2606 29538
rect 2658 29486 2660 29538
rect 2156 29428 2212 29438
rect 2492 29428 2548 29438
rect 2156 29426 2548 29428
rect 2156 29374 2158 29426
rect 2210 29374 2494 29426
rect 2546 29374 2548 29426
rect 2156 29372 2548 29374
rect 2156 29362 2212 29372
rect 2044 29204 2100 29214
rect 2044 29110 2100 29148
rect 2044 28420 2100 28430
rect 1932 28364 2044 28420
rect 2044 28354 2100 28364
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 27010 1876 27022
rect 1708 25618 1764 25630
rect 1708 25566 1710 25618
rect 1762 25566 1764 25618
rect 1708 24948 1764 25566
rect 1708 24882 1764 24892
rect 2380 24724 2436 29372
rect 2492 29362 2548 29372
rect 2604 28532 2660 29486
rect 2604 27636 2660 28476
rect 2828 29426 2884 29438
rect 2828 29374 2830 29426
rect 2882 29374 2884 29426
rect 2828 27972 2884 29374
rect 3052 29428 3108 29438
rect 3052 29334 3108 29372
rect 3164 29204 3220 29214
rect 3276 29204 3332 30156
rect 3836 30100 3892 30110
rect 3836 30006 3892 30044
rect 4396 29538 4452 30380
rect 4620 30324 4676 30334
rect 4620 30212 4676 30268
rect 4620 30210 4900 30212
rect 4620 30158 4622 30210
rect 4674 30158 4900 30210
rect 4620 30156 4900 30158
rect 4620 30146 4676 30156
rect 4396 29486 4398 29538
rect 4450 29486 4452 29538
rect 4396 29474 4452 29486
rect 3724 29428 3780 29438
rect 3724 29334 3780 29372
rect 4844 29428 4900 30156
rect 3164 29202 3332 29204
rect 3164 29150 3166 29202
rect 3218 29150 3332 29202
rect 3164 29148 3332 29150
rect 3164 29138 3220 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28868 4900 29372
rect 4620 28812 4900 28868
rect 4620 28642 4676 28812
rect 4620 28590 4622 28642
rect 4674 28590 4676 28642
rect 4620 28578 4676 28590
rect 3836 28530 3892 28542
rect 3836 28478 3838 28530
rect 3890 28478 3892 28530
rect 3836 28082 3892 28478
rect 3836 28030 3838 28082
rect 3890 28030 3892 28082
rect 3836 28018 3892 28030
rect 4956 28420 5012 28430
rect 2828 27906 2884 27916
rect 3164 27972 3220 27982
rect 3500 27972 3556 27982
rect 3164 27970 3332 27972
rect 3164 27918 3166 27970
rect 3218 27918 3332 27970
rect 3164 27916 3332 27918
rect 3164 27906 3220 27916
rect 2604 27570 2660 27580
rect 3052 27858 3108 27870
rect 3052 27806 3054 27858
rect 3106 27806 3108 27858
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2492 26628 2548 26910
rect 2492 26562 2548 26572
rect 3052 26740 3108 27806
rect 3164 27634 3220 27646
rect 3164 27582 3166 27634
rect 3218 27582 3220 27634
rect 3164 26852 3220 27582
rect 3276 27636 3332 27916
rect 3500 27858 3556 27916
rect 3500 27806 3502 27858
rect 3554 27806 3556 27858
rect 3500 27794 3556 27806
rect 3948 27860 4004 27870
rect 3948 27766 4004 27804
rect 4172 27858 4228 27870
rect 4172 27806 4174 27858
rect 4226 27806 4228 27858
rect 3276 27570 3332 27580
rect 4172 27076 4228 27806
rect 4620 27860 4676 27870
rect 4620 27858 4900 27860
rect 4620 27806 4622 27858
rect 4674 27806 4900 27858
rect 4620 27804 4900 27806
rect 4620 27794 4676 27804
rect 4732 27636 4788 27674
rect 4732 27570 4788 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 27300 4900 27804
rect 4956 27858 5012 28364
rect 4956 27806 4958 27858
rect 5010 27806 5012 27858
rect 4956 27794 5012 27806
rect 5180 27858 5236 30492
rect 5628 30324 5684 31054
rect 5740 31892 5796 31902
rect 5740 31554 5796 31836
rect 5740 31502 5742 31554
rect 5794 31502 5796 31554
rect 5740 30548 5796 31502
rect 5852 31666 5908 31678
rect 5852 31614 5854 31666
rect 5906 31614 5908 31666
rect 5852 31444 5908 31614
rect 5852 31378 5908 31388
rect 5740 30482 5796 30492
rect 5628 30258 5684 30268
rect 5852 30212 5908 30222
rect 5852 30118 5908 30156
rect 5628 30098 5684 30110
rect 5628 30046 5630 30098
rect 5682 30046 5684 30098
rect 5516 29540 5572 29550
rect 5516 28980 5572 29484
rect 5628 29204 5684 30046
rect 5740 30100 5796 30110
rect 5740 30006 5796 30044
rect 5628 29138 5684 29148
rect 5516 28924 5684 28980
rect 5628 28530 5684 28924
rect 5628 28478 5630 28530
rect 5682 28478 5684 28530
rect 5628 28466 5684 28478
rect 5740 28420 5796 28430
rect 5740 28082 5796 28364
rect 5740 28030 5742 28082
rect 5794 28030 5796 28082
rect 5740 28018 5796 28030
rect 5964 28418 6020 28430
rect 5964 28366 5966 28418
rect 6018 28366 6020 28418
rect 5292 27972 5348 27982
rect 5292 27878 5348 27916
rect 5180 27806 5182 27858
rect 5234 27806 5236 27858
rect 5180 27794 5236 27806
rect 5516 27860 5572 27870
rect 5516 27766 5572 27804
rect 5852 27858 5908 27870
rect 5852 27806 5854 27858
rect 5906 27806 5908 27858
rect 3164 26786 3220 26796
rect 3724 27020 4228 27076
rect 3052 26402 3108 26684
rect 3164 26516 3220 26526
rect 3164 26422 3220 26460
rect 3052 26350 3054 26402
rect 3106 26350 3108 26402
rect 3052 26338 3108 26350
rect 3724 26290 3780 27020
rect 3836 26852 3892 26862
rect 3836 26402 3892 26796
rect 3948 26628 4004 26638
rect 3948 26514 4004 26572
rect 3948 26462 3950 26514
rect 4002 26462 4004 26514
rect 3948 26450 4004 26462
rect 3836 26350 3838 26402
rect 3890 26350 3892 26402
rect 3836 26338 3892 26350
rect 3724 26238 3726 26290
rect 3778 26238 3780 26290
rect 3724 26226 3780 26238
rect 3164 26066 3220 26078
rect 3164 26014 3166 26066
rect 3218 26014 3220 26066
rect 3164 25172 3220 26014
rect 3164 25106 3220 25116
rect 3836 25394 3892 25406
rect 3836 25342 3838 25394
rect 3890 25342 3892 25394
rect 3276 24948 3332 24958
rect 3276 24854 3332 24892
rect 3836 24946 3892 25342
rect 3836 24894 3838 24946
rect 3890 24894 3892 24946
rect 3836 24882 3892 24894
rect 3948 25172 4004 25182
rect 2380 24658 2436 24668
rect 3164 24724 3220 24734
rect 3164 24630 3220 24668
rect 3500 24724 3556 24734
rect 3724 24724 3780 24734
rect 3500 24722 3780 24724
rect 3500 24670 3502 24722
rect 3554 24670 3726 24722
rect 3778 24670 3780 24722
rect 3500 24668 3780 24670
rect 3500 24658 3556 24668
rect 3724 24658 3780 24668
rect 3948 24722 4004 25116
rect 3948 24670 3950 24722
rect 4002 24670 4004 24722
rect 3948 24658 4004 24670
rect 4172 24722 4228 27020
rect 4620 27244 4900 27300
rect 4620 27186 4676 27244
rect 4620 27134 4622 27186
rect 4674 27134 4676 27186
rect 4620 26516 4676 27134
rect 5852 26740 5908 27806
rect 4620 26422 4676 26460
rect 5628 26684 5852 26740
rect 4396 26402 4452 26414
rect 4396 26350 4398 26402
rect 4450 26350 4452 26402
rect 4284 26292 4340 26302
rect 4396 26292 4452 26350
rect 4284 26290 4452 26292
rect 4284 26238 4286 26290
rect 4338 26238 4452 26290
rect 4284 26236 4452 26238
rect 4732 26292 4788 26302
rect 4732 26290 4900 26292
rect 4732 26238 4734 26290
rect 4786 26238 4900 26290
rect 4732 26236 4900 26238
rect 4284 26226 4340 26236
rect 4732 26226 4788 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4508 25732 4564 25742
rect 4508 25506 4564 25676
rect 4508 25454 4510 25506
rect 4562 25454 4564 25506
rect 4508 25442 4564 25454
rect 4172 24670 4174 24722
rect 4226 24670 4228 24722
rect 3836 24500 3892 24510
rect 3836 23938 3892 24444
rect 3836 23886 3838 23938
rect 3890 23886 3892 23938
rect 3836 23874 3892 23886
rect 4060 23940 4116 23950
rect 4172 23940 4228 24670
rect 4620 24836 4676 24846
rect 4844 24836 4900 26236
rect 5628 25396 5684 26684
rect 5852 26674 5908 26684
rect 5964 27860 6020 28366
rect 5740 26292 5796 26302
rect 5740 25732 5796 26236
rect 5740 25666 5796 25676
rect 5516 25394 5684 25396
rect 5516 25342 5630 25394
rect 5682 25342 5684 25394
rect 5516 25340 5684 25342
rect 4956 24948 5012 24958
rect 5404 24948 5460 24958
rect 5012 24892 5124 24948
rect 4956 24882 5012 24892
rect 4620 24834 4900 24836
rect 4620 24782 4622 24834
rect 4674 24782 4900 24834
rect 4620 24780 4900 24782
rect 4620 24724 4676 24780
rect 4620 24658 4676 24668
rect 4956 24724 5012 24734
rect 4956 24630 5012 24668
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4060 23938 5012 23940
rect 4060 23886 4062 23938
rect 4114 23886 5012 23938
rect 4060 23884 5012 23886
rect 4060 23874 4116 23884
rect 3500 23826 3556 23838
rect 3500 23774 3502 23826
rect 3554 23774 3556 23826
rect 2492 23716 2548 23726
rect 2492 23266 2548 23660
rect 3500 23380 3556 23774
rect 3612 23716 3668 23726
rect 3612 23622 3668 23660
rect 4396 23714 4452 23726
rect 4396 23662 4398 23714
rect 4450 23662 4452 23714
rect 3500 23314 3556 23324
rect 2492 23214 2494 23266
rect 2546 23214 2548 23266
rect 2492 23202 2548 23214
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 21586 1876 23102
rect 4396 23156 4452 23662
rect 4732 23716 4788 23726
rect 4732 23622 4788 23660
rect 4956 23378 5012 23884
rect 4956 23326 4958 23378
rect 5010 23326 5012 23378
rect 4956 23314 5012 23326
rect 4396 23090 4452 23100
rect 4620 23268 4676 23278
rect 4620 23042 4676 23212
rect 5068 23156 5124 24892
rect 5404 24854 5460 24892
rect 5516 24834 5572 25340
rect 5628 25330 5684 25340
rect 5852 25508 5908 25518
rect 5964 25508 6020 27804
rect 5852 25506 6020 25508
rect 5852 25454 5854 25506
rect 5906 25454 6020 25506
rect 5852 25452 6020 25454
rect 5516 24782 5518 24834
rect 5570 24782 5572 24834
rect 5516 24770 5572 24782
rect 5404 24500 5460 24510
rect 5404 24406 5460 24444
rect 5740 23716 5796 23726
rect 5740 23622 5796 23660
rect 5852 23492 5908 25452
rect 6076 24388 6132 32732
rect 7532 32562 7588 33516
rect 7532 32510 7534 32562
rect 7586 32510 7588 32562
rect 7532 32498 7588 32510
rect 7980 32452 8036 33852
rect 8540 33458 8596 33470
rect 8540 33406 8542 33458
rect 8594 33406 8596 33458
rect 8540 32452 8596 33406
rect 7980 32450 8596 32452
rect 7980 32398 7982 32450
rect 8034 32398 8596 32450
rect 7980 32396 8596 32398
rect 7980 32386 8036 32396
rect 8764 32338 8820 32350
rect 8764 32286 8766 32338
rect 8818 32286 8820 32338
rect 7644 31780 7700 31790
rect 8428 31780 8484 31790
rect 6300 31666 6356 31678
rect 6300 31614 6302 31666
rect 6354 31614 6356 31666
rect 6188 31556 6244 31566
rect 6188 30772 6244 31500
rect 6300 31444 6356 31614
rect 6636 31668 6692 31678
rect 6860 31668 6916 31678
rect 6636 31666 6916 31668
rect 6636 31614 6638 31666
rect 6690 31614 6862 31666
rect 6914 31614 6916 31666
rect 6636 31612 6916 31614
rect 6636 31602 6692 31612
rect 6860 31602 6916 31612
rect 7196 31666 7252 31678
rect 7420 31668 7476 31678
rect 7196 31614 7198 31666
rect 7250 31614 7252 31666
rect 6412 31556 6468 31566
rect 6412 31554 6580 31556
rect 6412 31502 6414 31554
rect 6466 31502 6580 31554
rect 6412 31500 6580 31502
rect 6412 31490 6468 31500
rect 6300 31378 6356 31388
rect 6188 30716 6468 30772
rect 6188 30212 6244 30222
rect 6188 30118 6244 30156
rect 6412 30210 6468 30716
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 6524 29540 6580 31500
rect 6972 31554 7028 31566
rect 6972 31502 6974 31554
rect 7026 31502 7028 31554
rect 6972 30436 7028 31502
rect 7196 31220 7252 31614
rect 7196 31154 7252 31164
rect 7308 31612 7420 31668
rect 7308 30436 7364 31612
rect 7420 31574 7476 31612
rect 7644 30994 7700 31724
rect 8316 31724 8428 31780
rect 7644 30942 7646 30994
rect 7698 30942 7700 30994
rect 7644 30930 7700 30942
rect 7756 31666 7812 31678
rect 7756 31614 7758 31666
rect 7810 31614 7812 31666
rect 7756 31444 7812 31614
rect 6972 30370 7028 30380
rect 7084 30380 7308 30436
rect 6748 30324 6804 30334
rect 6636 29988 6692 29998
rect 6636 29894 6692 29932
rect 6524 29316 6580 29484
rect 6748 29428 6804 30268
rect 7084 30212 7140 30380
rect 7308 30342 7364 30380
rect 7420 30324 7476 30334
rect 7420 30230 7476 30268
rect 7756 30212 7812 31388
rect 7868 31554 7924 31566
rect 8092 31556 8148 31566
rect 7868 31502 7870 31554
rect 7922 31502 7924 31554
rect 7868 31108 7924 31502
rect 7868 30324 7924 31052
rect 7868 30258 7924 30268
rect 7980 31554 8148 31556
rect 7980 31502 8094 31554
rect 8146 31502 8148 31554
rect 7980 31500 8148 31502
rect 7084 30118 7140 30156
rect 7532 30156 7812 30212
rect 6860 30098 6916 30110
rect 6860 30046 6862 30098
rect 6914 30046 6916 30098
rect 6860 29652 6916 30046
rect 6860 29586 6916 29596
rect 7420 29538 7476 29550
rect 7420 29486 7422 29538
rect 7474 29486 7476 29538
rect 7308 29428 7364 29438
rect 6748 29372 6916 29428
rect 6524 29314 6804 29316
rect 6524 29262 6526 29314
rect 6578 29262 6804 29314
rect 6524 29260 6804 29262
rect 6524 29250 6580 29260
rect 6636 28756 6692 28766
rect 6636 28662 6692 28700
rect 6412 28642 6468 28654
rect 6412 28590 6414 28642
rect 6466 28590 6468 28642
rect 6412 28196 6468 28590
rect 6748 28644 6804 29260
rect 6860 28866 6916 29372
rect 7308 29334 7364 29372
rect 6860 28814 6862 28866
rect 6914 28814 6916 28866
rect 6860 28802 6916 28814
rect 7420 28756 7476 29486
rect 7196 28700 7420 28756
rect 6972 28644 7028 28654
rect 6748 28642 7028 28644
rect 6748 28590 6974 28642
rect 7026 28590 7028 28642
rect 6748 28588 7028 28590
rect 6972 28578 7028 28588
rect 6412 28130 6468 28140
rect 6524 28418 6580 28430
rect 6524 28366 6526 28418
rect 6578 28366 6580 28418
rect 6300 28082 6356 28094
rect 6300 28030 6302 28082
rect 6354 28030 6356 28082
rect 6188 27972 6244 27982
rect 6300 27972 6356 28030
rect 6244 27916 6356 27972
rect 6412 27972 6468 27982
rect 6524 27972 6580 28366
rect 7196 28082 7252 28700
rect 7420 28662 7476 28700
rect 7532 28532 7588 30156
rect 7868 29540 7924 29550
rect 7980 29540 8036 31500
rect 8092 31490 8148 31500
rect 8092 31220 8148 31230
rect 8148 31164 8260 31220
rect 8092 31154 8148 31164
rect 8204 31106 8260 31164
rect 8204 31054 8206 31106
rect 8258 31054 8260 31106
rect 8204 31042 8260 31054
rect 8316 30436 8372 31724
rect 8428 31686 8484 31724
rect 8428 31108 8484 31118
rect 8428 31014 8484 31052
rect 8540 30994 8596 31006
rect 8540 30942 8542 30994
rect 8594 30942 8596 30994
rect 8204 30380 8372 30436
rect 8428 30436 8484 30446
rect 8092 30100 8148 30110
rect 8092 29650 8148 30044
rect 8092 29598 8094 29650
rect 8146 29598 8148 29650
rect 8092 29586 8148 29598
rect 7868 29538 8036 29540
rect 7868 29486 7870 29538
rect 7922 29486 8036 29538
rect 7868 29484 8036 29486
rect 7868 29474 7924 29484
rect 7644 29426 7700 29438
rect 7644 29374 7646 29426
rect 7698 29374 7700 29426
rect 7644 29092 7700 29374
rect 8092 29426 8148 29438
rect 8092 29374 8094 29426
rect 8146 29374 8148 29426
rect 8092 29092 8148 29374
rect 7644 29036 8148 29092
rect 7196 28030 7198 28082
rect 7250 28030 7252 28082
rect 7196 28018 7252 28030
rect 7308 28476 7588 28532
rect 6412 27970 6580 27972
rect 6412 27918 6414 27970
rect 6466 27918 6580 27970
rect 6412 27916 6580 27918
rect 6188 27906 6244 27916
rect 6412 27906 6468 27916
rect 7084 27860 7140 27870
rect 7308 27860 7364 28476
rect 7420 28364 7924 28420
rect 7420 28082 7476 28364
rect 7420 28030 7422 28082
rect 7474 28030 7476 28082
rect 7420 28018 7476 28030
rect 7756 28196 7812 28206
rect 7756 28082 7812 28140
rect 7756 28030 7758 28082
rect 7810 28030 7812 28082
rect 7084 27858 7364 27860
rect 7084 27806 7086 27858
rect 7138 27806 7364 27858
rect 7084 27804 7364 27806
rect 7644 27860 7700 27870
rect 7084 27794 7140 27804
rect 6300 27634 6356 27646
rect 6300 27582 6302 27634
rect 6354 27582 6356 27634
rect 6076 24322 6132 24332
rect 6188 24724 6244 24734
rect 6076 23940 6132 23950
rect 6188 23940 6244 24668
rect 6132 23884 6244 23940
rect 6076 23826 6132 23884
rect 6076 23774 6078 23826
rect 6130 23774 6132 23826
rect 6076 23762 6132 23774
rect 5628 23436 5908 23492
rect 5516 23380 5572 23390
rect 5516 23286 5572 23324
rect 4620 22990 4622 23042
rect 4674 22990 4676 23042
rect 4620 22932 4676 22990
rect 4284 22876 4676 22932
rect 4956 23100 5124 23156
rect 5292 23154 5348 23166
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 2828 22372 2884 22382
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 19234 1876 21534
rect 2716 21700 2772 21710
rect 2492 21476 2548 21486
rect 2492 21382 2548 21420
rect 2380 20804 2436 20814
rect 2716 20804 2772 21644
rect 2380 20802 2772 20804
rect 2380 20750 2382 20802
rect 2434 20750 2718 20802
rect 2770 20750 2772 20802
rect 2380 20748 2772 20750
rect 2380 20738 2436 20748
rect 2044 20580 2100 20590
rect 2268 20580 2324 20590
rect 2044 20578 2212 20580
rect 2044 20526 2046 20578
rect 2098 20526 2212 20578
rect 2044 20524 2212 20526
rect 2044 20514 2100 20524
rect 2044 20356 2100 20366
rect 2044 20130 2100 20300
rect 2156 20188 2212 20524
rect 2268 20486 2324 20524
rect 2604 20188 2660 20748
rect 2716 20738 2772 20748
rect 2828 20690 2884 22316
rect 4060 22370 4116 22382
rect 4060 22318 4062 22370
rect 4114 22318 4116 22370
rect 3388 22258 3444 22270
rect 3388 22206 3390 22258
rect 3442 22206 3444 22258
rect 2828 20638 2830 20690
rect 2882 20638 2884 20690
rect 2828 20626 2884 20638
rect 3052 20692 3108 20702
rect 3052 20598 3108 20636
rect 3276 20690 3332 20702
rect 3276 20638 3278 20690
rect 3330 20638 3332 20690
rect 3276 20356 3332 20638
rect 3276 20290 3332 20300
rect 2156 20132 2324 20188
rect 2604 20132 2772 20188
rect 2044 20078 2046 20130
rect 2098 20078 2100 20130
rect 2044 20066 2100 20078
rect 2268 20130 2324 20132
rect 2268 20078 2270 20130
rect 2322 20078 2324 20130
rect 2268 20066 2324 20078
rect 2604 20020 2660 20030
rect 2604 19926 2660 19964
rect 2492 19906 2548 19918
rect 2492 19854 2494 19906
rect 2546 19854 2548 19906
rect 2492 19346 2548 19854
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2492 19282 2548 19294
rect 1820 19182 1822 19234
rect 1874 19182 1876 19234
rect 1820 18564 1876 19182
rect 1820 18450 1876 18508
rect 1820 18398 1822 18450
rect 1874 18398 1876 18450
rect 1820 16882 1876 18398
rect 2492 19124 2548 19134
rect 2492 18450 2548 19068
rect 2492 18398 2494 18450
rect 2546 18398 2548 18450
rect 2492 18386 2548 18398
rect 2716 17666 2772 20132
rect 3388 20132 3444 22206
rect 4060 22260 4116 22318
rect 4284 22372 4340 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4732 22484 4788 22494
rect 4732 22390 4788 22428
rect 4396 22372 4452 22382
rect 4284 22316 4396 22372
rect 4396 22278 4452 22316
rect 3948 22148 4004 22158
rect 3612 21476 3668 21486
rect 3500 20692 3556 20702
rect 3500 20598 3556 20636
rect 3612 20578 3668 21420
rect 3948 20802 4004 22092
rect 3948 20750 3950 20802
rect 4002 20750 4004 20802
rect 3948 20738 4004 20750
rect 4060 21476 4116 22204
rect 4956 22258 5012 23100
rect 4956 22206 4958 22258
rect 5010 22206 5012 22258
rect 4956 22194 5012 22206
rect 5292 21812 5348 23102
rect 5516 22148 5572 22158
rect 5516 22054 5572 22092
rect 5292 21746 5348 21756
rect 4956 21700 5012 21710
rect 4956 21606 5012 21644
rect 5292 21588 5348 21598
rect 5628 21588 5684 23436
rect 5740 23268 5796 23278
rect 5740 23174 5796 23212
rect 5852 23156 5908 23166
rect 6300 23156 6356 27582
rect 7084 27076 7140 27086
rect 6748 27074 7140 27076
rect 6748 27022 7086 27074
rect 7138 27022 7140 27074
rect 6748 27020 7140 27022
rect 6412 26178 6468 26190
rect 6412 26126 6414 26178
rect 6466 26126 6468 26178
rect 6412 25730 6468 26126
rect 6412 25678 6414 25730
rect 6466 25678 6468 25730
rect 6412 25666 6468 25678
rect 6748 25620 6804 27020
rect 7084 27010 7140 27020
rect 7196 26908 7252 27804
rect 7644 27766 7700 27804
rect 6860 26852 7252 26908
rect 6860 26850 6916 26852
rect 6860 26798 6862 26850
rect 6914 26798 6916 26850
rect 6860 26786 6916 26798
rect 6636 25564 6804 25620
rect 6524 25282 6580 25294
rect 6524 25230 6526 25282
rect 6578 25230 6580 25282
rect 6524 25060 6580 25230
rect 6524 24994 6580 25004
rect 6524 24836 6580 24846
rect 6524 24742 6580 24780
rect 6636 24612 6692 25564
rect 6748 25396 6804 25406
rect 6748 25394 7364 25396
rect 6748 25342 6750 25394
rect 6802 25342 7364 25394
rect 6748 25340 7364 25342
rect 6748 25330 6804 25340
rect 7196 25172 7252 25182
rect 7084 25060 7140 25070
rect 6412 24556 6692 24612
rect 6748 24722 6804 24734
rect 6748 24670 6750 24722
rect 6802 24670 6804 24722
rect 6412 23826 6468 24556
rect 6748 24276 6804 24670
rect 6412 23774 6414 23826
rect 6466 23774 6468 23826
rect 6412 23604 6468 23774
rect 6412 23538 6468 23548
rect 6524 24220 6804 24276
rect 6524 23716 6580 24220
rect 7084 24164 7140 25004
rect 7196 24946 7252 25116
rect 7196 24894 7198 24946
rect 7250 24894 7252 24946
rect 7196 24882 7252 24894
rect 7308 24946 7364 25340
rect 7756 25284 7812 28030
rect 7868 28084 7924 28364
rect 7868 28028 8148 28084
rect 7980 27860 8036 27870
rect 7980 27766 8036 27804
rect 8092 27858 8148 28028
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 8092 27794 8148 27806
rect 8204 26908 8260 30380
rect 8428 29538 8484 30380
rect 8428 29486 8430 29538
rect 8482 29486 8484 29538
rect 8428 29474 8484 29486
rect 8540 29428 8596 30942
rect 8764 29764 8820 32286
rect 8876 31778 8932 35532
rect 9100 34356 9156 34366
rect 9212 34356 9268 37212
rect 9324 37202 9380 37212
rect 9884 37268 9940 38108
rect 10108 38052 10164 38062
rect 10108 37958 10164 37996
rect 11116 38050 11172 38220
rect 11340 38162 11396 38668
rect 11340 38110 11342 38162
rect 11394 38110 11396 38162
rect 11340 38098 11396 38110
rect 11564 38276 11620 38286
rect 11116 37998 11118 38050
rect 11170 37998 11172 38050
rect 11116 37986 11172 37998
rect 11564 38050 11620 38220
rect 11564 37998 11566 38050
rect 11618 37998 11620 38050
rect 11564 37986 11620 37998
rect 11788 38050 11844 39116
rect 11788 37998 11790 38050
rect 11842 37998 11844 38050
rect 11788 37986 11844 37998
rect 11900 38724 11956 38734
rect 12572 38668 12628 39340
rect 13132 39172 13188 39182
rect 13132 39058 13188 39116
rect 13132 39006 13134 39058
rect 13186 39006 13188 39058
rect 13020 38836 13076 38846
rect 11900 37940 11956 38668
rect 10892 37716 10948 37726
rect 9884 37174 9940 37212
rect 10444 37378 10500 37390
rect 10444 37326 10446 37378
rect 10498 37326 10500 37378
rect 10108 37156 10164 37166
rect 10444 37156 10500 37326
rect 10780 37268 10836 37278
rect 10892 37268 10948 37660
rect 10780 37266 10948 37268
rect 10780 37214 10782 37266
rect 10834 37214 10948 37266
rect 10780 37212 10948 37214
rect 10780 37202 10836 37212
rect 10108 37154 10500 37156
rect 10108 37102 10110 37154
rect 10162 37102 10500 37154
rect 10108 37100 10500 37102
rect 9660 36482 9716 36494
rect 9660 36430 9662 36482
rect 9714 36430 9716 36482
rect 9436 35700 9492 35710
rect 9100 34354 9268 34356
rect 9100 34302 9102 34354
rect 9154 34302 9268 34354
rect 9100 34300 9268 34302
rect 9324 34802 9380 34814
rect 9324 34750 9326 34802
rect 9378 34750 9380 34802
rect 9100 34290 9156 34300
rect 9324 33460 9380 34750
rect 9436 34130 9492 35644
rect 9660 35588 9716 36430
rect 9772 35588 9828 35598
rect 9660 35532 9772 35588
rect 9772 35494 9828 35532
rect 10108 35252 10164 37100
rect 10108 35186 10164 35196
rect 10332 36370 10388 36382
rect 10332 36318 10334 36370
rect 10386 36318 10388 36370
rect 9884 35140 9940 35150
rect 9660 35028 9716 35038
rect 9660 34244 9716 34972
rect 9884 34356 9940 35084
rect 9884 34262 9940 34300
rect 9996 34804 10052 34814
rect 9996 34354 10052 34748
rect 10332 34468 10388 36318
rect 10332 34402 10388 34412
rect 10780 34468 10836 34478
rect 9996 34302 9998 34354
rect 10050 34302 10052 34354
rect 9996 34290 10052 34302
rect 10444 34356 10500 34366
rect 10444 34262 10500 34300
rect 9660 34178 9716 34188
rect 9436 34078 9438 34130
rect 9490 34078 9492 34130
rect 9436 34066 9492 34078
rect 10108 34130 10164 34142
rect 10556 34132 10612 34142
rect 10108 34078 10110 34130
rect 10162 34078 10164 34130
rect 10108 33684 10164 34078
rect 9996 33628 10164 33684
rect 10220 34130 10612 34132
rect 10220 34078 10558 34130
rect 10610 34078 10612 34130
rect 10220 34076 10612 34078
rect 9436 33460 9492 33470
rect 9324 33458 9492 33460
rect 9324 33406 9438 33458
rect 9490 33406 9492 33458
rect 9324 33404 9492 33406
rect 9436 33394 9492 33404
rect 9996 33348 10052 33628
rect 9996 33254 10052 33292
rect 9548 32340 9604 32350
rect 9548 31890 9604 32284
rect 9548 31838 9550 31890
rect 9602 31838 9604 31890
rect 9548 31826 9604 31838
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 8876 31714 8932 31726
rect 9548 31668 9604 31678
rect 9548 31218 9604 31612
rect 9548 31166 9550 31218
rect 9602 31166 9604 31218
rect 9548 31154 9604 31166
rect 10220 31668 10276 34076
rect 10556 34066 10612 34076
rect 10780 33570 10836 34412
rect 10892 33796 10948 37212
rect 11788 37268 11844 37278
rect 11788 37174 11844 37212
rect 11900 37156 11956 37884
rect 12460 38612 12628 38668
rect 12684 38834 13076 38836
rect 12684 38782 13022 38834
rect 13074 38782 13076 38834
rect 12684 38780 13076 38782
rect 12684 38722 12740 38780
rect 13020 38770 13076 38780
rect 12684 38670 12686 38722
rect 12738 38670 12740 38722
rect 12684 38658 12740 38670
rect 12348 37828 12404 37838
rect 12348 37734 12404 37772
rect 12460 37268 12516 38612
rect 13132 38276 13188 39006
rect 13804 38946 13860 38958
rect 13804 38894 13806 38946
rect 13858 38894 13860 38946
rect 13468 38836 13524 38846
rect 13132 38210 13188 38220
rect 13244 38834 13524 38836
rect 13244 38782 13470 38834
rect 13522 38782 13524 38834
rect 13244 38780 13524 38782
rect 12572 37938 12628 37950
rect 12572 37886 12574 37938
rect 12626 37886 12628 37938
rect 12572 37492 12628 37886
rect 12796 37940 12852 37950
rect 12796 37846 12852 37884
rect 12684 37826 12740 37838
rect 12684 37774 12686 37826
rect 12738 37774 12740 37826
rect 12684 37716 12740 37774
rect 12684 37650 12740 37660
rect 12908 37492 12964 37502
rect 13244 37492 13300 38780
rect 13468 38770 13524 38780
rect 12572 37436 12740 37492
rect 12572 37268 12628 37278
rect 12460 37266 12628 37268
rect 12460 37214 12574 37266
rect 12626 37214 12628 37266
rect 12460 37212 12628 37214
rect 12572 37202 12628 37212
rect 12684 37268 12740 37436
rect 12908 37490 13300 37492
rect 12908 37438 12910 37490
rect 12962 37438 13300 37490
rect 12908 37436 13300 37438
rect 13692 37940 13748 37950
rect 12908 37426 12964 37436
rect 12012 37156 12068 37166
rect 12348 37156 12404 37166
rect 11900 37154 12292 37156
rect 11900 37102 12014 37154
rect 12066 37102 12292 37154
rect 11900 37100 12292 37102
rect 12012 37090 12068 37100
rect 11452 37044 11508 37054
rect 11452 36950 11508 36988
rect 11788 34802 11844 34814
rect 11788 34750 11790 34802
rect 11842 34750 11844 34802
rect 11116 34356 11172 34366
rect 11116 34262 11172 34300
rect 11788 34356 11844 34750
rect 11788 34290 11844 34300
rect 11900 34580 11956 34590
rect 11900 34354 11956 34524
rect 11900 34302 11902 34354
rect 11954 34302 11956 34354
rect 11900 34290 11956 34302
rect 12012 34468 12068 34478
rect 12012 34354 12068 34412
rect 12012 34302 12014 34354
rect 12066 34302 12068 34354
rect 11452 34244 11508 34254
rect 11676 34244 11732 34254
rect 11452 34150 11508 34188
rect 11564 34188 11676 34244
rect 11004 34020 11060 34030
rect 11004 33926 11060 33964
rect 10892 33740 11172 33796
rect 10780 33518 10782 33570
rect 10834 33518 10836 33570
rect 10780 33506 10836 33518
rect 10332 33346 10388 33358
rect 10332 33294 10334 33346
rect 10386 33294 10388 33346
rect 10332 32452 10388 33294
rect 10892 33122 10948 33134
rect 10892 33070 10894 33122
rect 10946 33070 10948 33122
rect 10892 32562 10948 33070
rect 11116 33122 11172 33740
rect 11116 33070 11118 33122
rect 11170 33070 11172 33122
rect 11116 33058 11172 33070
rect 11340 32788 11396 32798
rect 11564 32788 11620 34188
rect 11676 34150 11732 34188
rect 11900 34132 11956 34142
rect 11788 34020 11844 34030
rect 11788 33926 11844 33964
rect 11340 32786 11620 32788
rect 11340 32734 11342 32786
rect 11394 32734 11620 32786
rect 11340 32732 11620 32734
rect 11788 33572 11844 33582
rect 11788 33458 11844 33516
rect 11788 33406 11790 33458
rect 11842 33406 11844 33458
rect 11340 32722 11396 32732
rect 10892 32510 10894 32562
rect 10946 32510 10948 32562
rect 10892 32498 10948 32510
rect 11116 32564 11172 32574
rect 11116 32470 11172 32508
rect 11564 32562 11620 32574
rect 11564 32510 11566 32562
rect 11618 32510 11620 32562
rect 10332 32386 10388 32396
rect 10556 32450 10612 32462
rect 10556 32398 10558 32450
rect 10610 32398 10612 32450
rect 10444 32340 10500 32350
rect 10556 32340 10612 32398
rect 11004 32450 11060 32462
rect 11004 32398 11006 32450
rect 11058 32398 11060 32450
rect 11004 32340 11060 32398
rect 11564 32452 11620 32510
rect 11788 32564 11844 33406
rect 11788 32498 11844 32508
rect 11900 33348 11956 34076
rect 12012 33908 12068 34302
rect 12012 33842 12068 33852
rect 11620 32396 11732 32452
rect 11564 32386 11620 32396
rect 10556 32284 11060 32340
rect 10444 32246 10500 32284
rect 11676 31890 11732 32396
rect 11900 32450 11956 33292
rect 11900 32398 11902 32450
rect 11954 32398 11956 32450
rect 11900 32386 11956 32398
rect 12236 33122 12292 37100
rect 12348 37062 12404 37100
rect 12684 37044 12740 37212
rect 13468 37268 13524 37278
rect 13692 37268 13748 37884
rect 13468 37266 13748 37268
rect 13468 37214 13470 37266
rect 13522 37214 13748 37266
rect 13468 37212 13748 37214
rect 12460 36988 12740 37044
rect 13132 37044 13188 37054
rect 12460 36594 12516 36988
rect 12460 36542 12462 36594
rect 12514 36542 12516 36594
rect 12460 36530 12516 36542
rect 12572 36372 12628 36382
rect 12572 34914 12628 36316
rect 13020 36258 13076 36270
rect 13020 36206 13022 36258
rect 13074 36206 13076 36258
rect 12572 34862 12574 34914
rect 12626 34862 12628 34914
rect 12572 34850 12628 34862
rect 12684 35588 12740 35598
rect 12572 34580 12628 34590
rect 12572 34354 12628 34524
rect 12572 34302 12574 34354
rect 12626 34302 12628 34354
rect 12572 34290 12628 34302
rect 12236 33070 12238 33122
rect 12290 33070 12292 33122
rect 12236 32004 12292 33070
rect 12236 31938 12292 31948
rect 11676 31838 11678 31890
rect 11730 31838 11732 31890
rect 11676 31826 11732 31838
rect 9100 30996 9156 31006
rect 9100 30902 9156 30940
rect 9884 30996 9940 31006
rect 9884 30902 9940 30940
rect 10220 30884 10276 31612
rect 11900 31556 11956 31566
rect 10668 30996 10724 31006
rect 10444 30884 10500 30894
rect 10220 30882 10500 30884
rect 10220 30830 10446 30882
rect 10498 30830 10500 30882
rect 10220 30828 10500 30830
rect 10444 30818 10500 30828
rect 10332 30324 10388 30334
rect 10332 30210 10388 30268
rect 10332 30158 10334 30210
rect 10386 30158 10388 30210
rect 9548 30100 9604 30110
rect 9548 30006 9604 30044
rect 8764 29708 9268 29764
rect 8652 29652 8708 29662
rect 8652 29558 8708 29596
rect 8876 29540 8932 29550
rect 8876 29446 8932 29484
rect 8540 29362 8596 29372
rect 8988 29428 9044 29438
rect 8988 29334 9044 29372
rect 8316 28644 8372 28654
rect 8316 28082 8372 28588
rect 8316 28030 8318 28082
rect 8370 28030 8372 28082
rect 8316 28018 8372 28030
rect 8764 28196 8820 28206
rect 8764 27970 8820 28140
rect 8764 27918 8766 27970
rect 8818 27918 8820 27970
rect 8764 27906 8820 27918
rect 8540 27860 8596 27870
rect 8540 27766 8596 27804
rect 8204 26852 8372 26908
rect 8316 25620 8372 26852
rect 9212 26628 9268 29708
rect 9548 28644 9604 28654
rect 9548 28550 9604 28588
rect 10332 28642 10388 30158
rect 10332 28590 10334 28642
rect 10386 28590 10388 28642
rect 10332 28578 10388 28590
rect 10668 29988 10724 30940
rect 10444 28308 10500 28318
rect 9660 28196 9716 28206
rect 9660 28082 9716 28140
rect 9660 28030 9662 28082
rect 9714 28030 9716 28082
rect 9660 28018 9716 28030
rect 10444 28082 10500 28252
rect 10444 28030 10446 28082
rect 10498 28030 10500 28082
rect 10444 28018 10500 28030
rect 10332 27746 10388 27758
rect 10332 27694 10334 27746
rect 10386 27694 10388 27746
rect 10220 27636 10276 27646
rect 10108 27634 10276 27636
rect 10108 27582 10222 27634
rect 10274 27582 10276 27634
rect 10108 27580 10276 27582
rect 10108 27188 10164 27580
rect 10220 27570 10276 27580
rect 9996 27132 10164 27188
rect 9212 26562 9268 26572
rect 9436 27074 9492 27086
rect 9436 27022 9438 27074
rect 9490 27022 9492 27074
rect 9436 26292 9492 27022
rect 9996 26908 10052 27132
rect 10332 27076 10388 27694
rect 10220 27020 10388 27076
rect 9884 26852 10052 26908
rect 10108 26964 10164 26974
rect 10220 26964 10276 27020
rect 10108 26962 10276 26964
rect 10108 26910 10110 26962
rect 10162 26910 10276 26962
rect 10108 26908 10276 26910
rect 10108 26898 10164 26908
rect 8316 25506 8372 25564
rect 8316 25454 8318 25506
rect 8370 25454 8372 25506
rect 8316 25442 8372 25454
rect 8540 26178 8596 26190
rect 8540 26126 8542 26178
rect 8594 26126 8596 26178
rect 7756 25218 7812 25228
rect 8540 25284 8596 26126
rect 9436 25396 9492 26236
rect 9660 26516 9716 26526
rect 9660 26290 9716 26460
rect 9660 26238 9662 26290
rect 9714 26238 9716 26290
rect 9660 26226 9716 26238
rect 9884 26402 9940 26852
rect 10332 26516 10388 26526
rect 10668 26516 10724 29932
rect 10892 30996 10948 31006
rect 10892 30324 10948 30940
rect 10892 29426 10948 30268
rect 11228 30210 11284 30222
rect 11228 30158 11230 30210
rect 11282 30158 11284 30210
rect 11228 29540 11284 30158
rect 11900 30210 11956 31500
rect 12572 31554 12628 31566
rect 12572 31502 12574 31554
rect 12626 31502 12628 31554
rect 12572 31444 12628 31502
rect 12572 31378 12628 31388
rect 12572 30884 12628 30894
rect 12012 30882 12628 30884
rect 12012 30830 12574 30882
rect 12626 30830 12628 30882
rect 12012 30828 12628 30830
rect 12012 30434 12068 30828
rect 12572 30818 12628 30828
rect 12012 30382 12014 30434
rect 12066 30382 12068 30434
rect 12012 30370 12068 30382
rect 11900 30158 11902 30210
rect 11954 30158 11956 30210
rect 11900 30146 11956 30158
rect 12460 29988 12516 29998
rect 12460 29894 12516 29932
rect 11228 29474 11284 29484
rect 10892 29374 10894 29426
rect 10946 29374 10948 29426
rect 10892 29362 10948 29374
rect 11564 29314 11620 29326
rect 11564 29262 11566 29314
rect 11618 29262 11620 29314
rect 11116 28756 11172 28766
rect 11116 28662 11172 28700
rect 11564 28756 11620 29262
rect 11564 28690 11620 28700
rect 12236 28868 12292 28878
rect 10780 28644 10836 28654
rect 10780 28550 10836 28588
rect 11004 28642 11060 28654
rect 11004 28590 11006 28642
rect 11058 28590 11060 28642
rect 11004 28308 11060 28590
rect 11340 28642 11396 28654
rect 12236 28644 12292 28812
rect 11340 28590 11342 28642
rect 11394 28590 11396 28642
rect 11340 28420 11396 28590
rect 11900 28642 12292 28644
rect 11900 28590 12238 28642
rect 12290 28590 12292 28642
rect 11900 28588 12292 28590
rect 11676 28532 11732 28542
rect 11676 28438 11732 28476
rect 11564 28420 11620 28430
rect 11340 28364 11564 28420
rect 11564 28326 11620 28364
rect 11788 28418 11844 28430
rect 11788 28366 11790 28418
rect 11842 28366 11844 28418
rect 11004 28242 11060 28252
rect 11788 28308 11844 28366
rect 11788 28242 11844 28252
rect 10332 26514 10668 26516
rect 10332 26462 10334 26514
rect 10386 26462 10668 26514
rect 10332 26460 10668 26462
rect 10332 26450 10388 26460
rect 10668 26450 10724 26460
rect 11676 28196 11732 28206
rect 9884 26350 9886 26402
rect 9938 26350 9940 26402
rect 9436 25330 9492 25340
rect 8540 25218 8596 25228
rect 9772 25284 9828 25294
rect 9884 25284 9940 26350
rect 10780 26292 10836 26302
rect 10780 26198 10836 26236
rect 11452 26178 11508 26190
rect 11452 26126 11454 26178
rect 11506 26126 11508 26178
rect 11004 25396 11060 25406
rect 9884 25228 10164 25284
rect 7308 24894 7310 24946
rect 7362 24894 7364 24946
rect 7308 24882 7364 24894
rect 7420 24948 7476 24958
rect 7420 24946 8036 24948
rect 7420 24894 7422 24946
rect 7474 24894 8036 24946
rect 7420 24892 8036 24894
rect 7420 24882 7476 24892
rect 7980 24834 8036 24892
rect 9772 24946 9828 25228
rect 9772 24894 9774 24946
rect 9826 24894 9828 24946
rect 9772 24882 9828 24894
rect 7980 24782 7982 24834
rect 8034 24782 8036 24834
rect 7084 24098 7140 24108
rect 7756 24164 7812 24174
rect 7980 24164 8036 24782
rect 6412 23156 6468 23166
rect 6300 23154 6468 23156
rect 6300 23102 6414 23154
rect 6466 23102 6468 23154
rect 6300 23100 6468 23102
rect 5740 22260 5796 22270
rect 5740 22166 5796 22204
rect 5852 22258 5908 23100
rect 6412 23090 6468 23100
rect 5852 22206 5854 22258
rect 5906 22206 5908 22258
rect 5852 21924 5908 22206
rect 5292 21586 5684 21588
rect 5292 21534 5294 21586
rect 5346 21534 5684 21586
rect 5292 21532 5684 21534
rect 5740 21868 5908 21924
rect 5964 22932 6020 22942
rect 4620 21476 4676 21486
rect 4060 21474 4676 21476
rect 4060 21422 4622 21474
rect 4674 21422 4676 21474
rect 4060 21420 4676 21422
rect 3612 20526 3614 20578
rect 3666 20526 3668 20578
rect 3612 20514 3668 20526
rect 3948 20580 4004 20590
rect 4060 20580 4116 21420
rect 4620 21410 4676 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4620 20802 4676 20814
rect 4620 20750 4622 20802
rect 4674 20750 4676 20802
rect 4004 20524 4116 20580
rect 4172 20690 4228 20702
rect 4172 20638 4174 20690
rect 4226 20638 4228 20690
rect 3948 20514 4004 20524
rect 3388 20076 3556 20132
rect 3388 19906 3444 19918
rect 3388 19854 3390 19906
rect 3442 19854 3444 19906
rect 3052 19796 3108 19806
rect 2716 17614 2718 17666
rect 2770 17614 2772 17666
rect 2716 17602 2772 17614
rect 2828 19348 2884 19358
rect 2828 17554 2884 19292
rect 3052 17666 3108 19740
rect 3388 18564 3444 19854
rect 3500 19348 3556 20076
rect 3500 19282 3556 19292
rect 3388 18498 3444 18508
rect 3836 19012 3892 19022
rect 3052 17614 3054 17666
rect 3106 17614 3108 17666
rect 3052 17602 3108 17614
rect 3836 17666 3892 18956
rect 3836 17614 3838 17666
rect 3890 17614 3892 17666
rect 3836 17602 3892 17614
rect 4172 17666 4228 20638
rect 4508 20690 4564 20702
rect 4508 20638 4510 20690
rect 4562 20638 4564 20690
rect 4284 20578 4340 20590
rect 4284 20526 4286 20578
rect 4338 20526 4340 20578
rect 4284 19124 4340 20526
rect 4508 19796 4564 20638
rect 4620 20356 4676 20750
rect 4620 19908 4676 20300
rect 4620 19842 4676 19852
rect 4508 19730 4564 19740
rect 5292 19796 5348 21532
rect 5740 21476 5796 21868
rect 5964 21812 6020 22876
rect 6300 22146 6356 22158
rect 6300 22094 6302 22146
rect 6354 22094 6356 22146
rect 6300 21812 6356 22094
rect 5964 21810 6132 21812
rect 5964 21758 5966 21810
rect 6018 21758 6132 21810
rect 5964 21756 6132 21758
rect 5964 21746 6020 21756
rect 5852 21700 5908 21710
rect 5852 21606 5908 21644
rect 5740 21420 5908 21476
rect 5292 19730 5348 19740
rect 5516 20020 5572 20030
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4732 19460 4788 19470
rect 4620 19348 4676 19358
rect 4620 19254 4676 19292
rect 4284 19058 4340 19068
rect 4620 18340 4676 18350
rect 4732 18340 4788 19404
rect 5516 19234 5572 19964
rect 5516 19182 5518 19234
rect 5570 19182 5572 19234
rect 5516 19170 5572 19182
rect 5740 19348 5796 19358
rect 5740 19122 5796 19292
rect 5740 19070 5742 19122
rect 5794 19070 5796 19122
rect 5740 19058 5796 19070
rect 5852 19122 5908 21420
rect 5852 19070 5854 19122
rect 5906 19070 5908 19122
rect 5852 19012 5908 19070
rect 5852 18946 5908 18956
rect 5964 20802 6020 20814
rect 5964 20750 5966 20802
rect 6018 20750 6020 20802
rect 5740 18900 5796 18910
rect 5292 18564 5348 18574
rect 5292 18450 5348 18508
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5292 18386 5348 18398
rect 4172 17614 4174 17666
rect 4226 17614 4228 17666
rect 4172 17602 4228 17614
rect 4284 18338 4788 18340
rect 4284 18286 4622 18338
rect 4674 18286 4788 18338
rect 4284 18284 4788 18286
rect 2828 17502 2830 17554
rect 2882 17502 2884 17554
rect 2828 17490 2884 17502
rect 3948 17444 4004 17454
rect 4284 17444 4340 18284
rect 4620 18274 4676 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5740 17554 5796 18844
rect 5852 18564 5908 18574
rect 5964 18564 6020 20750
rect 6076 19460 6132 21756
rect 6188 21586 6244 21598
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 6188 20244 6244 21534
rect 6300 20580 6356 21756
rect 6300 20514 6356 20524
rect 6188 20188 6468 20244
rect 6300 20020 6356 20030
rect 6076 19394 6132 19404
rect 6188 19908 6244 19918
rect 6188 19234 6244 19852
rect 6188 19182 6190 19234
rect 6242 19182 6244 19234
rect 6188 18900 6244 19182
rect 6188 18834 6244 18844
rect 5908 18508 6020 18564
rect 5852 18498 5908 18508
rect 6076 18450 6132 18462
rect 6076 18398 6078 18450
rect 6130 18398 6132 18450
rect 6076 17892 6132 18398
rect 5740 17502 5742 17554
rect 5794 17502 5796 17554
rect 5740 17490 5796 17502
rect 5964 17836 6132 17892
rect 3948 17442 4340 17444
rect 3948 17390 3950 17442
rect 4002 17390 4340 17442
rect 3948 17388 4340 17390
rect 3948 17378 4004 17388
rect 5964 17108 6020 17836
rect 6300 17780 6356 19964
rect 6412 19234 6468 20188
rect 6412 19182 6414 19234
rect 6466 19182 6468 19234
rect 6412 19170 6468 19182
rect 6524 19124 6580 23660
rect 6636 24052 6692 24062
rect 6636 23154 6692 23996
rect 7196 24052 7252 24062
rect 7644 24052 7700 24062
rect 7196 24050 7700 24052
rect 7196 23998 7198 24050
rect 7250 23998 7646 24050
rect 7698 23998 7700 24050
rect 7196 23996 7700 23998
rect 7196 23986 7252 23996
rect 7644 23986 7700 23996
rect 7756 24050 7812 24108
rect 7756 23998 7758 24050
rect 7810 23998 7812 24050
rect 7756 23986 7812 23998
rect 7868 24108 8036 24164
rect 8092 24834 8148 24846
rect 8092 24782 8094 24834
rect 8146 24782 8148 24834
rect 6860 23938 6916 23950
rect 6860 23886 6862 23938
rect 6914 23886 6916 23938
rect 6860 23380 6916 23886
rect 7084 23938 7140 23950
rect 7084 23886 7086 23938
rect 7138 23886 7140 23938
rect 7084 23716 7140 23886
rect 7308 23828 7364 23838
rect 7308 23734 7364 23772
rect 7084 23650 7140 23660
rect 6860 23324 7700 23380
rect 7644 23266 7700 23324
rect 7644 23214 7646 23266
rect 7698 23214 7700 23266
rect 7644 23202 7700 23214
rect 6860 23156 6916 23166
rect 6636 23102 6638 23154
rect 6690 23102 6692 23154
rect 6636 23090 6692 23102
rect 6748 23100 6860 23156
rect 6748 22482 6804 23100
rect 6860 23062 6916 23100
rect 7196 23156 7252 23166
rect 7532 23156 7588 23166
rect 7196 23154 7588 23156
rect 7196 23102 7198 23154
rect 7250 23102 7534 23154
rect 7586 23102 7588 23154
rect 7196 23100 7588 23102
rect 7196 23090 7252 23100
rect 7532 23090 7588 23100
rect 7756 23154 7812 23166
rect 7756 23102 7758 23154
rect 7810 23102 7812 23154
rect 7084 22932 7140 22942
rect 7084 22838 7140 22876
rect 6748 22430 6750 22482
rect 6802 22430 6804 22482
rect 6748 22418 6804 22430
rect 7756 22484 7812 23102
rect 7756 22418 7812 22428
rect 7868 22260 7924 24108
rect 8092 24052 8148 24782
rect 8540 24836 8596 24846
rect 8316 24724 8372 24734
rect 8316 24630 8372 24668
rect 8092 23986 8148 23996
rect 7980 23940 8036 23978
rect 7980 23874 8036 23884
rect 8204 23828 8260 23838
rect 7980 23716 8036 23726
rect 8036 23660 8148 23716
rect 7980 23650 8036 23660
rect 8092 22932 8148 23660
rect 8204 23156 8260 23772
rect 8540 23492 8596 24780
rect 8652 24834 8708 24846
rect 8652 24782 8654 24834
rect 8706 24782 8708 24834
rect 8652 24052 8708 24782
rect 8652 23958 8708 23996
rect 8876 24722 8932 24734
rect 9436 24724 9492 24734
rect 8876 24670 8878 24722
rect 8930 24670 8932 24722
rect 8204 23062 8260 23100
rect 8316 23436 8596 23492
rect 7756 22204 7924 22260
rect 7980 22930 8148 22932
rect 7980 22878 8094 22930
rect 8146 22878 8148 22930
rect 7980 22876 8148 22878
rect 7084 21924 7140 21934
rect 6972 21812 7028 21822
rect 6972 21718 7028 21756
rect 7084 21698 7140 21868
rect 7084 21646 7086 21698
rect 7138 21646 7140 21698
rect 7084 21634 7140 21646
rect 7756 21698 7812 22204
rect 7868 21812 7924 21822
rect 7980 21812 8036 22876
rect 8092 22866 8148 22876
rect 7924 21756 8036 21812
rect 8316 21924 8372 23436
rect 7868 21718 7924 21756
rect 7756 21646 7758 21698
rect 7810 21646 7812 21698
rect 6748 21586 6804 21598
rect 6748 21534 6750 21586
rect 6802 21534 6804 21586
rect 6636 20690 6692 20702
rect 6636 20638 6638 20690
rect 6690 20638 6692 20690
rect 6636 19346 6692 20638
rect 6636 19294 6638 19346
rect 6690 19294 6692 19346
rect 6636 19282 6692 19294
rect 6748 19234 6804 21534
rect 7756 20692 7812 21646
rect 8316 21698 8372 21868
rect 8428 23268 8484 23278
rect 8540 23268 8596 23436
rect 8652 23268 8708 23278
rect 8540 23266 8708 23268
rect 8540 23214 8654 23266
rect 8706 23214 8708 23266
rect 8540 23212 8708 23214
rect 8428 21810 8484 23212
rect 8652 23202 8708 23212
rect 8764 23266 8820 23278
rect 8764 23214 8766 23266
rect 8818 23214 8820 23266
rect 8764 23156 8820 23214
rect 8876 23156 8932 24670
rect 8988 24722 9492 24724
rect 8988 24670 9438 24722
rect 9490 24670 9492 24722
rect 8988 24668 9492 24670
rect 8988 23378 9044 24668
rect 9436 24658 9492 24668
rect 9772 24724 9828 24734
rect 9772 24630 9828 24668
rect 10108 24722 10164 25228
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 8988 23326 8990 23378
rect 9042 23326 9044 23378
rect 8988 23314 9044 23326
rect 9772 23828 9828 23838
rect 9772 23378 9828 23772
rect 9772 23326 9774 23378
rect 9826 23326 9828 23378
rect 9772 23314 9828 23326
rect 9436 23156 9492 23166
rect 8876 23154 9492 23156
rect 8876 23102 9438 23154
rect 9490 23102 9492 23154
rect 8876 23100 9492 23102
rect 8764 22708 8820 23100
rect 9436 23090 9492 23100
rect 9884 23156 9940 23166
rect 9884 23062 9940 23100
rect 10108 23154 10164 24670
rect 11004 24722 11060 25340
rect 11004 24670 11006 24722
rect 11058 24670 11060 24722
rect 11004 24658 11060 24670
rect 11452 24164 11508 26126
rect 11452 24098 11508 24108
rect 11452 23938 11508 23950
rect 11452 23886 11454 23938
rect 11506 23886 11508 23938
rect 10780 23828 10836 23838
rect 10780 23734 10836 23772
rect 10556 23268 10612 23278
rect 10556 23174 10612 23212
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 8764 22642 8820 22652
rect 9660 22372 9716 22382
rect 9996 22372 10052 22382
rect 9660 22370 9996 22372
rect 9660 22318 9662 22370
rect 9714 22318 9996 22370
rect 9660 22316 9996 22318
rect 9660 22306 9716 22316
rect 8876 22260 8932 22270
rect 8876 22258 9604 22260
rect 8876 22206 8878 22258
rect 8930 22206 9604 22258
rect 8876 22204 9604 22206
rect 8876 22194 8932 22204
rect 8428 21758 8430 21810
rect 8482 21758 8484 21810
rect 8428 21746 8484 21758
rect 8540 21812 8596 21822
rect 9548 21812 9604 22204
rect 9660 21812 9716 21822
rect 9548 21810 9716 21812
rect 9548 21758 9662 21810
rect 9714 21758 9716 21810
rect 9548 21756 9716 21758
rect 8316 21646 8318 21698
rect 8370 21646 8372 21698
rect 8316 21634 8372 21646
rect 8092 21588 8148 21598
rect 8092 21494 8148 21532
rect 7756 20626 7812 20636
rect 8428 21476 8484 21486
rect 8092 20132 8148 20142
rect 8092 19458 8148 20076
rect 8204 20018 8260 20030
rect 8204 19966 8206 20018
rect 8258 19966 8260 20018
rect 8204 19908 8260 19966
rect 8204 19842 8260 19852
rect 8092 19406 8094 19458
rect 8146 19406 8148 19458
rect 8092 19394 8148 19406
rect 8428 19460 8484 21420
rect 8540 20916 8596 21756
rect 9660 21746 9716 21756
rect 8652 21588 8708 21598
rect 9436 21588 9492 21598
rect 8652 21586 9492 21588
rect 8652 21534 8654 21586
rect 8706 21534 9438 21586
rect 9490 21534 9492 21586
rect 8652 21532 9492 21534
rect 8652 21522 8708 21532
rect 9436 21522 9492 21532
rect 9772 21588 9828 21598
rect 9772 21494 9828 21532
rect 9996 21476 10052 22316
rect 10108 21698 10164 23102
rect 10332 23156 10388 23166
rect 10332 23062 10388 23100
rect 10668 23154 10724 23166
rect 10668 23102 10670 23154
rect 10722 23102 10724 23154
rect 10108 21646 10110 21698
rect 10162 21646 10164 21698
rect 10108 21634 10164 21646
rect 9996 21420 10164 21476
rect 8764 20916 8820 20926
rect 8540 20914 8820 20916
rect 8540 20862 8766 20914
rect 8818 20862 8820 20914
rect 8540 20860 8820 20862
rect 8764 20850 8820 20860
rect 9436 20692 9492 20702
rect 9436 20598 9492 20636
rect 9100 20580 9156 20590
rect 8876 20578 9156 20580
rect 8876 20526 9102 20578
rect 9154 20526 9156 20578
rect 8876 20524 9156 20526
rect 8540 20130 8596 20142
rect 8540 20078 8542 20130
rect 8594 20078 8596 20130
rect 8540 19796 8596 20078
rect 8876 20132 8932 20524
rect 9100 20514 9156 20524
rect 8876 20038 8932 20076
rect 10108 20132 10164 21420
rect 10668 20692 10724 23102
rect 11452 22372 11508 23886
rect 11452 22306 11508 22316
rect 10780 22258 10836 22270
rect 10780 22206 10782 22258
rect 10834 22206 10836 22258
rect 10780 21812 10836 22206
rect 10780 21746 10836 21756
rect 10668 20626 10724 20636
rect 10892 20914 10948 20926
rect 10892 20862 10894 20914
rect 10946 20862 10948 20914
rect 9772 19908 9828 19918
rect 9772 19814 9828 19852
rect 8540 19730 8596 19740
rect 8540 19460 8596 19470
rect 8428 19458 8596 19460
rect 8428 19406 8542 19458
rect 8594 19406 8596 19458
rect 8428 19404 8596 19406
rect 8540 19394 8596 19404
rect 6748 19182 6750 19234
rect 6802 19182 6804 19234
rect 6748 19170 6804 19182
rect 7532 19234 7588 19246
rect 7532 19182 7534 19234
rect 7586 19182 7588 19234
rect 6524 19068 6692 19124
rect 6524 17780 6580 17790
rect 6076 17778 6580 17780
rect 6076 17726 6526 17778
rect 6578 17726 6580 17778
rect 6076 17724 6580 17726
rect 6076 17666 6132 17724
rect 6524 17714 6580 17724
rect 6076 17614 6078 17666
rect 6130 17614 6132 17666
rect 6076 17602 6132 17614
rect 5964 17052 6356 17108
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 15314 1876 16830
rect 6188 16882 6244 16894
rect 6188 16830 6190 16882
rect 6242 16830 6244 16882
rect 2492 16770 2548 16782
rect 2492 16718 2494 16770
rect 2546 16718 2548 16770
rect 2492 16324 2548 16718
rect 4620 16772 4676 16782
rect 4620 16678 4676 16716
rect 5516 16772 5572 16782
rect 4956 16660 5012 16670
rect 4844 16658 5012 16660
rect 4844 16606 4958 16658
rect 5010 16606 5012 16658
rect 4844 16604 5012 16606
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2492 16258 2548 16268
rect 4732 16324 4788 16334
rect 4732 16230 4788 16268
rect 4060 16098 4116 16110
rect 4060 16046 4062 16098
rect 4114 16046 4116 16098
rect 3500 15874 3556 15886
rect 3500 15822 3502 15874
rect 3554 15822 3556 15874
rect 3500 15652 3556 15822
rect 3500 15586 3556 15596
rect 3724 15874 3780 15886
rect 3724 15822 3726 15874
rect 3778 15822 3780 15874
rect 1820 15262 1822 15314
rect 1874 15262 1876 15314
rect 1820 15250 1876 15262
rect 2492 15204 2548 15214
rect 2492 15202 3220 15204
rect 2492 15150 2494 15202
rect 2546 15150 3220 15202
rect 2492 15148 3220 15150
rect 3724 15148 3780 15822
rect 2492 15138 2548 15148
rect 3164 14754 3220 15148
rect 3612 15092 3780 15148
rect 3836 15652 3892 15662
rect 4060 15652 4116 16046
rect 3892 15596 4116 15652
rect 4284 16098 4340 16110
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 3612 14756 3668 15092
rect 3164 14702 3166 14754
rect 3218 14702 3220 14754
rect 3164 14690 3220 14702
rect 3276 14700 3668 14756
rect 3276 14418 3332 14700
rect 3276 14366 3278 14418
rect 3330 14366 3332 14418
rect 3276 14354 3332 14366
rect 3388 14084 3444 14700
rect 3500 14420 3556 14430
rect 3500 14418 3780 14420
rect 3500 14366 3502 14418
rect 3554 14366 3780 14418
rect 3500 14364 3780 14366
rect 3500 14354 3556 14364
rect 3724 14084 3780 14364
rect 3836 14306 3892 15596
rect 4284 15092 4340 16046
rect 4844 15986 4900 16604
rect 4956 16594 5012 16604
rect 5292 16658 5348 16670
rect 5292 16606 5294 16658
rect 5346 16606 5348 16658
rect 4844 15934 4846 15986
rect 4898 15934 4900 15986
rect 4732 15652 4788 15662
rect 4844 15652 4900 15934
rect 5068 15986 5124 15998
rect 5068 15934 5070 15986
rect 5122 15934 5124 15986
rect 5068 15764 5124 15934
rect 5292 15876 5348 16606
rect 5516 16436 5572 16716
rect 5516 16380 5908 16436
rect 5852 16098 5908 16380
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5852 16034 5908 16046
rect 5628 15876 5684 15886
rect 5292 15874 5684 15876
rect 5292 15822 5630 15874
rect 5682 15822 5684 15874
rect 5292 15820 5684 15822
rect 5628 15764 5684 15820
rect 5068 15708 5572 15764
rect 4844 15596 5012 15652
rect 4620 15202 4676 15214
rect 4620 15150 4622 15202
rect 4674 15150 4676 15202
rect 4620 15092 4676 15150
rect 4732 15148 4788 15596
rect 4732 15092 4900 15148
rect 4284 15036 4676 15092
rect 4060 14532 4116 14542
rect 4284 14532 4340 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14642 4900 15092
rect 4844 14590 4846 14642
rect 4898 14590 4900 14642
rect 4844 14578 4900 14590
rect 4060 14530 4340 14532
rect 4060 14478 4062 14530
rect 4114 14478 4340 14530
rect 4060 14476 4340 14478
rect 4396 14532 4452 14542
rect 4060 14466 4116 14476
rect 4396 14438 4452 14476
rect 3836 14254 3838 14306
rect 3890 14254 3892 14306
rect 3836 14242 3892 14254
rect 3948 14306 4004 14318
rect 3948 14254 3950 14306
rect 4002 14254 4004 14306
rect 3948 14084 4004 14254
rect 3388 14028 3668 14084
rect 3724 14028 4004 14084
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 12178 1876 13694
rect 3612 13748 3668 14028
rect 4956 13860 5012 15596
rect 5516 15540 5572 15708
rect 5628 15698 5684 15708
rect 5740 15874 5796 15886
rect 6076 15876 6132 15886
rect 5740 15822 5742 15874
rect 5794 15822 5796 15874
rect 5740 15540 5796 15822
rect 5964 15874 6132 15876
rect 5964 15822 6078 15874
rect 6130 15822 6132 15874
rect 5964 15820 6132 15822
rect 5964 15540 6020 15820
rect 6076 15810 6132 15820
rect 5516 15484 5796 15540
rect 5852 15484 6020 15540
rect 5852 14532 5908 15484
rect 6076 15316 6132 15326
rect 6188 15316 6244 16830
rect 6132 15260 6244 15316
rect 6076 15222 6132 15260
rect 6300 15148 6356 17052
rect 5628 14420 5684 14430
rect 5628 14326 5684 14364
rect 5852 13972 5908 14476
rect 5964 15092 6356 15148
rect 5964 14418 6020 15092
rect 5964 14366 5966 14418
rect 6018 14366 6020 14418
rect 5964 14354 6020 14366
rect 6636 14418 6692 19068
rect 7196 19012 7252 19022
rect 7532 19012 7588 19182
rect 7756 19236 7812 19246
rect 7756 19142 7812 19180
rect 8652 19236 8708 19246
rect 7196 19010 7532 19012
rect 7196 18958 7198 19010
rect 7250 18958 7532 19010
rect 7196 18956 7532 18958
rect 7196 18946 7252 18956
rect 7532 18946 7588 18956
rect 8540 19012 8596 19022
rect 8540 18564 8596 18956
rect 8652 18674 8708 19180
rect 10108 19234 10164 20076
rect 10332 20580 10388 20590
rect 10332 20020 10388 20524
rect 10108 19182 10110 19234
rect 10162 19182 10164 19234
rect 9100 19012 9156 19022
rect 9100 18918 9156 18956
rect 8652 18622 8654 18674
rect 8706 18622 8708 18674
rect 8652 18610 8708 18622
rect 8092 18508 8596 18564
rect 6860 16772 6916 16782
rect 6860 16678 6916 16716
rect 6636 14366 6638 14418
rect 6690 14366 6692 14418
rect 6300 14308 6356 14318
rect 6188 14306 6356 14308
rect 6188 14254 6302 14306
rect 6354 14254 6356 14306
rect 6188 14252 6356 14254
rect 6188 14084 6244 14252
rect 6300 14242 6356 14252
rect 5852 13970 6132 13972
rect 5852 13918 5854 13970
rect 5906 13918 6132 13970
rect 5852 13916 6132 13918
rect 5852 13906 5908 13916
rect 4956 13804 5124 13860
rect 1820 12126 1822 12178
rect 1874 12126 1876 12178
rect 1820 10612 1876 12126
rect 2268 13636 2324 13646
rect 2044 10612 2100 10622
rect 1820 10610 2100 10612
rect 1820 10558 2046 10610
rect 2098 10558 2100 10610
rect 1820 10556 2100 10558
rect 1820 9828 1876 9838
rect 2044 9828 2100 10556
rect 1820 9826 2100 9828
rect 1820 9774 1822 9826
rect 1874 9774 2100 9826
rect 1820 9772 2100 9774
rect 1820 8484 1876 9772
rect 1708 7362 1764 7374
rect 1708 7310 1710 7362
rect 1762 7310 1764 7362
rect 1708 6692 1764 7310
rect 1708 6626 1764 6636
rect 1820 5906 1876 8428
rect 2268 9266 2324 13580
rect 2492 13636 2548 13646
rect 2492 13634 2996 13636
rect 2492 13582 2494 13634
rect 2546 13582 2996 13634
rect 2492 13580 2996 13582
rect 2492 13570 2548 13580
rect 2940 13186 2996 13580
rect 2940 13134 2942 13186
rect 2994 13134 2996 13186
rect 2940 13122 2996 13134
rect 3052 13076 3108 13086
rect 3052 12852 3108 13020
rect 3276 12852 3332 12862
rect 3052 12850 3220 12852
rect 3052 12798 3054 12850
rect 3106 12798 3220 12850
rect 3052 12796 3220 12798
rect 3052 12786 3108 12796
rect 2492 12066 2548 12078
rect 2492 12014 2494 12066
rect 2546 12014 2548 12066
rect 2492 10836 2548 12014
rect 3164 11844 3220 12796
rect 3276 12758 3332 12796
rect 3612 12738 3668 13692
rect 4620 13636 4676 13646
rect 4956 13636 5012 13646
rect 4620 13634 5012 13636
rect 4620 13582 4622 13634
rect 4674 13582 4958 13634
rect 5010 13582 5012 13634
rect 4620 13580 5012 13582
rect 4620 13524 4676 13580
rect 4956 13570 5012 13580
rect 4284 13468 4676 13524
rect 3836 12964 3892 12974
rect 4284 12964 4340 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 5068 13300 5124 13804
rect 5180 13748 5236 13758
rect 5180 13654 5236 13692
rect 5516 13524 5572 13534
rect 5516 13522 5796 13524
rect 5516 13470 5518 13522
rect 5570 13470 5796 13522
rect 5516 13468 5796 13470
rect 5516 13458 5572 13468
rect 4476 13290 4740 13300
rect 4844 13244 5684 13300
rect 4732 13188 4788 13198
rect 4844 13188 4900 13244
rect 4732 13186 4900 13188
rect 4732 13134 4734 13186
rect 4786 13134 4900 13186
rect 4732 13132 4900 13134
rect 4732 13122 4788 13132
rect 3836 12962 4340 12964
rect 3836 12910 3838 12962
rect 3890 12910 4340 12962
rect 3836 12908 4340 12910
rect 4508 12964 4564 12974
rect 4564 12908 4676 12964
rect 3836 12898 3892 12908
rect 4508 12870 4564 12908
rect 3724 12852 3780 12862
rect 3724 12758 3780 12796
rect 3612 12686 3614 12738
rect 3666 12686 3668 12738
rect 3612 12674 3668 12686
rect 4060 12738 4116 12750
rect 4060 12686 4062 12738
rect 4114 12686 4116 12738
rect 4060 12628 4116 12686
rect 4172 12628 4228 12638
rect 4060 12572 4172 12628
rect 4172 12562 4228 12572
rect 4620 12066 4676 12908
rect 5628 12962 5684 13244
rect 5740 13076 5796 13468
rect 5740 13010 5796 13020
rect 5628 12910 5630 12962
rect 5682 12910 5684 12962
rect 5628 12898 5684 12910
rect 5852 12964 5908 12974
rect 5852 12870 5908 12908
rect 6076 12850 6132 13916
rect 6188 13970 6244 14028
rect 6188 13918 6190 13970
rect 6242 13918 6244 13970
rect 6188 13906 6244 13918
rect 6636 13636 6692 14366
rect 6748 15202 6804 15214
rect 6748 15150 6750 15202
rect 6802 15150 6804 15202
rect 6748 13972 6804 15150
rect 7084 15092 7140 15102
rect 7084 14530 7140 15036
rect 8092 14756 8148 18508
rect 8204 18340 8260 18350
rect 8540 18340 8596 18350
rect 8204 18338 8596 18340
rect 8204 18286 8206 18338
rect 8258 18286 8542 18338
rect 8594 18286 8596 18338
rect 8204 18284 8596 18286
rect 8204 18274 8260 18284
rect 8540 18274 8596 18284
rect 10108 17668 10164 19182
rect 9660 17666 10164 17668
rect 9660 17614 10110 17666
rect 10162 17614 10164 17666
rect 9660 17612 10164 17614
rect 9660 16884 9716 17612
rect 10108 17602 10164 17612
rect 10220 19964 10388 20020
rect 9660 16790 9716 16828
rect 10108 17108 10164 17118
rect 8988 16770 9044 16782
rect 8988 16718 8990 16770
rect 9042 16718 9044 16770
rect 8988 16324 9044 16718
rect 8652 16268 9828 16324
rect 8652 16210 8708 16268
rect 8652 16158 8654 16210
rect 8706 16158 8708 16210
rect 8652 16146 8708 16158
rect 8876 16100 8932 16110
rect 8876 16006 8932 16044
rect 9548 16100 9604 16110
rect 9548 16006 9604 16044
rect 9772 16098 9828 16268
rect 9772 16046 9774 16098
rect 9826 16046 9828 16098
rect 9772 16034 9828 16046
rect 10108 16098 10164 17052
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 10108 16034 10164 16046
rect 9660 15988 9716 15998
rect 9660 15894 9716 15932
rect 9212 15876 9268 15886
rect 9212 15782 9268 15820
rect 10108 15876 10164 15886
rect 10108 15538 10164 15820
rect 10220 15764 10276 19964
rect 10780 19122 10836 19134
rect 10780 19070 10782 19122
rect 10834 19070 10836 19122
rect 10780 18452 10836 19070
rect 10780 18386 10836 18396
rect 10892 18340 10948 20862
rect 11228 20690 11284 20702
rect 11228 20638 11230 20690
rect 11282 20638 11284 20690
rect 11004 20580 11060 20590
rect 11004 20486 11060 20524
rect 11228 19460 11284 20638
rect 11228 19394 11284 19404
rect 11004 18732 11396 18788
rect 11004 18674 11060 18732
rect 11004 18622 11006 18674
rect 11058 18622 11060 18674
rect 11004 18610 11060 18622
rect 10892 18284 11060 18340
rect 10780 17780 10836 17790
rect 11004 17780 11060 18284
rect 10780 17778 11060 17780
rect 10780 17726 10782 17778
rect 10834 17726 11060 17778
rect 10780 17724 11060 17726
rect 11116 18338 11172 18350
rect 11116 18286 11118 18338
rect 11170 18286 11172 18338
rect 10780 17714 10836 17724
rect 11116 17444 11172 18286
rect 10332 17388 11172 17444
rect 11228 18226 11284 18238
rect 11228 18174 11230 18226
rect 11282 18174 11284 18226
rect 10332 16994 10388 17388
rect 10332 16942 10334 16994
rect 10386 16942 10388 16994
rect 10332 16930 10388 16942
rect 10780 17108 10836 17118
rect 10556 16772 10612 16782
rect 10556 16210 10612 16716
rect 10556 16158 10558 16210
rect 10610 16158 10612 16210
rect 10556 16146 10612 16158
rect 10444 15988 10500 15998
rect 10444 15894 10500 15932
rect 10668 15876 10724 15886
rect 10668 15782 10724 15820
rect 10220 15708 10500 15764
rect 10108 15486 10110 15538
rect 10162 15486 10164 15538
rect 8876 15316 8932 15326
rect 8876 15202 8932 15260
rect 8876 15150 8878 15202
rect 8930 15150 8932 15202
rect 8876 15138 8932 15150
rect 8988 15204 9044 15214
rect 10108 15148 10164 15486
rect 10332 15316 10388 15326
rect 7756 14644 7812 14654
rect 7756 14550 7812 14588
rect 7084 14478 7086 14530
rect 7138 14478 7140 14530
rect 6748 13906 6804 13916
rect 6972 14420 7028 14430
rect 6972 13970 7028 14364
rect 7084 14308 7140 14478
rect 7084 14242 7140 14252
rect 7980 13972 8036 13982
rect 8092 13972 8148 14700
rect 6972 13918 6974 13970
rect 7026 13918 7028 13970
rect 6972 13906 7028 13918
rect 7532 13970 8148 13972
rect 7532 13918 7982 13970
rect 8034 13918 8148 13970
rect 7532 13916 8148 13918
rect 8428 14308 8484 14318
rect 7532 13746 7588 13916
rect 7980 13906 8036 13916
rect 7532 13694 7534 13746
rect 7586 13694 7588 13746
rect 7532 13682 7588 13694
rect 6636 13570 6692 13580
rect 6748 13634 6804 13646
rect 6748 13582 6750 13634
rect 6802 13582 6804 13634
rect 6748 13524 6804 13582
rect 6748 13458 6804 13468
rect 7308 13524 7364 13534
rect 7308 13430 7364 13468
rect 8428 13076 8484 14252
rect 8876 13972 8932 13982
rect 8876 13878 8932 13916
rect 8764 13860 8820 13870
rect 8764 13766 8820 13804
rect 8988 13858 9044 15148
rect 9996 15092 10164 15148
rect 10220 15204 10276 15242
rect 10220 15138 10276 15148
rect 9884 14642 9940 14654
rect 9884 14590 9886 14642
rect 9938 14590 9940 14642
rect 9884 14532 9940 14590
rect 9884 14466 9940 14476
rect 9548 13972 9604 13982
rect 9548 13878 9604 13916
rect 8988 13806 8990 13858
rect 9042 13806 9044 13858
rect 8988 13794 9044 13806
rect 9884 13748 9940 13758
rect 9996 13748 10052 15092
rect 10332 14868 10388 15260
rect 9884 13746 10052 13748
rect 9884 13694 9886 13746
rect 9938 13694 10052 13746
rect 9884 13692 10052 13694
rect 10108 14812 10388 14868
rect 10108 13746 10164 14812
rect 10220 14644 10276 14654
rect 10220 14550 10276 14588
rect 10332 14420 10388 14430
rect 10332 14326 10388 14364
rect 10444 14196 10500 15708
rect 10780 15316 10836 17052
rect 11116 16884 11172 16894
rect 10780 15314 11060 15316
rect 10780 15262 10782 15314
rect 10834 15262 11060 15314
rect 10780 15260 11060 15262
rect 10780 15250 10836 15260
rect 10892 14532 10948 14542
rect 10668 14476 10892 14532
rect 10108 13694 10110 13746
rect 10162 13694 10164 13746
rect 9884 13682 9940 13692
rect 10108 13682 10164 13694
rect 10220 14140 10500 14196
rect 10556 14418 10612 14430
rect 10556 14366 10558 14418
rect 10610 14366 10612 14418
rect 9772 13524 9828 13534
rect 8428 13074 8932 13076
rect 8428 13022 8430 13074
rect 8482 13022 8932 13074
rect 8428 13020 8932 13022
rect 8428 13010 8484 13020
rect 6076 12798 6078 12850
rect 6130 12798 6132 12850
rect 5068 12740 5124 12750
rect 5068 12646 5124 12684
rect 5740 12738 5796 12750
rect 5740 12686 5742 12738
rect 5794 12686 5796 12738
rect 4620 12014 4622 12066
rect 4674 12014 4676 12066
rect 4620 12002 4676 12014
rect 5068 12460 5684 12516
rect 3164 11788 3444 11844
rect 2492 10770 2548 10780
rect 2828 11172 2884 11182
rect 2828 10722 2884 11116
rect 2828 10670 2830 10722
rect 2882 10670 2884 10722
rect 2828 10658 2884 10670
rect 2492 9716 2548 9726
rect 2492 9714 2660 9716
rect 2492 9662 2494 9714
rect 2546 9662 2660 9714
rect 2492 9660 2660 9662
rect 2492 9650 2548 9660
rect 2268 9214 2270 9266
rect 2322 9214 2324 9266
rect 2268 8036 2324 9214
rect 2604 8930 2660 9660
rect 2604 8878 2606 8930
rect 2658 8878 2660 8930
rect 2604 8866 2660 8878
rect 2716 9154 2772 9166
rect 2716 9102 2718 9154
rect 2770 9102 2772 9154
rect 2716 8428 2772 9102
rect 2940 8820 2996 8830
rect 2940 8818 3332 8820
rect 2940 8766 2942 8818
rect 2994 8766 3332 8818
rect 2940 8764 3332 8766
rect 2940 8754 2996 8764
rect 2716 8372 3108 8428
rect 3052 8258 3108 8372
rect 3276 8372 3332 8764
rect 3276 8306 3332 8316
rect 3052 8206 3054 8258
rect 3106 8206 3108 8258
rect 3052 8148 3108 8206
rect 3052 8082 3108 8092
rect 2604 8036 2660 8046
rect 2268 8034 2660 8036
rect 2268 7982 2270 8034
rect 2322 7982 2606 8034
rect 2658 7982 2660 8034
rect 2268 7980 2660 7982
rect 2268 7970 2324 7980
rect 2492 6916 2548 6926
rect 2492 6018 2548 6860
rect 2604 6804 2660 7980
rect 2604 6738 2660 6748
rect 2828 8034 2884 8046
rect 2828 7982 2830 8034
rect 2882 7982 2884 8034
rect 2828 6692 2884 7982
rect 2940 8034 2996 8046
rect 2940 7982 2942 8034
rect 2994 7982 2996 8034
rect 2940 7588 2996 7982
rect 3388 8036 3444 11788
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11396 4900 11406
rect 4508 11284 4564 11294
rect 4508 11190 4564 11228
rect 4620 11172 4676 11182
rect 4620 11078 4676 11116
rect 4844 10500 4900 11340
rect 5068 11394 5124 12460
rect 5628 12402 5684 12460
rect 5628 12350 5630 12402
rect 5682 12350 5684 12402
rect 5628 12338 5684 12350
rect 5740 12404 5796 12686
rect 6076 12628 6132 12798
rect 6076 12562 6132 12572
rect 6524 12740 6580 12750
rect 5740 12348 5908 12404
rect 5068 11342 5070 11394
rect 5122 11342 5124 11394
rect 5068 11330 5124 11342
rect 5516 12292 5572 12302
rect 5516 11284 5572 12236
rect 5740 12180 5796 12190
rect 5740 12086 5796 12124
rect 5292 10836 5348 10846
rect 4956 10500 5012 10510
rect 4844 10498 5012 10500
rect 4844 10446 4958 10498
rect 5010 10446 5012 10498
rect 4844 10444 5012 10446
rect 4956 10434 5012 10444
rect 5292 10498 5348 10780
rect 5404 10836 5460 10846
rect 5516 10836 5572 11228
rect 5852 11172 5908 12348
rect 5404 10834 5572 10836
rect 5404 10782 5406 10834
rect 5458 10782 5572 10834
rect 5404 10780 5572 10782
rect 5628 11116 5908 11172
rect 5964 12180 6020 12190
rect 5964 11396 6020 12124
rect 6188 12178 6244 12190
rect 6188 12126 6190 12178
rect 6242 12126 6244 12178
rect 6188 11844 6244 12126
rect 6188 11778 6244 11788
rect 6412 12178 6468 12190
rect 6412 12126 6414 12178
rect 6466 12126 6468 12178
rect 6076 11506 6132 11518
rect 6076 11454 6078 11506
rect 6130 11454 6132 11506
rect 6076 11396 6132 11454
rect 6412 11396 6468 12126
rect 6076 11340 6468 11396
rect 5404 10770 5460 10780
rect 5628 10722 5684 11116
rect 5628 10670 5630 10722
rect 5682 10670 5684 10722
rect 5628 10658 5684 10670
rect 5964 10612 6020 11340
rect 6412 10722 6468 11340
rect 6412 10670 6414 10722
rect 6466 10670 6468 10722
rect 6412 10658 6468 10670
rect 6524 10722 6580 12684
rect 7532 12740 7588 12750
rect 7084 12292 7140 12302
rect 7308 12292 7364 12302
rect 7140 12290 7364 12292
rect 7140 12238 7310 12290
rect 7362 12238 7364 12290
rect 7140 12236 7364 12238
rect 6636 12180 6692 12190
rect 6636 12086 6692 12124
rect 7084 12178 7140 12236
rect 7308 12226 7364 12236
rect 7084 12126 7086 12178
rect 7138 12126 7140 12178
rect 7084 12114 7140 12126
rect 7532 12178 7588 12684
rect 7532 12126 7534 12178
rect 7586 12126 7588 12178
rect 7532 12114 7588 12126
rect 6860 12066 6916 12078
rect 6860 12014 6862 12066
rect 6914 12014 6916 12066
rect 6524 10670 6526 10722
rect 6578 10670 6580 10722
rect 6524 10658 6580 10670
rect 6748 11844 6804 11854
rect 6188 10612 6244 10622
rect 5964 10610 6244 10612
rect 5964 10558 6190 10610
rect 6242 10558 6244 10610
rect 5964 10556 6244 10558
rect 6188 10546 6244 10556
rect 5292 10446 5294 10498
rect 5346 10446 5348 10498
rect 5292 10434 5348 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 6748 10164 6804 11788
rect 6860 11284 6916 12014
rect 8876 11396 8932 13020
rect 9660 12404 9716 12414
rect 9548 12348 9660 12404
rect 9324 11396 9380 11406
rect 8876 11394 9380 11396
rect 8876 11342 8878 11394
rect 8930 11342 9326 11394
rect 9378 11342 9380 11394
rect 8876 11340 9380 11342
rect 8876 11330 8932 11340
rect 9324 11330 9380 11340
rect 8204 11284 8260 11294
rect 6860 11228 7812 11284
rect 7756 10610 7812 11228
rect 8092 11282 8260 11284
rect 8092 11230 8206 11282
rect 8258 11230 8260 11282
rect 8092 11228 8260 11230
rect 7756 10558 7758 10610
rect 7810 10558 7812 10610
rect 7756 10546 7812 10558
rect 7980 10724 8036 10734
rect 7980 10610 8036 10668
rect 8092 10722 8148 11228
rect 8204 11218 8260 11228
rect 8092 10670 8094 10722
rect 8146 10670 8148 10722
rect 8092 10658 8148 10670
rect 8540 10724 8596 10734
rect 8540 10630 8596 10668
rect 7980 10558 7982 10610
rect 8034 10558 8036 10610
rect 7980 10546 8036 10558
rect 9436 10500 9492 10510
rect 6972 10388 7028 10398
rect 7644 10388 7700 10398
rect 6972 10386 7812 10388
rect 6972 10334 6974 10386
rect 7026 10334 7646 10386
rect 7698 10334 7812 10386
rect 6972 10332 7812 10334
rect 6972 10322 7028 10332
rect 7644 10322 7700 10332
rect 6748 10108 7140 10164
rect 4620 9940 4676 9950
rect 4620 9938 4900 9940
rect 4620 9886 4622 9938
rect 4674 9886 4900 9938
rect 4620 9884 4900 9886
rect 4620 9874 4676 9884
rect 3612 8930 3668 8942
rect 3612 8878 3614 8930
rect 3666 8878 3668 8930
rect 3612 8484 3668 8878
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4844 8428 4900 9884
rect 7084 9828 7140 10108
rect 7084 9734 7140 9772
rect 7532 9604 7588 9614
rect 7532 9510 7588 9548
rect 7644 9602 7700 9614
rect 7644 9550 7646 9602
rect 7698 9550 7700 9602
rect 7644 9156 7700 9550
rect 7756 9602 7812 10332
rect 9436 9938 9492 10444
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 8764 9828 8820 9838
rect 8764 9826 9268 9828
rect 8764 9774 8766 9826
rect 8818 9774 9268 9826
rect 8764 9772 9268 9774
rect 8764 9762 8820 9772
rect 7756 9550 7758 9602
rect 7810 9550 7812 9602
rect 7756 9492 7812 9550
rect 7756 9426 7812 9436
rect 8428 9604 8484 9614
rect 7644 9090 7700 9100
rect 3500 8372 3556 8382
rect 3500 8278 3556 8316
rect 3612 8260 3668 8428
rect 3612 8194 3668 8204
rect 3724 8372 4900 8428
rect 3500 8036 3556 8046
rect 3388 8034 3500 8036
rect 3388 7982 3390 8034
rect 3442 7982 3500 8034
rect 3388 7980 3500 7982
rect 3388 7942 3444 7980
rect 3500 7970 3556 7980
rect 3612 8036 3668 8046
rect 3724 8036 3780 8372
rect 4844 8370 4900 8372
rect 4844 8318 4846 8370
rect 4898 8318 4900 8370
rect 4844 8306 4900 8318
rect 6412 8932 6468 8942
rect 6412 8370 6468 8876
rect 8428 8596 8484 9548
rect 8540 9042 8596 9054
rect 8540 8990 8542 9042
rect 8594 8990 8596 9042
rect 8540 8932 8596 8990
rect 9100 9044 9156 9054
rect 8988 8932 9044 8942
rect 8540 8930 9044 8932
rect 8540 8878 8990 8930
rect 9042 8878 9044 8930
rect 8540 8876 9044 8878
rect 8428 8428 8484 8540
rect 8876 8708 8932 8718
rect 8428 8372 8596 8428
rect 6412 8318 6414 8370
rect 6466 8318 6468 8370
rect 6412 8306 6468 8318
rect 8540 8370 8596 8372
rect 8540 8318 8542 8370
rect 8594 8318 8596 8370
rect 8540 8306 8596 8318
rect 4060 8258 4116 8270
rect 4060 8206 4062 8258
rect 4114 8206 4116 8258
rect 3612 8034 3780 8036
rect 3612 7982 3614 8034
rect 3666 7982 3780 8034
rect 3612 7980 3780 7982
rect 3948 8148 4004 8158
rect 3612 7970 3668 7980
rect 2940 7522 2996 7532
rect 3836 7364 3892 7374
rect 3836 7270 3892 7308
rect 3836 6916 3892 6926
rect 3948 6916 4004 8092
rect 3836 6914 4004 6916
rect 3836 6862 3838 6914
rect 3890 6862 4004 6914
rect 3836 6860 4004 6862
rect 3836 6850 3892 6860
rect 3276 6804 3332 6814
rect 3276 6710 3332 6748
rect 4060 6804 4116 8206
rect 4508 8260 4564 8270
rect 4284 8148 4340 8158
rect 4284 8054 4340 8092
rect 4508 7476 4564 8204
rect 4620 8258 4676 8270
rect 4620 8206 4622 8258
rect 4674 8206 4676 8258
rect 4620 8036 4676 8206
rect 4620 7970 4676 7980
rect 5628 8258 5684 8270
rect 5628 8206 5630 8258
rect 5682 8206 5684 8258
rect 4956 7588 5012 7598
rect 4956 7494 5012 7532
rect 5180 7586 5236 7598
rect 5180 7534 5182 7586
rect 5234 7534 5236 7586
rect 4508 7382 4564 7420
rect 5068 7364 5124 7374
rect 5068 7270 5124 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4060 6738 4116 6748
rect 4396 6804 4452 6814
rect 2828 6626 2884 6636
rect 3612 6692 3668 6702
rect 3612 6598 3668 6636
rect 4172 6692 4228 6702
rect 4172 6598 4228 6636
rect 4396 6690 4452 6748
rect 4956 6804 5012 6814
rect 4956 6710 5012 6748
rect 4396 6638 4398 6690
rect 4450 6638 4452 6690
rect 4396 6626 4452 6638
rect 5068 6692 5124 6702
rect 5180 6692 5236 7534
rect 5628 7476 5684 8206
rect 8876 8260 8932 8652
rect 8988 8484 9044 8876
rect 8988 8418 9044 8428
rect 8876 8204 9044 8260
rect 5628 7382 5684 7420
rect 8876 8034 8932 8046
rect 8876 7982 8878 8034
rect 8930 7982 8932 8034
rect 6412 7362 6468 7374
rect 6412 7310 6414 7362
rect 6466 7310 6468 7362
rect 5740 6916 5796 6926
rect 5628 6804 5684 6814
rect 5628 6710 5684 6748
rect 5740 6802 5796 6860
rect 5740 6750 5742 6802
rect 5794 6750 5796 6802
rect 5740 6738 5796 6750
rect 6412 6802 6468 7310
rect 6412 6750 6414 6802
rect 6466 6750 6468 6802
rect 6412 6738 6468 6750
rect 8540 7362 8596 7374
rect 8540 7310 8542 7362
rect 8594 7310 8596 7362
rect 5124 6636 5236 6692
rect 5068 6598 5124 6636
rect 4844 6468 4900 6478
rect 4844 6466 5012 6468
rect 4844 6414 4846 6466
rect 4898 6414 5012 6466
rect 4844 6412 5012 6414
rect 4844 6402 4900 6412
rect 2492 5966 2494 6018
rect 2546 5966 2548 6018
rect 2492 5954 2548 5966
rect 4956 5908 5012 6412
rect 1820 5854 1822 5906
rect 1874 5854 1876 5906
rect 1820 5842 1876 5854
rect 4620 5906 5012 5908
rect 4620 5854 4958 5906
rect 5010 5854 5012 5906
rect 4620 5852 5012 5854
rect 4620 5794 4676 5852
rect 4956 5842 5012 5852
rect 5180 5906 5236 6636
rect 5964 6692 6020 6702
rect 6188 6692 6244 6702
rect 5964 6690 6244 6692
rect 5964 6638 5966 6690
rect 6018 6638 6190 6690
rect 6242 6638 6244 6690
rect 5964 6636 6244 6638
rect 5964 6626 6020 6636
rect 6188 6132 6244 6636
rect 6860 6692 6916 6702
rect 7308 6692 7364 6702
rect 6860 6690 7364 6692
rect 6860 6638 6862 6690
rect 6914 6638 7310 6690
rect 7362 6638 7364 6690
rect 6860 6636 7364 6638
rect 6860 6626 6916 6636
rect 7308 6626 7364 6636
rect 7868 6690 7924 6702
rect 7868 6638 7870 6690
rect 7922 6638 7924 6690
rect 6188 6038 6244 6076
rect 6636 6578 6692 6590
rect 6636 6526 6638 6578
rect 6690 6526 6692 6578
rect 6636 6468 6692 6526
rect 5180 5854 5182 5906
rect 5234 5854 5236 5906
rect 5180 5842 5236 5854
rect 5964 5906 6020 5918
rect 5964 5854 5966 5906
rect 6018 5854 6020 5906
rect 4620 5742 4622 5794
rect 4674 5742 4676 5794
rect 4620 5730 4676 5742
rect 4844 5684 4900 5694
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4172 5236 4228 5246
rect 4172 4226 4228 5180
rect 4844 5122 4900 5628
rect 5516 5684 5572 5694
rect 5516 5590 5572 5628
rect 5964 5684 6020 5854
rect 5964 5618 6020 5628
rect 4844 5070 4846 5122
rect 4898 5070 4900 5122
rect 4844 5058 4900 5070
rect 4956 5572 5012 5582
rect 4956 5010 5012 5516
rect 6636 5572 6692 6412
rect 7196 6466 7252 6478
rect 7196 6414 7198 6466
rect 7250 6414 7252 6466
rect 7084 6244 7140 6254
rect 7084 5906 7140 6188
rect 7196 6244 7252 6414
rect 7420 6468 7476 6478
rect 7420 6374 7476 6412
rect 7196 6188 7588 6244
rect 7196 6132 7252 6188
rect 7196 6066 7252 6076
rect 7084 5854 7086 5906
rect 7138 5854 7140 5906
rect 7084 5842 7140 5854
rect 7196 5906 7252 5918
rect 7196 5854 7198 5906
rect 7250 5854 7252 5906
rect 6636 5506 6692 5516
rect 7084 5572 7140 5582
rect 7196 5572 7252 5854
rect 7140 5516 7252 5572
rect 7308 5906 7364 5918
rect 7308 5854 7310 5906
rect 7362 5854 7364 5906
rect 7084 5506 7140 5516
rect 6300 5236 6356 5246
rect 5180 5124 5236 5134
rect 5180 5030 5236 5068
rect 6076 5124 6132 5134
rect 6076 5030 6132 5068
rect 6300 5122 6356 5180
rect 7308 5236 7364 5854
rect 7532 5906 7588 6188
rect 7868 6020 7924 6638
rect 8204 6692 8260 6702
rect 8540 6692 8596 7310
rect 8876 6804 8932 7982
rect 8988 7364 9044 8204
rect 9100 7476 9156 8988
rect 9212 7588 9268 9772
rect 9436 9492 9492 9502
rect 9436 9044 9492 9436
rect 9324 9042 9492 9044
rect 9324 8990 9438 9042
rect 9490 8990 9492 9042
rect 9324 8988 9492 8990
rect 9324 8258 9380 8988
rect 9436 8978 9492 8988
rect 9548 9044 9604 12348
rect 9660 12310 9716 12348
rect 9772 12292 9828 13468
rect 10108 12404 10164 12414
rect 10220 12404 10276 14140
rect 10444 13972 10500 13982
rect 10444 13878 10500 13916
rect 10556 13970 10612 14366
rect 10556 13918 10558 13970
rect 10610 13918 10612 13970
rect 10556 13906 10612 13918
rect 10668 13970 10724 14476
rect 10892 14438 10948 14476
rect 10668 13918 10670 13970
rect 10722 13918 10724 13970
rect 10668 13906 10724 13918
rect 11004 13748 11060 15260
rect 11116 15314 11172 16828
rect 11228 16772 11284 18174
rect 11228 16706 11284 16716
rect 11228 16324 11284 16334
rect 11340 16324 11396 18732
rect 11228 16322 11396 16324
rect 11228 16270 11230 16322
rect 11282 16270 11396 16322
rect 11228 16268 11396 16270
rect 11564 16996 11620 17006
rect 11564 16322 11620 16940
rect 11564 16270 11566 16322
rect 11618 16270 11620 16322
rect 11228 16100 11284 16268
rect 11564 16258 11620 16270
rect 11228 16034 11284 16044
rect 11116 15262 11118 15314
rect 11170 15262 11172 15314
rect 11116 15250 11172 15262
rect 11116 14530 11172 14542
rect 11116 14478 11118 14530
rect 11170 14478 11172 14530
rect 11116 13972 11172 14478
rect 11452 14308 11508 14318
rect 11452 14306 11620 14308
rect 11452 14254 11454 14306
rect 11506 14254 11620 14306
rect 11452 14252 11620 14254
rect 11452 14242 11508 14252
rect 11116 13906 11172 13916
rect 11452 13972 11508 13982
rect 11452 13878 11508 13916
rect 11564 13860 11620 14252
rect 11564 13766 11620 13804
rect 11116 13748 11172 13758
rect 11004 13692 11116 13748
rect 11116 13654 11172 13692
rect 11452 13522 11508 13534
rect 11452 13470 11454 13522
rect 11506 13470 11508 13522
rect 10164 12348 10276 12404
rect 11340 12404 11396 12414
rect 10108 12310 10164 12348
rect 9772 12236 9940 12292
rect 9548 8978 9604 8988
rect 9772 9042 9828 9054
rect 9772 8990 9774 9042
rect 9826 8990 9828 9042
rect 9660 8932 9716 8942
rect 9660 8838 9716 8876
rect 9324 8206 9326 8258
rect 9378 8206 9380 8258
rect 9324 8194 9380 8206
rect 9436 8596 9492 8606
rect 9772 8596 9828 8990
rect 9492 8540 9828 8596
rect 9884 8932 9940 12236
rect 11340 12178 11396 12348
rect 11340 12126 11342 12178
rect 11394 12126 11396 12178
rect 11340 12114 11396 12126
rect 10108 12066 10164 12078
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 10108 11506 10164 12014
rect 10332 12068 10388 12078
rect 10668 12068 10724 12078
rect 10332 12066 10724 12068
rect 10332 12014 10334 12066
rect 10386 12014 10670 12066
rect 10722 12014 10724 12066
rect 10332 12012 10724 12014
rect 10332 12002 10388 12012
rect 10668 12002 10724 12012
rect 11452 12066 11508 13470
rect 11452 12014 11454 12066
rect 11506 12014 11508 12066
rect 11452 12002 11508 12014
rect 10108 11454 10110 11506
rect 10162 11454 10164 11506
rect 10108 11442 10164 11454
rect 11340 10780 11620 10836
rect 11228 10724 11284 10734
rect 11340 10724 11396 10780
rect 11228 10722 11396 10724
rect 11228 10670 11230 10722
rect 11282 10670 11396 10722
rect 11228 10668 11396 10670
rect 10892 10612 10948 10622
rect 10892 10518 10948 10556
rect 11004 10500 11060 10510
rect 11004 10406 11060 10444
rect 11228 9268 11284 10668
rect 11452 10610 11508 10622
rect 11452 10558 11454 10610
rect 11506 10558 11508 10610
rect 11452 9940 11508 10558
rect 11452 9874 11508 9884
rect 11564 9938 11620 10780
rect 11564 9886 11566 9938
rect 11618 9886 11620 9938
rect 11564 9874 11620 9886
rect 11228 9174 11284 9212
rect 10108 9156 10164 9166
rect 10108 9062 10164 9100
rect 11340 9156 11396 9166
rect 11676 9156 11732 28140
rect 11788 28084 11844 28094
rect 11900 28084 11956 28588
rect 12236 28578 12292 28588
rect 11788 28082 11956 28084
rect 11788 28030 11790 28082
rect 11842 28030 11956 28082
rect 11788 28028 11956 28030
rect 11788 28018 11844 28028
rect 11788 24610 11844 24622
rect 11788 24558 11790 24610
rect 11842 24558 11844 24610
rect 11788 24276 11844 24558
rect 11788 24210 11844 24220
rect 11900 21364 11956 28028
rect 12124 28308 12180 28318
rect 12124 27970 12180 28252
rect 12124 27918 12126 27970
rect 12178 27918 12180 27970
rect 12124 27636 12180 27918
rect 12460 27860 12516 27870
rect 12124 27570 12180 27580
rect 12236 27804 12460 27860
rect 12236 27186 12292 27804
rect 12460 27766 12516 27804
rect 12236 27134 12238 27186
rect 12290 27134 12292 27186
rect 12236 27122 12292 27134
rect 12684 24836 12740 35532
rect 13020 35364 13076 36206
rect 13020 35298 13076 35308
rect 13020 34356 13076 34366
rect 13020 34262 13076 34300
rect 12796 34020 12852 34030
rect 12796 33458 12852 33964
rect 12796 33406 12798 33458
rect 12850 33406 12852 33458
rect 12796 33394 12852 33406
rect 12908 33124 12964 33134
rect 12908 33030 12964 33068
rect 13020 31554 13076 31566
rect 13020 31502 13022 31554
rect 13074 31502 13076 31554
rect 13020 31444 13076 31502
rect 13020 31378 13076 31388
rect 13020 28756 13076 28766
rect 13020 28662 13076 28700
rect 12796 27634 12852 27646
rect 12796 27582 12798 27634
rect 12850 27582 12852 27634
rect 12796 26908 12852 27582
rect 13132 26908 13188 36988
rect 13468 36482 13524 37212
rect 13804 37156 13860 38894
rect 13916 38164 13972 40908
rect 14140 39620 14196 39630
rect 14140 39526 14196 39564
rect 14028 39396 14084 39406
rect 14028 39060 14084 39340
rect 14140 39060 14196 39070
rect 14028 39058 14196 39060
rect 14028 39006 14142 39058
rect 14194 39006 14196 39058
rect 14028 39004 14196 39006
rect 14140 38994 14196 39004
rect 13916 38098 13972 38108
rect 14252 37940 14308 43484
rect 14364 42756 14420 44268
rect 15148 44098 15204 44110
rect 15148 44046 15150 44098
rect 15202 44046 15204 44098
rect 15148 43764 15204 44046
rect 15820 43708 15876 44382
rect 18172 44436 18228 45164
rect 20076 44436 20132 44446
rect 17500 44324 17556 44334
rect 17500 44230 17556 44268
rect 18172 44322 18228 44380
rect 19068 44434 20132 44436
rect 19068 44382 20078 44434
rect 20130 44382 20132 44434
rect 19068 44380 20132 44382
rect 18172 44270 18174 44322
rect 18226 44270 18228 44322
rect 18172 44258 18228 44270
rect 18732 44322 18788 44334
rect 18732 44270 18734 44322
rect 18786 44270 18788 44322
rect 16156 44210 16212 44222
rect 16156 44158 16158 44210
rect 16210 44158 16212 44210
rect 15036 43652 15204 43708
rect 15372 43652 15876 43708
rect 15932 44098 15988 44110
rect 15932 44046 15934 44098
rect 15986 44046 15988 44098
rect 14700 43426 14756 43438
rect 14700 43374 14702 43426
rect 14754 43374 14756 43426
rect 14700 42980 14756 43374
rect 14812 42980 14868 42990
rect 14700 42978 14868 42980
rect 14700 42926 14814 42978
rect 14866 42926 14868 42978
rect 14700 42924 14868 42926
rect 14812 42914 14868 42924
rect 14364 42690 14420 42700
rect 14924 42754 14980 42766
rect 14924 42702 14926 42754
rect 14978 42702 14980 42754
rect 14924 42084 14980 42702
rect 14476 42028 14980 42084
rect 14364 39620 14420 39630
rect 14364 39172 14420 39564
rect 14476 39396 14532 42028
rect 14924 41860 14980 41870
rect 15036 41860 15092 43652
rect 14980 41804 15092 41860
rect 15148 42756 15204 42766
rect 14924 41794 14980 41804
rect 14700 41300 14756 41310
rect 14700 41186 14756 41244
rect 14924 41300 14980 41310
rect 15148 41300 15204 42700
rect 15372 42754 15428 43652
rect 15932 43428 15988 44046
rect 16156 43708 16212 44158
rect 17948 44098 18004 44110
rect 17948 44046 17950 44098
rect 18002 44046 18004 44098
rect 17948 43876 18004 44046
rect 17948 43708 18004 43820
rect 18732 43708 18788 44270
rect 16156 43652 16660 43708
rect 17948 43652 18228 43708
rect 15932 43362 15988 43372
rect 15372 42702 15374 42754
rect 15426 42702 15428 42754
rect 15372 42690 15428 42702
rect 15820 42756 15876 42766
rect 15820 42662 15876 42700
rect 16492 42642 16548 42654
rect 16492 42590 16494 42642
rect 16546 42590 16548 42642
rect 15820 42196 15876 42206
rect 16380 42196 16436 42206
rect 16492 42196 16548 42590
rect 15820 42194 16324 42196
rect 15820 42142 15822 42194
rect 15874 42142 16324 42194
rect 15820 42140 16324 42142
rect 15820 42130 15876 42140
rect 15484 41970 15540 41982
rect 15484 41918 15486 41970
rect 15538 41918 15540 41970
rect 15484 41636 15540 41918
rect 15260 41300 15316 41310
rect 14924 41298 15316 41300
rect 14924 41246 14926 41298
rect 14978 41246 15262 41298
rect 15314 41246 15316 41298
rect 14924 41244 15316 41246
rect 14924 41234 14980 41244
rect 15260 41234 15316 41244
rect 14700 41134 14702 41186
rect 14754 41134 14756 41186
rect 14700 41122 14756 41134
rect 15036 40516 15092 40526
rect 14700 40460 15036 40516
rect 14700 40290 14756 40460
rect 15036 40422 15092 40460
rect 15484 40402 15540 41580
rect 15708 41970 15764 41982
rect 15708 41918 15710 41970
rect 15762 41918 15764 41970
rect 15596 41188 15652 41198
rect 15596 41094 15652 41132
rect 15708 41076 15764 41918
rect 15932 41970 15988 41982
rect 15932 41918 15934 41970
rect 15986 41918 15988 41970
rect 15820 41076 15876 41086
rect 15708 41074 15876 41076
rect 15708 41022 15822 41074
rect 15874 41022 15876 41074
rect 15708 41020 15876 41022
rect 15708 40516 15764 41020
rect 15820 41010 15876 41020
rect 15708 40422 15764 40460
rect 15820 40516 15876 40526
rect 15932 40516 15988 41918
rect 16268 41972 16324 42140
rect 16380 42194 16548 42196
rect 16380 42142 16382 42194
rect 16434 42142 16548 42194
rect 16380 42140 16548 42142
rect 16380 42130 16436 42140
rect 16492 41972 16548 41982
rect 16268 41970 16548 41972
rect 16268 41918 16494 41970
rect 16546 41918 16548 41970
rect 16268 41916 16548 41918
rect 16492 41906 16548 41916
rect 16268 41748 16324 41758
rect 16156 41524 16212 41534
rect 16156 41074 16212 41468
rect 16268 41298 16324 41692
rect 16268 41246 16270 41298
rect 16322 41246 16324 41298
rect 16268 41234 16324 41246
rect 16380 41748 16436 41758
rect 16604 41748 16660 43652
rect 17612 43538 17668 43550
rect 17612 43486 17614 43538
rect 17666 43486 17668 43538
rect 16828 43428 16884 43438
rect 16828 42084 16884 43372
rect 16828 42018 16884 42028
rect 17276 42420 17332 42430
rect 16380 41746 16660 41748
rect 16380 41694 16382 41746
rect 16434 41694 16660 41746
rect 16380 41692 16660 41694
rect 16716 41746 16772 41758
rect 16716 41694 16718 41746
rect 16770 41694 16772 41746
rect 16156 41022 16158 41074
rect 16210 41022 16212 41074
rect 16156 41010 16212 41022
rect 16268 40628 16324 40638
rect 16380 40628 16436 41692
rect 16268 40626 16436 40628
rect 16268 40574 16270 40626
rect 16322 40574 16436 40626
rect 16268 40572 16436 40574
rect 16492 41188 16548 41198
rect 16268 40562 16324 40572
rect 15820 40514 15988 40516
rect 15820 40462 15822 40514
rect 15874 40462 15988 40514
rect 15820 40460 15988 40462
rect 15484 40350 15486 40402
rect 15538 40350 15540 40402
rect 15484 40338 15540 40350
rect 14700 40238 14702 40290
rect 14754 40238 14756 40290
rect 14700 40226 14756 40238
rect 15148 40178 15204 40190
rect 15148 40126 15150 40178
rect 15202 40126 15204 40178
rect 15148 39620 15204 40126
rect 15708 39732 15764 39742
rect 15820 39732 15876 40460
rect 15708 39730 16212 39732
rect 15708 39678 15710 39730
rect 15762 39678 16212 39730
rect 15708 39676 16212 39678
rect 15484 39620 15540 39630
rect 15148 39564 15484 39620
rect 15484 39526 15540 39564
rect 14588 39508 14644 39518
rect 14812 39508 14868 39518
rect 14644 39506 14868 39508
rect 14644 39454 14814 39506
rect 14866 39454 14868 39506
rect 14644 39452 14868 39454
rect 14588 39442 14644 39452
rect 14812 39442 14868 39452
rect 14476 39302 14532 39340
rect 15260 39396 15316 39406
rect 14364 39116 14532 39172
rect 14476 38834 14532 39116
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14252 37874 14308 37884
rect 14364 38724 14420 38734
rect 14364 37716 14420 38668
rect 14476 38668 14532 38782
rect 15148 38724 15204 38734
rect 14476 38612 14644 38668
rect 15148 38630 15204 38668
rect 15260 38724 15316 39340
rect 15596 38836 15652 38846
rect 15484 38780 15596 38836
rect 15260 38722 15428 38724
rect 15260 38670 15262 38722
rect 15314 38670 15428 38722
rect 15260 38668 15428 38670
rect 15260 38658 15316 38668
rect 14252 37660 14420 37716
rect 14252 37378 14308 37660
rect 14252 37326 14254 37378
rect 14306 37326 14308 37378
rect 14252 37314 14308 37326
rect 13804 37100 14308 37156
rect 14252 36594 14308 37100
rect 14252 36542 14254 36594
rect 14306 36542 14308 36594
rect 14252 36530 14308 36542
rect 13468 36430 13470 36482
rect 13522 36430 13524 36482
rect 13468 36372 13524 36430
rect 13468 36306 13524 36316
rect 14588 36260 14644 38612
rect 14588 36194 14644 36204
rect 14700 38052 14756 38062
rect 14700 35698 14756 37996
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 13692 35028 13748 35038
rect 13692 34934 13748 34972
rect 13804 34468 13860 34478
rect 13804 34354 13860 34412
rect 13804 34302 13806 34354
rect 13858 34302 13860 34354
rect 13804 34290 13860 34302
rect 14700 34356 14756 35646
rect 15372 35698 15428 38668
rect 15484 38722 15540 38780
rect 15596 38770 15652 38780
rect 15708 38834 15764 39676
rect 16156 39506 16212 39676
rect 16156 39454 16158 39506
rect 16210 39454 16212 39506
rect 16156 39442 16212 39454
rect 16492 39394 16548 41132
rect 16716 40852 16772 41694
rect 17276 41186 17332 42364
rect 17500 42084 17556 42094
rect 17612 42084 17668 43486
rect 17556 42028 17668 42084
rect 17836 43426 17892 43438
rect 17836 43374 17838 43426
rect 17890 43374 17892 43426
rect 17500 41990 17556 42028
rect 17276 41134 17278 41186
rect 17330 41134 17332 41186
rect 17276 41122 17332 41134
rect 17388 41636 17444 41646
rect 16604 40796 16772 40852
rect 16604 39508 16660 40796
rect 16716 40628 16772 40638
rect 16716 40626 16996 40628
rect 16716 40574 16718 40626
rect 16770 40574 16996 40626
rect 16716 40572 16996 40574
rect 16716 40562 16772 40572
rect 16828 40402 16884 40414
rect 16828 40350 16830 40402
rect 16882 40350 16884 40402
rect 16604 39442 16660 39452
rect 16716 40178 16772 40190
rect 16716 40126 16718 40178
rect 16770 40126 16772 40178
rect 16492 39342 16494 39394
rect 16546 39342 16548 39394
rect 16492 39172 16548 39342
rect 16716 39396 16772 40126
rect 16828 39396 16884 40350
rect 16940 39620 16996 40572
rect 17276 39730 17332 39742
rect 17276 39678 17278 39730
rect 17330 39678 17332 39730
rect 17164 39620 17220 39630
rect 16996 39618 17220 39620
rect 16996 39566 17166 39618
rect 17218 39566 17220 39618
rect 16996 39564 17220 39566
rect 16940 39526 16996 39564
rect 17164 39554 17220 39564
rect 17276 39396 17332 39678
rect 16828 39340 17332 39396
rect 16716 39330 16772 39340
rect 16492 39116 16772 39172
rect 16604 38946 16660 38958
rect 16604 38894 16606 38946
rect 16658 38894 16660 38946
rect 15708 38782 15710 38834
rect 15762 38782 15764 38834
rect 15708 38770 15764 38782
rect 16044 38836 16100 38846
rect 16492 38836 16548 38846
rect 16044 38834 16324 38836
rect 16044 38782 16046 38834
rect 16098 38782 16324 38834
rect 16044 38780 16324 38782
rect 16044 38770 16100 38780
rect 15484 38670 15486 38722
rect 15538 38670 15540 38722
rect 15484 38658 15540 38670
rect 16156 38612 16212 38622
rect 16156 38518 16212 38556
rect 16268 38500 16324 38780
rect 16492 38722 16548 38780
rect 16492 38670 16494 38722
rect 16546 38670 16548 38722
rect 16492 38658 16548 38670
rect 16604 38500 16660 38894
rect 16268 38444 16660 38500
rect 16380 37156 16436 37166
rect 16604 37156 16660 38444
rect 16716 37828 16772 39116
rect 16716 37762 16772 37772
rect 16828 38722 16884 38734
rect 16828 38670 16830 38722
rect 16882 38670 16884 38722
rect 16436 37100 16660 37156
rect 16380 37062 16436 37100
rect 16380 36594 16436 36606
rect 16380 36542 16382 36594
rect 16434 36542 16436 36594
rect 15372 35646 15374 35698
rect 15426 35646 15428 35698
rect 15372 35634 15428 35646
rect 15596 36148 15652 36158
rect 15596 35698 15652 36092
rect 16380 36036 16436 36542
rect 16716 36482 16772 36494
rect 16716 36430 16718 36482
rect 16770 36430 16772 36482
rect 16436 35980 16548 36036
rect 16380 35970 16436 35980
rect 15708 35924 15764 35934
rect 15708 35922 15876 35924
rect 15708 35870 15710 35922
rect 15762 35870 15876 35922
rect 15708 35868 15876 35870
rect 15708 35858 15764 35868
rect 15596 35646 15598 35698
rect 15650 35646 15652 35698
rect 15596 35634 15652 35646
rect 15708 35700 15764 35710
rect 15708 35606 15764 35644
rect 15820 35026 15876 35868
rect 16492 35922 16548 35980
rect 16492 35870 16494 35922
rect 16546 35870 16548 35922
rect 16492 35858 16548 35870
rect 15820 34974 15822 35026
rect 15874 34974 15876 35026
rect 15820 34962 15876 34974
rect 15932 35364 15988 35374
rect 14700 34290 14756 34300
rect 14924 34468 14980 34478
rect 14924 34354 14980 34412
rect 14924 34302 14926 34354
rect 14978 34302 14980 34354
rect 13580 34244 13636 34254
rect 13356 34132 13412 34142
rect 13356 34038 13412 34076
rect 13580 34130 13636 34188
rect 13580 34078 13582 34130
rect 13634 34078 13636 34130
rect 13468 33346 13524 33358
rect 13468 33294 13470 33346
rect 13522 33294 13524 33346
rect 13468 31892 13524 33294
rect 13356 31836 13524 31892
rect 13356 30996 13412 31836
rect 13468 31668 13524 31678
rect 13468 31574 13524 31612
rect 13580 31556 13636 34078
rect 13916 34130 13972 34142
rect 13916 34078 13918 34130
rect 13970 34078 13972 34130
rect 13692 34020 13748 34030
rect 13692 33926 13748 33964
rect 13916 33908 13972 34078
rect 14588 34018 14644 34030
rect 14588 33966 14590 34018
rect 14642 33966 14644 34018
rect 13916 33842 13972 33852
rect 14476 33908 14532 33918
rect 14252 33236 14308 33246
rect 14252 33142 14308 33180
rect 14028 33124 14084 33134
rect 14028 32674 14084 33068
rect 14028 32622 14030 32674
rect 14082 32622 14084 32674
rect 14028 32610 14084 32622
rect 13916 31892 13972 31902
rect 13916 31778 13972 31836
rect 13916 31726 13918 31778
rect 13970 31726 13972 31778
rect 13916 31714 13972 31726
rect 14140 31778 14196 31790
rect 14140 31726 14142 31778
rect 14194 31726 14196 31778
rect 13692 31556 13748 31566
rect 13580 31554 13748 31556
rect 13580 31502 13694 31554
rect 13746 31502 13748 31554
rect 13580 31500 13748 31502
rect 13692 31220 13748 31500
rect 13804 31556 13860 31566
rect 13804 31462 13860 31500
rect 14140 31444 14196 31726
rect 14476 31666 14532 33852
rect 14476 31614 14478 31666
rect 14530 31614 14532 31666
rect 14476 31602 14532 31614
rect 14588 31892 14644 33966
rect 14924 34020 14980 34302
rect 15260 34020 15316 34030
rect 15484 34020 15540 34030
rect 14924 33964 15204 34020
rect 14812 32564 14868 32574
rect 14812 32470 14868 32508
rect 14140 31378 14196 31388
rect 14588 31332 14644 31836
rect 14812 31554 14868 31566
rect 14812 31502 14814 31554
rect 14866 31502 14868 31554
rect 14812 31444 14868 31502
rect 15148 31556 15204 33964
rect 15316 34018 15540 34020
rect 15316 33966 15486 34018
rect 15538 33966 15540 34018
rect 15316 33964 15540 33966
rect 15260 31780 15316 33964
rect 15484 33954 15540 33964
rect 15932 34018 15988 35308
rect 16716 35028 16772 36430
rect 16828 36148 16884 38670
rect 17164 38500 17220 38510
rect 17276 38500 17332 39340
rect 17388 39058 17444 41580
rect 17836 41412 17892 43374
rect 17948 43316 18004 43326
rect 17948 43314 18116 43316
rect 17948 43262 17950 43314
rect 18002 43262 18116 43314
rect 17948 43260 18116 43262
rect 17948 43250 18004 43260
rect 18060 41972 18116 43260
rect 18172 42532 18228 43652
rect 18508 43652 18788 43708
rect 18396 43538 18452 43550
rect 18396 43486 18398 43538
rect 18450 43486 18452 43538
rect 18396 42756 18452 43486
rect 18396 42690 18452 42700
rect 18172 42466 18228 42476
rect 18060 41878 18116 41916
rect 18396 41970 18452 41982
rect 18396 41918 18398 41970
rect 18450 41918 18452 41970
rect 18172 41858 18228 41870
rect 18172 41806 18174 41858
rect 18226 41806 18228 41858
rect 17836 41346 17892 41356
rect 18060 41748 18116 41758
rect 18060 41300 18116 41692
rect 18060 41186 18116 41244
rect 18060 41134 18062 41186
rect 18114 41134 18116 41186
rect 18060 41122 18116 41134
rect 18172 41188 18228 41806
rect 18396 41636 18452 41918
rect 18396 41570 18452 41580
rect 18172 41122 18228 41132
rect 18396 41412 18452 41422
rect 18396 41186 18452 41356
rect 18396 41134 18398 41186
rect 18450 41134 18452 41186
rect 18396 41122 18452 41134
rect 17500 40514 17556 40526
rect 17500 40462 17502 40514
rect 17554 40462 17556 40514
rect 17500 40404 17556 40462
rect 17500 40338 17556 40348
rect 17612 40516 17668 40526
rect 17612 40290 17668 40460
rect 17612 40238 17614 40290
rect 17666 40238 17668 40290
rect 17612 40226 17668 40238
rect 17724 40180 17780 40190
rect 17724 40086 17780 40124
rect 18284 39842 18340 39854
rect 18284 39790 18286 39842
rect 18338 39790 18340 39842
rect 17388 39006 17390 39058
rect 17442 39006 17444 39058
rect 17388 38994 17444 39006
rect 18172 39618 18228 39630
rect 18172 39566 18174 39618
rect 18226 39566 18228 39618
rect 18060 38948 18116 38958
rect 17724 38836 17780 38846
rect 17724 38742 17780 38780
rect 17220 38444 17332 38500
rect 17164 38434 17220 38444
rect 17948 38052 18004 38062
rect 17500 37828 17556 37838
rect 17500 37490 17556 37772
rect 17500 37438 17502 37490
rect 17554 37438 17556 37490
rect 17500 37426 17556 37438
rect 17724 37604 17780 37614
rect 16940 37268 16996 37278
rect 16940 37174 16996 37212
rect 17724 37266 17780 37548
rect 17724 37214 17726 37266
rect 17778 37214 17780 37266
rect 17052 36708 17108 36718
rect 17052 36482 17108 36652
rect 17052 36430 17054 36482
rect 17106 36430 17108 36482
rect 17052 36418 17108 36430
rect 17388 36484 17444 36522
rect 17388 36418 17444 36428
rect 17612 36484 17668 36494
rect 17500 36372 17556 36382
rect 17164 36260 17220 36270
rect 16828 36082 16884 36092
rect 16940 36258 17220 36260
rect 16940 36206 17166 36258
rect 17218 36206 17220 36258
rect 16940 36204 17220 36206
rect 16940 36036 16996 36204
rect 17164 36194 17220 36204
rect 17276 36258 17332 36270
rect 17276 36206 17278 36258
rect 17330 36206 17332 36258
rect 16940 35970 16996 35980
rect 17164 36036 17220 36046
rect 17052 35924 17108 35934
rect 16828 35812 16884 35822
rect 16828 35718 16884 35756
rect 16940 35028 16996 35038
rect 16716 34972 16940 35028
rect 16604 34916 16660 34926
rect 16604 34822 16660 34860
rect 16940 34914 16996 34972
rect 16940 34862 16942 34914
rect 16994 34862 16996 34914
rect 16940 34850 16996 34862
rect 16492 34468 16548 34478
rect 16492 34354 16548 34412
rect 16492 34302 16494 34354
rect 16546 34302 16548 34354
rect 16492 34290 16548 34302
rect 17052 34356 17108 35868
rect 17052 34290 17108 34300
rect 15932 33966 15934 34018
rect 15986 33966 15988 34018
rect 15372 33236 15428 33246
rect 15372 32786 15428 33180
rect 15372 32734 15374 32786
rect 15426 32734 15428 32786
rect 15372 32722 15428 32734
rect 15596 32674 15652 32686
rect 15596 32622 15598 32674
rect 15650 32622 15652 32674
rect 15484 32564 15540 32574
rect 15596 32564 15652 32622
rect 15484 32562 15652 32564
rect 15484 32510 15486 32562
rect 15538 32510 15652 32562
rect 15484 32508 15652 32510
rect 15484 32498 15540 32508
rect 15260 31714 15316 31724
rect 15372 32004 15428 32014
rect 15148 31500 15316 31556
rect 14812 31378 14868 31388
rect 14588 31266 14644 31276
rect 13692 31164 14196 31220
rect 13356 30902 13412 30940
rect 14028 30996 14084 31006
rect 14028 30322 14084 30940
rect 14028 30270 14030 30322
rect 14082 30270 14084 30322
rect 13692 29316 13748 29326
rect 13692 29314 13860 29316
rect 13692 29262 13694 29314
rect 13746 29262 13860 29314
rect 13692 29260 13860 29262
rect 13692 29250 13748 29260
rect 13468 28420 13524 28430
rect 13244 27858 13300 27870
rect 13244 27806 13246 27858
rect 13298 27806 13300 27858
rect 13244 27188 13300 27806
rect 13356 27860 13412 27870
rect 13468 27860 13524 28364
rect 13804 28418 13860 29260
rect 13804 28366 13806 28418
rect 13858 28366 13860 28418
rect 13356 27858 13524 27860
rect 13356 27806 13358 27858
rect 13410 27806 13524 27858
rect 13356 27804 13524 27806
rect 13580 27860 13636 27870
rect 13356 27748 13412 27804
rect 13356 27682 13412 27692
rect 13244 27122 13300 27132
rect 13580 27076 13636 27804
rect 13804 27298 13860 28366
rect 13804 27246 13806 27298
rect 13858 27246 13860 27298
rect 13804 27234 13860 27246
rect 14028 27860 14084 30270
rect 14140 29538 14196 31164
rect 14700 31108 14756 31118
rect 14700 31014 14756 31052
rect 15260 30212 15316 31500
rect 15260 30146 15316 30156
rect 14140 29486 14142 29538
rect 14194 29486 14196 29538
rect 14140 29474 14196 29486
rect 14476 29426 14532 29438
rect 14476 29374 14478 29426
rect 14530 29374 14532 29426
rect 14476 29316 14532 29374
rect 14924 29428 14980 29438
rect 14924 29426 15092 29428
rect 14924 29374 14926 29426
rect 14978 29374 15092 29426
rect 14924 29372 15092 29374
rect 14924 29362 14980 29372
rect 14476 28756 14532 29260
rect 15036 29204 15092 29372
rect 15372 29426 15428 31948
rect 15820 31666 15876 31678
rect 15820 31614 15822 31666
rect 15874 31614 15876 31666
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15260 29204 15316 29214
rect 15036 29148 15260 29204
rect 15260 29138 15316 29148
rect 14476 28690 14532 28700
rect 14700 27972 14756 27982
rect 14700 27878 14756 27916
rect 13916 27188 13972 27198
rect 13916 27076 13972 27132
rect 13580 27010 13636 27020
rect 13804 27020 13972 27076
rect 12796 26852 12964 26908
rect 13132 26852 13748 26908
rect 12796 25620 12852 25630
rect 12796 25526 12852 25564
rect 12684 24780 12852 24836
rect 12684 24612 12740 24622
rect 12348 24164 12404 24174
rect 12348 24070 12404 24108
rect 12684 24162 12740 24556
rect 12684 24110 12686 24162
rect 12738 24110 12740 24162
rect 12684 24098 12740 24110
rect 12460 23938 12516 23950
rect 12460 23886 12462 23938
rect 12514 23886 12516 23938
rect 12012 23828 12068 23838
rect 12012 23734 12068 23772
rect 12460 23828 12516 23886
rect 12460 23762 12516 23772
rect 12796 22148 12852 24780
rect 12908 23940 12964 26852
rect 13692 26850 13748 26852
rect 13692 26798 13694 26850
rect 13746 26798 13748 26850
rect 13692 26786 13748 26798
rect 13580 26180 13636 26190
rect 13804 26180 13860 27020
rect 14028 26908 14084 27804
rect 14476 27748 14532 27758
rect 14140 27298 14196 27310
rect 14140 27246 14142 27298
rect 14194 27246 14196 27298
rect 14140 27074 14196 27246
rect 14140 27022 14142 27074
rect 14194 27022 14196 27074
rect 14140 27010 14196 27022
rect 14252 27076 14308 27086
rect 14252 26982 14308 27020
rect 13916 26852 14084 26908
rect 13916 26292 13972 26852
rect 13916 26198 13972 26236
rect 13580 26178 13860 26180
rect 13580 26126 13582 26178
rect 13634 26126 13860 26178
rect 13580 26124 13860 26126
rect 13580 26114 13636 26124
rect 13580 25506 13636 25518
rect 13580 25454 13582 25506
rect 13634 25454 13636 25506
rect 13580 24724 13636 25454
rect 14252 25394 14308 25406
rect 14252 25342 14254 25394
rect 14306 25342 14308 25394
rect 14252 25284 14308 25342
rect 14252 25218 14308 25228
rect 13580 24658 13636 24668
rect 14476 24722 14532 27692
rect 14588 27636 14644 27646
rect 14588 24836 14644 27580
rect 15036 27188 15092 27198
rect 14700 26180 14756 26190
rect 14700 26086 14756 26124
rect 14588 24780 14868 24836
rect 14476 24670 14478 24722
rect 14530 24670 14532 24722
rect 14476 24658 14532 24670
rect 14812 24722 14868 24780
rect 14812 24670 14814 24722
rect 14866 24670 14868 24722
rect 14812 24658 14868 24670
rect 15036 24722 15092 27132
rect 15372 26908 15428 29374
rect 15484 31554 15540 31566
rect 15484 31502 15486 31554
rect 15538 31502 15540 31554
rect 15484 31444 15540 31502
rect 15484 29204 15540 31388
rect 15708 31554 15764 31566
rect 15708 31502 15710 31554
rect 15762 31502 15764 31554
rect 15708 31108 15764 31502
rect 15708 31042 15764 31052
rect 15820 29652 15876 31614
rect 15820 29586 15876 29596
rect 15820 29316 15876 29326
rect 15820 29222 15876 29260
rect 15484 29138 15540 29148
rect 15484 27860 15540 27870
rect 15484 27074 15540 27804
rect 15932 27412 15988 33966
rect 16940 34018 16996 34030
rect 16940 33966 16942 34018
rect 16994 33966 16996 34018
rect 16940 33572 16996 33966
rect 17164 33908 17220 35980
rect 17276 35924 17332 36206
rect 17276 35858 17332 35868
rect 17388 36036 17444 36046
rect 17276 34692 17332 34702
rect 17276 34598 17332 34636
rect 17388 34354 17444 35980
rect 17500 35810 17556 36316
rect 17500 35758 17502 35810
rect 17554 35758 17556 35810
rect 17500 35746 17556 35758
rect 17612 35698 17668 36428
rect 17612 35646 17614 35698
rect 17666 35646 17668 35698
rect 17612 35364 17668 35646
rect 17724 35476 17780 37214
rect 17836 36258 17892 36270
rect 17836 36206 17838 36258
rect 17890 36206 17892 36258
rect 17836 36148 17892 36206
rect 17836 36082 17892 36092
rect 17948 36036 18004 37996
rect 17948 35970 18004 35980
rect 18060 38050 18116 38892
rect 18172 38276 18228 39566
rect 18284 39060 18340 39790
rect 18284 38994 18340 39004
rect 18396 39730 18452 39742
rect 18396 39678 18398 39730
rect 18450 39678 18452 39730
rect 18396 38724 18452 39678
rect 18396 38658 18452 38668
rect 18172 38210 18228 38220
rect 18060 37998 18062 38050
rect 18114 37998 18116 38050
rect 17948 35812 18004 35822
rect 17948 35698 18004 35756
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35634 18004 35646
rect 17724 35410 17780 35420
rect 17612 35298 17668 35308
rect 18060 35252 18116 37998
rect 18396 37378 18452 37390
rect 18396 37326 18398 37378
rect 18450 37326 18452 37378
rect 18172 37266 18228 37278
rect 18172 37214 18174 37266
rect 18226 37214 18228 37266
rect 18172 36148 18228 37214
rect 18396 36596 18452 37326
rect 18508 37380 18564 43652
rect 19068 43650 19124 44380
rect 20076 44370 20132 44380
rect 20412 44436 20468 44446
rect 20188 44212 20244 44222
rect 19292 44098 19348 44110
rect 19292 44046 19294 44098
rect 19346 44046 19348 44098
rect 19292 43764 19348 44046
rect 19852 44100 19908 44138
rect 20188 44118 20244 44156
rect 19852 44034 19908 44044
rect 20412 44100 20468 44380
rect 21980 44436 22036 44446
rect 21756 44324 21812 44334
rect 21756 44230 21812 44268
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19292 43652 19460 43708
rect 19068 43598 19070 43650
rect 19122 43598 19124 43650
rect 19068 43586 19124 43598
rect 19180 43428 19236 43438
rect 18620 42866 18676 42878
rect 18620 42814 18622 42866
rect 18674 42814 18676 42866
rect 18620 38836 18676 42814
rect 19180 42754 19236 43372
rect 19180 42702 19182 42754
rect 19234 42702 19236 42754
rect 19180 42420 19236 42702
rect 19180 42354 19236 42364
rect 19292 42866 19348 42878
rect 19292 42814 19294 42866
rect 19346 42814 19348 42866
rect 18844 42196 18900 42206
rect 18844 42194 19236 42196
rect 18844 42142 18846 42194
rect 18898 42142 19236 42194
rect 18844 42140 19236 42142
rect 18844 42130 18900 42140
rect 18956 40514 19012 40526
rect 18956 40462 18958 40514
rect 19010 40462 19012 40514
rect 18732 40402 18788 40414
rect 18732 40350 18734 40402
rect 18786 40350 18788 40402
rect 18732 39620 18788 40350
rect 18956 39844 19012 40462
rect 18956 39778 19012 39788
rect 19068 39620 19124 39630
rect 18732 39554 18788 39564
rect 18956 39618 19124 39620
rect 18956 39566 19070 39618
rect 19122 39566 19124 39618
rect 18956 39564 19124 39566
rect 18620 38724 18676 38780
rect 18732 38724 18788 38734
rect 18620 38722 18788 38724
rect 18620 38670 18734 38722
rect 18786 38670 18788 38722
rect 18620 38668 18788 38670
rect 18732 38658 18788 38668
rect 18508 37324 18900 37380
rect 18508 37156 18564 37166
rect 18508 37062 18564 37100
rect 18844 36596 18900 37324
rect 18956 37156 19012 39564
rect 19068 39554 19124 39564
rect 19180 38834 19236 42140
rect 19292 41748 19348 42814
rect 19292 41682 19348 41692
rect 19404 41970 19460 43652
rect 20076 42980 20132 42990
rect 20076 42886 20132 42924
rect 20412 42754 20468 44044
rect 20748 44210 20804 44222
rect 20748 44158 20750 44210
rect 20802 44158 20804 44210
rect 20748 43428 20804 44158
rect 21532 44210 21588 44222
rect 21532 44158 21534 44210
rect 21586 44158 21588 44210
rect 20860 44100 20916 44110
rect 20860 44006 20916 44044
rect 21084 44098 21140 44110
rect 21084 44046 21086 44098
rect 21138 44046 21140 44098
rect 21084 43652 21140 44046
rect 21532 43708 21588 44158
rect 21868 44212 21924 44222
rect 21868 44118 21924 44156
rect 21980 44098 22036 44380
rect 23100 44436 23156 44446
rect 23548 44436 23604 44446
rect 23100 44434 23604 44436
rect 23100 44382 23102 44434
rect 23154 44382 23550 44434
rect 23602 44382 23604 44434
rect 23100 44380 23604 44382
rect 23100 44370 23156 44380
rect 23548 44370 23604 44380
rect 27804 44434 27860 44446
rect 27804 44382 27806 44434
rect 27858 44382 27860 44434
rect 22428 44324 22484 44334
rect 21980 44046 21982 44098
rect 22034 44046 22036 44098
rect 21980 43876 22036 44046
rect 22092 44100 22148 44110
rect 22092 44006 22148 44044
rect 21980 43810 22036 43820
rect 21084 43586 21140 43596
rect 21196 43652 21588 43708
rect 22428 43764 22484 44268
rect 22764 44324 22820 44334
rect 22764 44230 22820 44268
rect 25004 44322 25060 44334
rect 25004 44270 25006 44322
rect 25058 44270 25060 44322
rect 22428 43698 22484 43708
rect 22540 44210 22596 44222
rect 22540 44158 22542 44210
rect 22594 44158 22596 44210
rect 21196 43428 21252 43652
rect 20748 43426 21252 43428
rect 20748 43374 21198 43426
rect 21250 43374 21252 43426
rect 20748 43372 21252 43374
rect 20412 42702 20414 42754
rect 20466 42702 20468 42754
rect 20412 42690 20468 42702
rect 20636 42756 20692 42766
rect 20748 42756 20804 43372
rect 21196 43362 21252 43372
rect 21644 43428 21700 43438
rect 21644 43334 21700 43372
rect 22540 43428 22596 44158
rect 22988 44098 23044 44110
rect 22988 44046 22990 44098
rect 23042 44046 23044 44098
rect 22652 43988 22708 43998
rect 22652 43708 22708 43932
rect 22988 43708 23044 44046
rect 23100 44100 23156 44110
rect 23156 44044 23380 44100
rect 23100 44006 23156 44044
rect 22652 43652 23044 43708
rect 22540 43362 22596 43372
rect 21868 42980 21924 42990
rect 20636 42754 20804 42756
rect 20636 42702 20638 42754
rect 20690 42702 20804 42754
rect 20636 42700 20804 42702
rect 21756 42866 21812 42878
rect 21756 42814 21758 42866
rect 21810 42814 21812 42866
rect 20636 42690 20692 42700
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 41918 19406 41970
rect 19458 41918 19460 41970
rect 19292 40292 19348 40302
rect 19292 39618 19348 40236
rect 19292 39566 19294 39618
rect 19346 39566 19348 39618
rect 19292 39172 19348 39566
rect 19292 39106 19348 39116
rect 19404 38948 19460 41918
rect 21308 41300 21364 41310
rect 21308 41298 21588 41300
rect 21308 41246 21310 41298
rect 21362 41246 21588 41298
rect 21308 41244 21588 41246
rect 21308 41234 21364 41244
rect 20412 41188 20468 41198
rect 20412 41094 20468 41132
rect 20636 41074 20692 41086
rect 20636 41022 20638 41074
rect 20690 41022 20692 41074
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20188 40516 20244 40526
rect 20188 40402 20244 40460
rect 20188 40350 20190 40402
rect 20242 40350 20244 40402
rect 20188 40338 20244 40350
rect 20076 39844 20132 39854
rect 20076 39618 20132 39788
rect 20076 39566 20078 39618
rect 20130 39566 20132 39618
rect 20076 39554 20132 39566
rect 20524 39620 20580 39630
rect 19404 38882 19460 38892
rect 19628 39506 19684 39518
rect 19628 39454 19630 39506
rect 19682 39454 19684 39506
rect 19180 38782 19182 38834
rect 19234 38782 19236 38834
rect 19180 38668 19236 38782
rect 19180 38612 19572 38668
rect 19404 38276 19460 38286
rect 19068 38052 19124 38062
rect 19068 37958 19124 37996
rect 19292 37826 19348 37838
rect 19292 37774 19294 37826
rect 19346 37774 19348 37826
rect 19180 37156 19236 37166
rect 18956 37154 19236 37156
rect 18956 37102 19182 37154
rect 19234 37102 19236 37154
rect 18956 37100 19236 37102
rect 19180 36932 19236 37100
rect 19180 36866 19236 36876
rect 18396 36540 18564 36596
rect 18844 36540 19124 36596
rect 18284 36484 18340 36494
rect 18284 36390 18340 36428
rect 18396 36372 18452 36382
rect 18396 36148 18452 36316
rect 18172 36092 18452 36148
rect 18396 35812 18452 36092
rect 18396 35746 18452 35756
rect 18508 36372 18564 36540
rect 18956 36372 19012 36382
rect 18508 36370 19012 36372
rect 18508 36318 18510 36370
rect 18562 36318 18958 36370
rect 19010 36318 19012 36370
rect 18508 36316 19012 36318
rect 18060 35186 18116 35196
rect 17836 35028 17892 35038
rect 17836 34934 17892 34972
rect 18508 34692 18564 36316
rect 18956 36306 19012 36316
rect 19068 35308 19124 36540
rect 19180 36372 19236 36382
rect 19180 36278 19236 36316
rect 19068 35252 19236 35308
rect 18508 34626 18564 34636
rect 19068 34692 19124 34702
rect 17388 34302 17390 34354
rect 17442 34302 17444 34354
rect 17388 34290 17444 34302
rect 18956 34356 19012 34366
rect 18620 34244 18676 34254
rect 17500 34018 17556 34030
rect 17500 33966 17502 34018
rect 17554 33966 17556 34018
rect 17164 33852 17444 33908
rect 16380 33460 16436 33470
rect 16380 33458 16772 33460
rect 16380 33406 16382 33458
rect 16434 33406 16772 33458
rect 16380 33404 16772 33406
rect 16380 33394 16436 33404
rect 16492 32788 16548 32798
rect 16044 32786 16548 32788
rect 16044 32734 16494 32786
rect 16546 32734 16548 32786
rect 16044 32732 16548 32734
rect 16044 32674 16100 32732
rect 16492 32722 16548 32732
rect 16044 32622 16046 32674
rect 16098 32622 16100 32674
rect 16044 32610 16100 32622
rect 16716 32676 16772 33404
rect 16828 33346 16884 33358
rect 16828 33294 16830 33346
rect 16882 33294 16884 33346
rect 16828 32788 16884 33294
rect 16828 32722 16884 32732
rect 16268 32562 16324 32574
rect 16268 32510 16270 32562
rect 16322 32510 16324 32562
rect 16268 32452 16324 32510
rect 16268 32386 16324 32396
rect 16380 32562 16436 32574
rect 16380 32510 16382 32562
rect 16434 32510 16436 32562
rect 16380 32116 16436 32510
rect 16604 32564 16660 32574
rect 16604 32470 16660 32508
rect 16716 32562 16772 32620
rect 16716 32510 16718 32562
rect 16770 32510 16772 32562
rect 16716 32498 16772 32510
rect 16380 32050 16436 32060
rect 16940 32116 16996 33516
rect 16940 32050 16996 32060
rect 17052 33684 17108 33694
rect 16268 32004 16324 32014
rect 16268 31890 16324 31948
rect 16268 31838 16270 31890
rect 16322 31838 16324 31890
rect 16268 31826 16324 31838
rect 16828 32002 16884 32014
rect 16828 31950 16830 32002
rect 16882 31950 16884 32002
rect 16828 31890 16884 31950
rect 16828 31838 16830 31890
rect 16882 31838 16884 31890
rect 16828 31826 16884 31838
rect 16828 30884 16884 30894
rect 17052 30884 17108 33628
rect 17388 32900 17444 33852
rect 17500 33684 17556 33966
rect 18060 34020 18116 34030
rect 18620 34020 18676 34188
rect 18956 34242 19012 34300
rect 19068 34354 19124 34636
rect 19068 34302 19070 34354
rect 19122 34302 19124 34354
rect 19068 34290 19124 34302
rect 18956 34190 18958 34242
rect 19010 34190 19012 34242
rect 18956 34178 19012 34190
rect 18060 34018 18340 34020
rect 18060 33966 18062 34018
rect 18114 33966 18340 34018
rect 18060 33964 18340 33966
rect 18060 33954 18116 33964
rect 17500 33618 17556 33628
rect 17948 33906 18004 33918
rect 17948 33854 17950 33906
rect 18002 33854 18004 33906
rect 17500 33460 17556 33470
rect 17500 33366 17556 33404
rect 17948 33460 18004 33854
rect 17948 33394 18004 33404
rect 18172 33684 18228 33694
rect 17276 32844 17444 32900
rect 17500 33124 17556 33134
rect 17276 32116 17332 32844
rect 17500 32786 17556 33068
rect 17500 32734 17502 32786
rect 17554 32734 17556 32786
rect 17500 32722 17556 32734
rect 17388 32676 17444 32686
rect 17388 32582 17444 32620
rect 17948 32562 18004 32574
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17948 32452 18004 32510
rect 18172 32564 18228 33628
rect 18284 32786 18340 33964
rect 18284 32734 18286 32786
rect 18338 32734 18340 32786
rect 18284 32722 18340 32734
rect 18508 34018 18676 34020
rect 18508 33966 18622 34018
rect 18674 33966 18676 34018
rect 18508 33964 18676 33966
rect 18396 32564 18452 32574
rect 18172 32562 18340 32564
rect 18172 32510 18174 32562
rect 18226 32510 18340 32562
rect 18172 32508 18340 32510
rect 18172 32498 18228 32508
rect 17276 32060 17444 32116
rect 17276 31780 17332 31790
rect 16828 30882 17220 30884
rect 16828 30830 16830 30882
rect 16882 30830 17220 30882
rect 16828 30828 17220 30830
rect 16828 30818 16884 30828
rect 16380 30212 16436 30222
rect 16380 29764 16436 30156
rect 17164 29876 17220 30828
rect 17276 30210 17332 31724
rect 17388 30882 17444 32060
rect 17836 31556 17892 31566
rect 17836 31462 17892 31500
rect 17388 30830 17390 30882
rect 17442 30830 17444 30882
rect 17388 30548 17444 30830
rect 17388 30482 17444 30492
rect 17276 30158 17278 30210
rect 17330 30158 17332 30210
rect 17276 30146 17332 30158
rect 17612 30212 17668 30222
rect 17164 29820 17444 29876
rect 16380 29650 16436 29708
rect 16380 29598 16382 29650
rect 16434 29598 16436 29650
rect 16380 29586 16436 29598
rect 17388 29538 17444 29820
rect 17612 29650 17668 30156
rect 17948 29988 18004 32396
rect 17836 29764 17892 29774
rect 17612 29598 17614 29650
rect 17666 29598 17668 29650
rect 17612 29586 17668 29598
rect 17724 29652 17780 29662
rect 17724 29558 17780 29596
rect 17836 29650 17892 29708
rect 17836 29598 17838 29650
rect 17890 29598 17892 29650
rect 17836 29586 17892 29598
rect 17948 29650 18004 29932
rect 17948 29598 17950 29650
rect 18002 29598 18004 29650
rect 17948 29586 18004 29598
rect 18060 32116 18116 32126
rect 17388 29486 17390 29538
rect 17442 29486 17444 29538
rect 17388 29474 17444 29486
rect 16940 29314 16996 29326
rect 16940 29262 16942 29314
rect 16994 29262 16996 29314
rect 16940 28644 16996 29262
rect 16940 28578 16996 28588
rect 17164 29316 17220 29326
rect 16380 28530 16436 28542
rect 16380 28478 16382 28530
rect 16434 28478 16436 28530
rect 15932 27346 15988 27356
rect 16268 27636 16324 27646
rect 16268 27186 16324 27580
rect 16268 27134 16270 27186
rect 16322 27134 16324 27186
rect 16268 27122 16324 27134
rect 15484 27022 15486 27074
rect 15538 27022 15540 27074
rect 15484 27010 15540 27022
rect 15372 26852 15540 26908
rect 15036 24670 15038 24722
rect 15090 24670 15092 24722
rect 15036 24658 15092 24670
rect 13916 24610 13972 24622
rect 13916 24558 13918 24610
rect 13970 24558 13972 24610
rect 13916 24276 13972 24558
rect 14700 24612 14756 24622
rect 14700 24518 14756 24556
rect 13692 24220 13972 24276
rect 14812 24276 14868 24286
rect 12908 23846 12964 23884
rect 13244 23940 13300 23950
rect 13020 23380 13076 23390
rect 13020 23154 13076 23324
rect 13020 23102 13022 23154
rect 13074 23102 13076 23154
rect 13020 23090 13076 23102
rect 13244 23154 13300 23884
rect 13244 23102 13246 23154
rect 13298 23102 13300 23154
rect 13244 23090 13300 23102
rect 13580 23716 13636 23726
rect 13580 23378 13636 23660
rect 13580 23326 13582 23378
rect 13634 23326 13636 23378
rect 12908 22484 12964 22494
rect 12908 22390 12964 22428
rect 12796 22082 12852 22092
rect 13244 21812 13300 21822
rect 13580 21812 13636 23326
rect 13692 23380 13748 24220
rect 13916 24052 13972 24062
rect 14700 24052 14756 24062
rect 13916 24050 14756 24052
rect 13916 23998 13918 24050
rect 13970 23998 14702 24050
rect 14754 23998 14756 24050
rect 13916 23996 14756 23998
rect 13916 23986 13972 23996
rect 14700 23986 14756 23996
rect 14812 24050 14868 24220
rect 14812 23998 14814 24050
rect 14866 23998 14868 24050
rect 14812 23986 14868 23998
rect 13804 23940 13860 23950
rect 13804 23846 13860 23884
rect 14028 23714 14084 23726
rect 14028 23662 14030 23714
rect 14082 23662 14084 23714
rect 14028 23380 14084 23662
rect 14252 23714 14308 23726
rect 14252 23662 14254 23714
rect 14306 23662 14308 23714
rect 13748 23324 14084 23380
rect 14140 23604 14196 23614
rect 13692 23286 13748 23324
rect 13692 22484 13748 22494
rect 13692 22370 13748 22428
rect 13692 22318 13694 22370
rect 13746 22318 13748 22370
rect 13692 21924 13748 22318
rect 13916 22260 13972 23324
rect 14028 23156 14084 23166
rect 14140 23156 14196 23548
rect 14028 23154 14196 23156
rect 14028 23102 14030 23154
rect 14082 23102 14196 23154
rect 14028 23100 14196 23102
rect 14028 23090 14084 23100
rect 14028 22260 14084 22270
rect 13916 22204 14028 22260
rect 14028 22194 14084 22204
rect 13804 22148 13860 22158
rect 13804 22054 13860 22092
rect 14140 21924 14196 21934
rect 13692 21868 14140 21924
rect 13580 21756 13972 21812
rect 13244 21474 13300 21756
rect 13244 21422 13246 21474
rect 13298 21422 13300 21474
rect 13244 21410 13300 21422
rect 13356 21698 13412 21710
rect 13356 21646 13358 21698
rect 13410 21646 13412 21698
rect 11900 21308 13188 21364
rect 12908 21028 12964 21038
rect 12908 20914 12964 20972
rect 12908 20862 12910 20914
rect 12962 20862 12964 20914
rect 12684 20804 12740 20814
rect 12684 20710 12740 20748
rect 11788 20580 11844 20590
rect 12348 20580 12404 20590
rect 11788 20486 11844 20524
rect 12012 20578 12404 20580
rect 12012 20526 12350 20578
rect 12402 20526 12404 20578
rect 12012 20524 12404 20526
rect 12012 19348 12068 20524
rect 12348 20514 12404 20524
rect 12012 18674 12068 19292
rect 12908 19346 12964 20862
rect 12908 19294 12910 19346
rect 12962 19294 12964 19346
rect 12908 19282 12964 19294
rect 13020 20018 13076 20030
rect 13020 19966 13022 20018
rect 13074 19966 13076 20018
rect 13020 19908 13076 19966
rect 12012 18622 12014 18674
rect 12066 18622 12068 18674
rect 12012 18610 12068 18622
rect 12236 19236 12292 19246
rect 11900 18452 11956 18462
rect 11900 18338 11956 18396
rect 12236 18450 12292 19180
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 12236 18386 12292 18398
rect 12908 19124 12964 19134
rect 11900 18286 11902 18338
rect 11954 18286 11956 18338
rect 11900 18274 11956 18286
rect 12572 18338 12628 18350
rect 12572 18286 12574 18338
rect 12626 18286 12628 18338
rect 12572 17668 12628 18286
rect 12908 17778 12964 19068
rect 13020 18564 13076 19852
rect 13020 18498 13076 18508
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17714 12964 17726
rect 12572 17602 12628 17612
rect 12796 16996 12852 17006
rect 12796 16902 12852 16940
rect 13020 16882 13076 16894
rect 13020 16830 13022 16882
rect 13074 16830 13076 16882
rect 12460 16770 12516 16782
rect 12460 16718 12462 16770
rect 12514 16718 12516 16770
rect 12460 16548 12516 16718
rect 12908 16772 12964 16782
rect 12908 16678 12964 16716
rect 13020 16548 13076 16830
rect 12460 16492 13076 16548
rect 11788 16212 11844 16222
rect 12460 16212 12516 16492
rect 11788 16210 12516 16212
rect 11788 16158 11790 16210
rect 11842 16158 12516 16210
rect 11788 16156 12516 16158
rect 11788 16146 11844 16156
rect 11900 15202 11956 15214
rect 11900 15150 11902 15202
rect 11954 15150 11956 15202
rect 11900 14644 11956 15150
rect 13132 14868 13188 21308
rect 13356 20804 13412 21646
rect 13916 21698 13972 21756
rect 14140 21810 14196 21868
rect 14140 21758 14142 21810
rect 14194 21758 14196 21810
rect 14140 21746 14196 21758
rect 13916 21646 13918 21698
rect 13970 21646 13972 21698
rect 13916 21634 13972 21646
rect 14252 21588 14308 23662
rect 14924 23716 14980 23726
rect 14980 23660 15092 23716
rect 14924 23622 14980 23660
rect 14700 23268 14756 23278
rect 14700 23174 14756 23212
rect 14812 22260 14868 22270
rect 14812 22258 14980 22260
rect 14812 22206 14814 22258
rect 14866 22206 14980 22258
rect 14812 22204 14980 22206
rect 14812 22194 14868 22204
rect 14812 21924 14868 21934
rect 14476 21588 14532 21598
rect 14252 21586 14532 21588
rect 14252 21534 14478 21586
rect 14530 21534 14532 21586
rect 14252 21532 14532 21534
rect 14028 21474 14084 21486
rect 14028 21422 14030 21474
rect 14082 21422 14084 21474
rect 13580 21364 13636 21374
rect 14028 21364 14084 21422
rect 13580 21362 14084 21364
rect 13580 21310 13582 21362
rect 13634 21310 14084 21362
rect 13580 21308 14084 21310
rect 13580 21298 13636 21308
rect 14252 21028 14308 21038
rect 13356 20738 13412 20748
rect 14028 20804 14084 20814
rect 14028 20710 14084 20748
rect 14252 20802 14308 20972
rect 14252 20750 14254 20802
rect 14306 20750 14308 20802
rect 14252 20738 14308 20750
rect 14140 20578 14196 20590
rect 14476 20580 14532 21532
rect 14812 21586 14868 21868
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14812 21522 14868 21534
rect 14140 20526 14142 20578
rect 14194 20526 14196 20578
rect 13580 19460 13636 19470
rect 13580 19234 13636 19404
rect 13804 19348 13860 19358
rect 13804 19254 13860 19292
rect 13580 19182 13582 19234
rect 13634 19182 13636 19234
rect 13580 19170 13636 19182
rect 14140 19236 14196 20526
rect 14140 19170 14196 19180
rect 14364 20578 14532 20580
rect 14364 20526 14478 20578
rect 14530 20526 14532 20578
rect 14364 20524 14532 20526
rect 14364 19012 14420 20524
rect 14476 20514 14532 20524
rect 14924 19796 14980 22204
rect 15036 21586 15092 23660
rect 15036 21534 15038 21586
rect 15090 21534 15092 21586
rect 15036 21522 15092 21534
rect 15372 21362 15428 21374
rect 15372 21310 15374 21362
rect 15426 21310 15428 21362
rect 15260 20802 15316 20814
rect 15260 20750 15262 20802
rect 15314 20750 15316 20802
rect 15260 20132 15316 20750
rect 15372 20804 15428 21310
rect 15372 20738 15428 20748
rect 15316 20076 15428 20132
rect 15260 20038 15316 20076
rect 14476 19740 14980 19796
rect 14476 19234 14532 19740
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19124 14532 19182
rect 14476 19058 14532 19068
rect 15036 19234 15092 19246
rect 15036 19182 15038 19234
rect 15090 19182 15092 19234
rect 14028 18956 14420 19012
rect 13916 17668 13972 17678
rect 14028 17668 14084 18956
rect 13916 17666 14084 17668
rect 13916 17614 13918 17666
rect 13970 17614 14084 17666
rect 13916 17612 14084 17614
rect 14140 18452 14196 18462
rect 13244 17108 13300 17118
rect 13244 17014 13300 17052
rect 13916 15540 13972 17612
rect 14028 16884 14084 16894
rect 14140 16884 14196 18396
rect 14700 18340 14756 18350
rect 14588 18338 14756 18340
rect 14588 18286 14702 18338
rect 14754 18286 14756 18338
rect 14588 18284 14756 18286
rect 14476 18116 14532 18126
rect 14252 17668 14308 17678
rect 14252 17574 14308 17612
rect 14476 17666 14532 18060
rect 14476 17614 14478 17666
rect 14530 17614 14532 17666
rect 14476 17602 14532 17614
rect 14028 16882 14196 16884
rect 14028 16830 14030 16882
rect 14082 16830 14196 16882
rect 14028 16828 14196 16830
rect 14364 17442 14420 17454
rect 14364 17390 14366 17442
rect 14418 17390 14420 17442
rect 14028 16818 14084 16828
rect 14364 16324 14420 17390
rect 14588 16772 14644 18284
rect 14700 18274 14756 18284
rect 15036 17668 15092 19182
rect 15260 19234 15316 19246
rect 15260 19182 15262 19234
rect 15314 19182 15316 19234
rect 15260 18116 15316 19182
rect 15372 18452 15428 20076
rect 15484 19124 15540 26852
rect 16380 25620 16436 28478
rect 16940 28420 16996 28430
rect 16828 27746 16884 27758
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 16828 27524 16884 27694
rect 16828 27458 16884 27468
rect 16828 26292 16884 26302
rect 16828 26178 16884 26236
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 26114 16884 26126
rect 16380 24724 16436 25564
rect 16492 25396 16548 25406
rect 16492 25282 16548 25340
rect 16492 25230 16494 25282
rect 16546 25230 16548 25282
rect 16492 25218 16548 25230
rect 16828 25284 16884 25294
rect 16828 24834 16884 25228
rect 16828 24782 16830 24834
rect 16882 24782 16884 24834
rect 16828 24770 16884 24782
rect 16380 24630 16436 24668
rect 15708 24612 15764 24622
rect 15708 23938 15764 24556
rect 16716 24500 16772 24510
rect 16380 24498 16772 24500
rect 16380 24446 16718 24498
rect 16770 24446 16772 24498
rect 16380 24444 16772 24446
rect 16380 24050 16436 24444
rect 16716 24434 16772 24444
rect 16380 23998 16382 24050
rect 16434 23998 16436 24050
rect 16380 23986 16436 23998
rect 15708 23886 15710 23938
rect 15762 23886 15764 23938
rect 15708 23604 15764 23886
rect 15708 23538 15764 23548
rect 16156 23828 16212 23838
rect 15708 22370 15764 22382
rect 15708 22318 15710 22370
rect 15762 22318 15764 22370
rect 15708 21028 15764 22318
rect 15932 21812 15988 21822
rect 15932 21718 15988 21756
rect 15708 20962 15764 20972
rect 16156 20804 16212 23772
rect 16828 23156 16884 23166
rect 16380 23044 16436 23054
rect 16380 22708 16436 22988
rect 16828 23042 16884 23100
rect 16828 22990 16830 23042
rect 16882 22990 16884 23042
rect 16828 22978 16884 22990
rect 16268 22260 16324 22270
rect 16268 22166 16324 22204
rect 16380 21474 16436 22652
rect 16380 21422 16382 21474
rect 16434 21422 16436 21474
rect 16380 21410 16436 21422
rect 16716 21586 16772 21598
rect 16716 21534 16718 21586
rect 16770 21534 16772 21586
rect 16716 21252 16772 21534
rect 16716 21186 16772 21196
rect 16156 20748 16324 20804
rect 16044 20692 16100 20702
rect 16044 20690 16212 20692
rect 16044 20638 16046 20690
rect 16098 20638 16212 20690
rect 16044 20636 16212 20638
rect 16044 20626 16100 20636
rect 16156 19458 16212 20636
rect 16156 19406 16158 19458
rect 16210 19406 16212 19458
rect 16156 19394 16212 19406
rect 16268 19458 16324 20748
rect 16268 19406 16270 19458
rect 16322 19406 16324 19458
rect 15484 19058 15540 19068
rect 15372 18358 15428 18396
rect 15596 19010 15652 19022
rect 15596 18958 15598 19010
rect 15650 18958 15652 19010
rect 15260 18050 15316 18060
rect 15036 17602 15092 17612
rect 15596 16996 15652 18958
rect 16268 18564 16324 19406
rect 16268 18498 16324 18508
rect 16492 20580 16548 20590
rect 16492 19458 16548 20524
rect 16716 20356 16772 20366
rect 16492 19406 16494 19458
rect 16546 19406 16548 19458
rect 16492 18452 16548 19406
rect 16604 20300 16716 20356
rect 16604 19012 16660 20300
rect 16716 20290 16772 20300
rect 16716 19908 16772 19918
rect 16716 19234 16772 19852
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 16716 19170 16772 19182
rect 16604 18956 16772 19012
rect 16604 18452 16660 18462
rect 16380 18450 16660 18452
rect 16380 18398 16606 18450
rect 16658 18398 16660 18450
rect 16380 18396 16660 18398
rect 15932 18340 15988 18350
rect 15932 17780 15988 18284
rect 16268 18228 16324 18238
rect 15932 17714 15988 17724
rect 16156 18226 16324 18228
rect 16156 18174 16270 18226
rect 16322 18174 16324 18226
rect 16156 18172 16324 18174
rect 16044 17666 16100 17678
rect 16044 17614 16046 17666
rect 16098 17614 16100 17666
rect 16044 17108 16100 17614
rect 16044 17042 16100 17052
rect 15652 16940 15876 16996
rect 15596 16930 15652 16940
rect 14588 16706 14644 16716
rect 14700 16772 14756 16782
rect 14700 16770 14980 16772
rect 14700 16718 14702 16770
rect 14754 16718 14980 16770
rect 14700 16716 14980 16718
rect 14700 16706 14756 16716
rect 14364 16258 14420 16268
rect 14924 16322 14980 16716
rect 14924 16270 14926 16322
rect 14978 16270 14980 16322
rect 14924 16258 14980 16270
rect 15036 16660 15092 16670
rect 15036 15986 15092 16604
rect 15596 16324 15652 16334
rect 15596 16230 15652 16268
rect 15036 15934 15038 15986
rect 15090 15934 15092 15986
rect 15036 15764 15092 15934
rect 15260 15988 15316 15998
rect 15260 15894 15316 15932
rect 15820 15874 15876 16940
rect 15932 16772 15988 16782
rect 15932 16322 15988 16716
rect 16156 16660 16212 18172
rect 16268 18162 16324 18172
rect 16380 17444 16436 18396
rect 16604 18386 16660 18396
rect 16156 16594 16212 16604
rect 16268 17388 16436 17444
rect 15932 16270 15934 16322
rect 15986 16270 15988 16322
rect 15932 16258 15988 16270
rect 15820 15822 15822 15874
rect 15874 15822 15876 15874
rect 15820 15810 15876 15822
rect 16268 15874 16324 17388
rect 16492 16772 16548 16782
rect 16492 16098 16548 16716
rect 16492 16046 16494 16098
rect 16546 16046 16548 16098
rect 16492 16034 16548 16046
rect 16380 15988 16436 15998
rect 16380 15894 16436 15932
rect 16268 15822 16270 15874
rect 16322 15822 16324 15874
rect 16268 15810 16324 15822
rect 15036 15698 15092 15708
rect 14364 15540 14420 15550
rect 13916 15538 14420 15540
rect 13916 15486 14366 15538
rect 14418 15486 14420 15538
rect 13916 15484 14420 15486
rect 14364 15474 14420 15484
rect 14700 15540 14756 15550
rect 15036 15540 15092 15550
rect 14700 15538 15092 15540
rect 14700 15486 14702 15538
rect 14754 15486 15038 15538
rect 15090 15486 15092 15538
rect 14700 15484 15092 15486
rect 14028 15202 14084 15214
rect 14028 15150 14030 15202
rect 14082 15150 14084 15202
rect 14028 15148 14084 15150
rect 14700 15148 14756 15484
rect 15036 15474 15092 15484
rect 12796 14812 13132 14868
rect 12012 14644 12068 14654
rect 11900 14642 12068 14644
rect 11900 14590 12014 14642
rect 12066 14590 12068 14642
rect 11900 14588 12068 14590
rect 12012 14578 12068 14588
rect 11788 14530 11844 14542
rect 12236 14532 12292 14542
rect 11788 14478 11790 14530
rect 11842 14478 11844 14530
rect 11788 14420 11844 14478
rect 11788 14354 11844 14364
rect 12124 14476 12236 14532
rect 12124 13972 12180 14476
rect 12236 14438 12292 14476
rect 12460 14420 12516 14430
rect 12460 14326 12516 14364
rect 12124 13858 12180 13916
rect 12124 13806 12126 13858
rect 12178 13806 12180 13858
rect 12124 13794 12180 13806
rect 12572 14308 12628 14318
rect 12012 13746 12068 13758
rect 12012 13694 12014 13746
rect 12066 13694 12068 13746
rect 12012 13636 12068 13694
rect 12012 13570 12068 13580
rect 12236 13746 12292 13758
rect 12236 13694 12238 13746
rect 12290 13694 12292 13746
rect 12236 12404 12292 13694
rect 12572 13746 12628 14252
rect 12572 13694 12574 13746
rect 12626 13694 12628 13746
rect 12572 13682 12628 13694
rect 12236 11506 12292 12348
rect 12684 12180 12740 12190
rect 12236 11454 12238 11506
rect 12290 11454 12292 11506
rect 12236 11442 12292 11454
rect 12348 12178 12740 12180
rect 12348 12126 12686 12178
rect 12738 12126 12740 12178
rect 12348 12124 12740 12126
rect 11788 10612 11844 10622
rect 11788 9828 11844 10556
rect 11900 10612 11956 10622
rect 12348 10612 12404 12124
rect 12684 12114 12740 12124
rect 12572 11506 12628 11518
rect 12572 11454 12574 11506
rect 12626 11454 12628 11506
rect 12572 10722 12628 11454
rect 12572 10670 12574 10722
rect 12626 10670 12628 10722
rect 12572 10658 12628 10670
rect 12684 11170 12740 11182
rect 12684 11118 12686 11170
rect 12738 11118 12740 11170
rect 11900 10610 12404 10612
rect 11900 10558 11902 10610
rect 11954 10558 12404 10610
rect 11900 10556 12404 10558
rect 11900 10546 11956 10556
rect 12348 10500 12404 10556
rect 12684 10612 12740 11118
rect 12684 10546 12740 10556
rect 12348 10434 12404 10444
rect 12012 9940 12068 9950
rect 12012 9846 12068 9884
rect 11900 9828 11956 9838
rect 11788 9772 11900 9828
rect 11900 9734 11956 9772
rect 12236 9828 12292 9838
rect 12124 9604 12180 9614
rect 12012 9602 12180 9604
rect 12012 9550 12126 9602
rect 12178 9550 12180 9602
rect 12012 9548 12180 9550
rect 11788 9268 11844 9278
rect 12012 9268 12068 9548
rect 12124 9538 12180 9548
rect 11844 9212 12068 9268
rect 11788 9202 11844 9212
rect 11340 9062 11396 9100
rect 11564 9100 11732 9156
rect 11900 9154 11956 9212
rect 11900 9102 11902 9154
rect 11954 9102 11956 9154
rect 9884 8708 9940 8876
rect 9436 8258 9492 8540
rect 9884 8428 9940 8652
rect 10668 8930 10724 8942
rect 10668 8878 10670 8930
rect 10722 8878 10724 8930
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 9436 8194 9492 8206
rect 9660 8372 9940 8428
rect 10108 8484 10164 8494
rect 9660 8258 9716 8372
rect 9660 8206 9662 8258
rect 9714 8206 9716 8258
rect 9660 8194 9716 8206
rect 9212 7532 9492 7588
rect 9436 7476 9492 7532
rect 9548 7476 9604 7486
rect 9100 7420 9268 7476
rect 9436 7474 9604 7476
rect 9436 7422 9550 7474
rect 9602 7422 9604 7474
rect 9436 7420 9604 7422
rect 8988 7362 9156 7364
rect 8988 7310 8990 7362
rect 9042 7310 9156 7362
rect 8988 7308 9156 7310
rect 8988 7298 9044 7308
rect 8876 6748 9044 6804
rect 8204 6598 8260 6636
rect 8316 6636 8596 6692
rect 8204 6468 8260 6478
rect 8316 6468 8372 6636
rect 8876 6580 8932 6590
rect 8260 6412 8372 6468
rect 8540 6578 8932 6580
rect 8540 6526 8878 6578
rect 8930 6526 8932 6578
rect 8540 6524 8932 6526
rect 8204 6402 8260 6412
rect 7868 5954 7924 5964
rect 8316 6244 8372 6254
rect 7532 5854 7534 5906
rect 7586 5854 7588 5906
rect 7532 5842 7588 5854
rect 7980 5908 8036 5918
rect 8204 5908 8260 5918
rect 7980 5906 8260 5908
rect 7980 5854 7982 5906
rect 8034 5854 8206 5906
rect 8258 5854 8260 5906
rect 7980 5852 8260 5854
rect 7980 5842 8036 5852
rect 8204 5842 8260 5852
rect 7308 5170 7364 5180
rect 8204 5236 8260 5246
rect 8316 5236 8372 6188
rect 8540 6130 8596 6524
rect 8876 6514 8932 6524
rect 8540 6078 8542 6130
rect 8594 6078 8596 6130
rect 8540 6066 8596 6078
rect 8764 6356 8820 6366
rect 8204 5234 8372 5236
rect 8204 5182 8206 5234
rect 8258 5182 8372 5234
rect 8204 5180 8372 5182
rect 8540 5236 8596 5246
rect 8204 5170 8260 5180
rect 8540 5142 8596 5180
rect 6300 5070 6302 5122
rect 6354 5070 6356 5122
rect 6300 5058 6356 5070
rect 4956 4958 4958 5010
rect 5010 4958 5012 5010
rect 4956 4946 5012 4958
rect 6972 5012 7028 5022
rect 7756 5012 7812 5022
rect 6972 5010 7476 5012
rect 6972 4958 6974 5010
rect 7026 4958 7476 5010
rect 6972 4956 7476 4958
rect 6972 4946 7028 4956
rect 7420 4450 7476 4956
rect 7420 4398 7422 4450
rect 7474 4398 7476 4450
rect 7420 4386 7476 4398
rect 7084 4340 7140 4350
rect 7084 4246 7140 4284
rect 7756 4338 7812 4956
rect 8652 4564 8708 4574
rect 8652 4470 8708 4508
rect 7756 4286 7758 4338
rect 7810 4286 7812 4338
rect 7756 4274 7812 4286
rect 8428 4338 8484 4350
rect 8428 4286 8430 4338
rect 8482 4286 8484 4338
rect 4172 4174 4174 4226
rect 4226 4174 4228 4226
rect 4172 4162 4228 4174
rect 6300 4228 6356 4238
rect 6300 4134 6356 4172
rect 7532 4228 7588 4238
rect 7532 4134 7588 4172
rect 8428 4116 8484 4286
rect 8764 4340 8820 6300
rect 8988 5124 9044 6748
rect 9100 6244 9156 7308
rect 9100 6178 9156 6188
rect 9100 6020 9156 6030
rect 9100 5926 9156 5964
rect 9100 5684 9156 5694
rect 9212 5684 9268 7420
rect 9156 5628 9268 5684
rect 9436 6580 9492 6590
rect 9100 5618 9156 5628
rect 8764 4274 8820 4284
rect 8876 5068 9044 5124
rect 8876 4116 8932 5068
rect 9436 5012 9492 6524
rect 9548 6356 9604 7420
rect 9548 6290 9604 6300
rect 10108 5906 10164 8428
rect 10668 8372 10724 8878
rect 11228 8818 11284 8830
rect 11228 8766 11230 8818
rect 11282 8766 11284 8818
rect 11228 8428 11284 8766
rect 10220 8316 10668 8372
rect 10220 8146 10276 8316
rect 10668 8306 10724 8316
rect 11116 8372 11284 8428
rect 11564 8428 11620 9100
rect 11900 9090 11956 9102
rect 12124 9154 12180 9166
rect 12124 9102 12126 9154
rect 12178 9102 12180 9154
rect 11788 9042 11844 9054
rect 11788 8990 11790 9042
rect 11842 8990 11844 9042
rect 11788 8932 11844 8990
rect 11788 8866 11844 8876
rect 12124 8428 12180 9102
rect 12236 9042 12292 9772
rect 12348 9716 12404 9726
rect 12348 9622 12404 9660
rect 12236 8990 12238 9042
rect 12290 8990 12292 9042
rect 12236 8978 12292 8990
rect 12684 9044 12740 9054
rect 12684 8950 12740 8988
rect 11564 8372 11732 8428
rect 11116 8370 11172 8372
rect 11116 8318 11118 8370
rect 11170 8318 11172 8370
rect 11116 8306 11172 8318
rect 11452 8260 11508 8270
rect 11452 8166 11508 8204
rect 10220 8094 10222 8146
rect 10274 8094 10276 8146
rect 10220 8082 10276 8094
rect 10444 8148 10500 8158
rect 10780 8148 10836 8158
rect 10444 8146 10836 8148
rect 10444 8094 10446 8146
rect 10498 8094 10782 8146
rect 10834 8094 10836 8146
rect 10444 8092 10836 8094
rect 10444 8082 10500 8092
rect 10780 8082 10836 8092
rect 10332 8034 10388 8046
rect 10332 7982 10334 8034
rect 10386 7982 10388 8034
rect 10332 7586 10388 7982
rect 10332 7534 10334 7586
rect 10386 7534 10388 7586
rect 10332 7522 10388 7534
rect 11004 7476 11060 7486
rect 10108 5854 10110 5906
rect 10162 5854 10164 5906
rect 10108 5842 10164 5854
rect 10780 6804 10836 6814
rect 9660 5796 9716 5806
rect 9660 5346 9716 5740
rect 9660 5294 9662 5346
rect 9714 5294 9716 5346
rect 9660 5282 9716 5294
rect 9548 5236 9604 5246
rect 9548 5142 9604 5180
rect 10780 5234 10836 6748
rect 11004 6802 11060 7420
rect 11676 7364 11732 8316
rect 12124 8372 12516 8428
rect 12124 8260 12180 8372
rect 12124 8194 12180 8204
rect 11676 7298 11732 7308
rect 12460 7362 12516 8372
rect 12460 7310 12462 7362
rect 12514 7310 12516 7362
rect 12460 7298 12516 7310
rect 12684 8036 12740 8046
rect 12236 6916 12292 6926
rect 12236 6822 12292 6860
rect 11004 6750 11006 6802
rect 11058 6750 11060 6802
rect 11004 6738 11060 6750
rect 12572 6804 12628 6814
rect 12572 6710 12628 6748
rect 12012 6692 12068 6702
rect 12012 6578 12068 6636
rect 12012 6526 12014 6578
rect 12066 6526 12068 6578
rect 12012 6514 12068 6526
rect 12684 6578 12740 7980
rect 12684 6526 12686 6578
rect 12738 6526 12740 6578
rect 12684 6514 12740 6526
rect 11004 6468 11060 6478
rect 10780 5182 10782 5234
rect 10834 5182 10836 5234
rect 10780 5170 10836 5182
rect 10892 6412 11004 6468
rect 9100 5010 9492 5012
rect 9100 4958 9438 5010
rect 9490 4958 9492 5010
rect 9100 4956 9492 4958
rect 8988 4900 9044 4910
rect 8988 4806 9044 4844
rect 8428 4060 8932 4116
rect 9100 4004 9156 4956
rect 9436 4946 9492 4956
rect 10108 5124 10164 5134
rect 9660 4452 9716 4462
rect 9660 4358 9716 4396
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 8540 3948 9156 4004
rect 9772 4340 9828 4350
rect 10108 4340 10164 5068
rect 9828 4338 10164 4340
rect 9828 4286 10110 4338
rect 10162 4286 10164 4338
rect 9828 4284 10164 4286
rect 8540 3442 8596 3948
rect 8764 3780 8820 3790
rect 8764 3686 8820 3724
rect 9772 3554 9828 4284
rect 10108 4274 10164 4284
rect 10556 4900 10612 4910
rect 9772 3502 9774 3554
rect 9826 3502 9828 3554
rect 9772 3490 9828 3502
rect 8540 3390 8542 3442
rect 8594 3390 8596 3442
rect 8540 3378 8596 3390
rect 8652 3444 8708 3454
rect 8652 3350 8708 3388
rect 10444 3444 10500 3454
rect 10444 3350 10500 3388
rect 2940 3332 2996 3342
rect 4508 3332 4564 3342
rect 6076 3332 6132 3342
rect 7532 3332 7588 3342
rect 2716 3330 2996 3332
rect 2716 3278 2942 3330
rect 2994 3278 2996 3330
rect 2716 3276 2996 3278
rect 2716 800 2772 3276
rect 2940 3266 2996 3276
rect 4284 3330 4564 3332
rect 4284 3278 4510 3330
rect 4562 3278 4564 3330
rect 4284 3276 4564 3278
rect 4284 800 4340 3276
rect 4508 3266 4564 3276
rect 5852 3330 6132 3332
rect 5852 3278 6078 3330
rect 6130 3278 6132 3330
rect 5852 3276 6132 3278
rect 5852 800 5908 3276
rect 6076 3266 6132 3276
rect 7420 3330 7588 3332
rect 7420 3278 7534 3330
rect 7586 3278 7588 3330
rect 7420 3276 7588 3278
rect 7420 800 7476 3276
rect 7532 3266 7588 3276
rect 8092 3332 8148 3342
rect 8092 3330 8484 3332
rect 8092 3278 8094 3330
rect 8146 3278 8484 3330
rect 8092 3276 8484 3278
rect 8092 3266 8148 3276
rect 8428 980 8484 3276
rect 8428 924 9044 980
rect 8988 800 9044 924
rect 10556 800 10612 4844
rect 10780 4452 10836 4462
rect 10892 4452 10948 6412
rect 11004 6402 11060 6412
rect 11564 6466 11620 6478
rect 11564 6414 11566 6466
rect 11618 6414 11620 6466
rect 10780 4450 10948 4452
rect 10780 4398 10782 4450
rect 10834 4398 10948 4450
rect 10780 4396 10948 4398
rect 10780 4386 10836 4396
rect 11564 3444 11620 6414
rect 12124 6468 12180 6478
rect 12124 6374 12180 6412
rect 12796 6020 12852 14812
rect 13132 14802 13188 14812
rect 13692 15092 14084 15148
rect 14140 15092 14196 15102
rect 13020 14644 13076 14654
rect 13020 14550 13076 14588
rect 13692 14532 13748 15092
rect 13692 14438 13748 14476
rect 14140 14644 14196 15036
rect 14140 14530 14196 14588
rect 14140 14478 14142 14530
rect 14194 14478 14196 14530
rect 14140 14466 14196 14478
rect 14588 15092 14756 15148
rect 14924 15316 14980 15326
rect 13580 14420 13636 14430
rect 13580 14326 13636 14364
rect 13468 14308 13524 14318
rect 13468 13970 13524 14252
rect 13468 13918 13470 13970
rect 13522 13918 13524 13970
rect 13468 13906 13524 13918
rect 14028 14084 14084 14094
rect 13132 13860 13188 13870
rect 13132 13766 13188 13804
rect 13804 13858 13860 13870
rect 13804 13806 13806 13858
rect 13858 13806 13860 13858
rect 13804 13636 13860 13806
rect 14028 13746 14084 14028
rect 14588 14084 14644 15092
rect 14924 14530 14980 15260
rect 15260 15316 15316 15326
rect 15260 15222 15316 15260
rect 16268 15204 16324 15214
rect 16716 15148 16772 18956
rect 16828 18338 16884 18350
rect 16828 18286 16830 18338
rect 16882 18286 16884 18338
rect 16828 16772 16884 18286
rect 16828 16678 16884 16716
rect 16940 16098 16996 28364
rect 17164 22372 17220 29260
rect 17948 28756 18004 28766
rect 17836 27972 17892 27982
rect 17836 27878 17892 27916
rect 17948 27970 18004 28700
rect 17948 27918 17950 27970
rect 18002 27918 18004 27970
rect 17948 27906 18004 27918
rect 17500 27748 17556 27758
rect 17500 27654 17556 27692
rect 17388 27636 17444 27646
rect 17388 27542 17444 27580
rect 18060 26908 18116 32060
rect 18284 32002 18340 32508
rect 18396 32470 18452 32508
rect 18508 32340 18564 33964
rect 18620 33954 18676 33964
rect 18620 33460 18676 33470
rect 18620 32674 18676 33404
rect 18620 32622 18622 32674
rect 18674 32622 18676 32674
rect 18620 32610 18676 32622
rect 19068 32674 19124 32686
rect 19068 32622 19070 32674
rect 19122 32622 19124 32674
rect 19068 32564 19124 32622
rect 19068 32498 19124 32508
rect 18284 31950 18286 32002
rect 18338 31950 18340 32002
rect 18172 31554 18228 31566
rect 18172 31502 18174 31554
rect 18226 31502 18228 31554
rect 18172 31332 18228 31502
rect 18172 30324 18228 31276
rect 18172 30258 18228 30268
rect 18284 27188 18340 31950
rect 18396 32284 18564 32340
rect 18396 28420 18452 32284
rect 18508 31666 18564 31678
rect 18508 31614 18510 31666
rect 18562 31614 18564 31666
rect 18508 30772 18564 31614
rect 19180 31668 19236 35252
rect 19292 34354 19348 37774
rect 19404 36596 19460 38220
rect 19516 37492 19572 38612
rect 19628 38052 19684 39454
rect 20188 39396 20244 39406
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20076 38836 20132 38846
rect 20076 38162 20132 38780
rect 20188 38834 20244 39340
rect 20188 38782 20190 38834
rect 20242 38782 20244 38834
rect 20188 38770 20244 38782
rect 20300 39060 20356 39070
rect 20300 38668 20356 39004
rect 20076 38110 20078 38162
rect 20130 38110 20132 38162
rect 20076 38098 20132 38110
rect 20188 38612 20356 38668
rect 20412 38724 20468 38734
rect 19628 37986 19684 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19516 37436 19908 37492
rect 19404 36540 19684 36596
rect 19516 36372 19572 36382
rect 19404 36258 19460 36270
rect 19404 36206 19406 36258
rect 19458 36206 19460 36258
rect 19404 35700 19460 36206
rect 19404 35634 19460 35644
rect 19516 34468 19572 36316
rect 19516 34402 19572 34412
rect 19292 34302 19294 34354
rect 19346 34302 19348 34354
rect 19292 34290 19348 34302
rect 19404 33572 19460 33582
rect 19404 32786 19460 33516
rect 19628 33460 19684 36540
rect 19852 36594 19908 37436
rect 19852 36542 19854 36594
rect 19906 36542 19908 36594
rect 19852 36530 19908 36542
rect 20188 36594 20244 38612
rect 20300 38276 20356 38286
rect 20300 38050 20356 38220
rect 20300 37998 20302 38050
rect 20354 37998 20356 38050
rect 20300 37986 20356 37998
rect 20412 37938 20468 38668
rect 20412 37886 20414 37938
rect 20466 37886 20468 37938
rect 20412 37874 20468 37886
rect 20188 36542 20190 36594
rect 20242 36542 20244 36594
rect 20188 36530 20244 36542
rect 20300 37268 20356 37278
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 34804 20020 34814
rect 19964 34710 20020 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19964 34020 20020 34030
rect 19964 33926 20020 33964
rect 19628 33366 19684 33404
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19404 32734 19406 32786
rect 19458 32734 19460 32786
rect 19404 32722 19460 32734
rect 19740 32788 19796 32798
rect 19516 32564 19572 32574
rect 19740 32564 19796 32732
rect 20300 32676 20356 37212
rect 20412 36260 20468 36270
rect 20412 36166 20468 36204
rect 20412 35698 20468 35710
rect 20412 35646 20414 35698
rect 20466 35646 20468 35698
rect 20412 35252 20468 35646
rect 20412 34354 20468 35196
rect 20412 34302 20414 34354
rect 20466 34302 20468 34354
rect 20412 34290 20468 34302
rect 20524 35028 20580 39564
rect 20636 38722 20692 41022
rect 21420 41076 21476 41086
rect 20860 40964 20916 40974
rect 20860 40870 20916 40908
rect 21420 39842 21476 41020
rect 21420 39790 21422 39842
rect 21474 39790 21476 39842
rect 21420 39778 21476 39790
rect 21308 39508 21364 39518
rect 21308 39414 21364 39452
rect 21532 39060 21588 41244
rect 21644 40628 21700 40638
rect 21644 40514 21700 40572
rect 21644 40462 21646 40514
rect 21698 40462 21700 40514
rect 21644 40450 21700 40462
rect 21756 40404 21812 42814
rect 21868 42754 21924 42924
rect 21868 42702 21870 42754
rect 21922 42702 21924 42754
rect 21868 42690 21924 42702
rect 21980 42756 22036 42766
rect 21980 41858 22036 42700
rect 21980 41806 21982 41858
rect 22034 41806 22036 41858
rect 21868 40404 21924 40414
rect 21756 40402 21924 40404
rect 21756 40350 21870 40402
rect 21922 40350 21924 40402
rect 21756 40348 21924 40350
rect 21868 40338 21924 40348
rect 21868 39620 21924 39630
rect 21980 39620 22036 41806
rect 22876 42754 22932 42766
rect 22876 42702 22878 42754
rect 22930 42702 22932 42754
rect 22876 40964 22932 42702
rect 22876 40898 22932 40908
rect 22988 40852 23044 43652
rect 23212 43764 23268 43774
rect 23212 42756 23268 43708
rect 23324 43708 23380 44044
rect 23660 44098 23716 44110
rect 23660 44046 23662 44098
rect 23714 44046 23716 44098
rect 23660 43708 23716 44046
rect 25004 43708 25060 44270
rect 23324 43652 23492 43708
rect 23436 42980 23492 43652
rect 22988 40786 23044 40796
rect 23100 42700 23212 42756
rect 22876 40740 22932 40750
rect 21868 39618 22036 39620
rect 21868 39566 21870 39618
rect 21922 39566 22036 39618
rect 21868 39564 22036 39566
rect 22204 40626 22260 40638
rect 22204 40574 22206 40626
rect 22258 40574 22260 40626
rect 21868 39554 21924 39564
rect 21532 38994 21588 39004
rect 20860 38836 20916 38874
rect 20860 38770 20916 38780
rect 21308 38836 21364 38846
rect 21308 38742 21364 38780
rect 20636 38670 20638 38722
rect 20690 38670 20692 38722
rect 20636 38658 20692 38670
rect 20748 38276 20804 38286
rect 20636 37268 20692 37278
rect 20636 36370 20692 37212
rect 20748 36484 20804 38220
rect 21756 38276 21812 38286
rect 21756 38182 21812 38220
rect 21308 38052 21364 38062
rect 21308 37958 21364 37996
rect 22204 38052 22260 40574
rect 22876 40514 22932 40684
rect 22876 40462 22878 40514
rect 22930 40462 22932 40514
rect 22876 40450 22932 40462
rect 22540 40292 22596 40302
rect 22204 37986 22260 37996
rect 22428 40290 22596 40292
rect 22428 40238 22542 40290
rect 22594 40238 22596 40290
rect 22428 40236 22596 40238
rect 21980 37266 22036 37278
rect 21980 37214 21982 37266
rect 22034 37214 22036 37266
rect 21308 37154 21364 37166
rect 21308 37102 21310 37154
rect 21362 37102 21364 37154
rect 21308 36596 21364 37102
rect 21420 36596 21476 36606
rect 21308 36594 21476 36596
rect 21308 36542 21422 36594
rect 21474 36542 21476 36594
rect 21308 36540 21476 36542
rect 21420 36530 21476 36540
rect 21868 36594 21924 36606
rect 21868 36542 21870 36594
rect 21922 36542 21924 36594
rect 20748 36482 21028 36484
rect 20748 36430 20750 36482
rect 20802 36430 21028 36482
rect 20748 36428 21028 36430
rect 20748 36418 20804 36428
rect 20636 36318 20638 36370
rect 20690 36318 20692 36370
rect 20636 36306 20692 36318
rect 20524 34244 20580 34972
rect 20636 34916 20692 34926
rect 20636 34822 20692 34860
rect 20860 34580 20916 34590
rect 20748 34244 20804 34254
rect 20524 34242 20804 34244
rect 20524 34190 20750 34242
rect 20802 34190 20804 34242
rect 20524 34188 20804 34190
rect 20748 34178 20804 34188
rect 20860 34244 20916 34524
rect 20860 34150 20916 34188
rect 20412 33236 20468 33246
rect 20412 33142 20468 33180
rect 20860 33124 20916 33134
rect 20748 33122 20916 33124
rect 20748 33070 20862 33122
rect 20914 33070 20916 33122
rect 20748 33068 20916 33070
rect 20300 32620 20468 32676
rect 19572 32508 19684 32564
rect 19516 32498 19572 32508
rect 19404 31668 19460 31678
rect 19180 31666 19460 31668
rect 19180 31614 19406 31666
rect 19458 31614 19460 31666
rect 19180 31612 19460 31614
rect 18620 31554 18676 31566
rect 18620 31502 18622 31554
rect 18674 31502 18676 31554
rect 18620 31444 18676 31502
rect 18620 31378 18676 31388
rect 18508 30706 18564 30716
rect 19292 31108 19348 31612
rect 19404 31602 19460 31612
rect 19404 31444 19460 31454
rect 19460 31388 19572 31444
rect 19404 31378 19460 31388
rect 19068 30548 19124 30558
rect 19068 30210 19124 30492
rect 19292 30436 19348 31052
rect 19516 31106 19572 31388
rect 19516 31054 19518 31106
rect 19570 31054 19572 31106
rect 19516 31042 19572 31054
rect 19068 30158 19070 30210
rect 19122 30158 19124 30210
rect 19068 30146 19124 30158
rect 19180 30380 19348 30436
rect 19404 30772 19460 30782
rect 18508 29764 18564 29774
rect 18508 29652 18564 29708
rect 18508 29650 18788 29652
rect 18508 29598 18510 29650
rect 18562 29598 18788 29650
rect 18508 29596 18788 29598
rect 18508 29586 18564 29596
rect 18396 28354 18452 28364
rect 18732 29092 18788 29596
rect 18844 29316 18900 29326
rect 18956 29316 19012 29326
rect 18844 29314 18956 29316
rect 18844 29262 18846 29314
rect 18898 29262 18956 29314
rect 18844 29260 18956 29262
rect 18844 29250 18900 29260
rect 18732 28084 18788 29036
rect 18844 28084 18900 28094
rect 18732 28082 18900 28084
rect 18732 28030 18846 28082
rect 18898 28030 18900 28082
rect 18732 28028 18900 28030
rect 18844 28018 18900 28028
rect 18284 27122 18340 27132
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 18396 27186 18452 27806
rect 18396 27134 18398 27186
rect 18450 27134 18452 27186
rect 18396 27076 18452 27134
rect 18396 27010 18452 27020
rect 18620 27858 18676 27870
rect 18620 27806 18622 27858
rect 18674 27806 18676 27858
rect 17500 26852 18116 26908
rect 18620 26908 18676 27806
rect 18732 27748 18788 27758
rect 18732 27654 18788 27692
rect 18956 27636 19012 29260
rect 19068 28420 19124 28430
rect 19068 27858 19124 28364
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27794 19124 27806
rect 18956 27580 19124 27636
rect 19068 27186 19124 27580
rect 19068 27134 19070 27186
rect 19122 27134 19124 27186
rect 19068 27122 19124 27134
rect 18956 27076 19012 27114
rect 18956 27010 19012 27020
rect 19068 26964 19124 26974
rect 18620 26852 19124 26908
rect 17500 25844 17556 26852
rect 17612 26628 17668 26638
rect 17612 26516 17668 26572
rect 17612 26514 18004 26516
rect 17612 26462 17614 26514
rect 17666 26462 18004 26514
rect 17612 26460 18004 26462
rect 17612 26450 17668 26460
rect 17500 25618 17556 25788
rect 17500 25566 17502 25618
rect 17554 25566 17556 25618
rect 17500 25554 17556 25566
rect 17948 26402 18004 26460
rect 17948 26350 17950 26402
rect 18002 26350 18004 26402
rect 17724 24724 17780 24734
rect 17724 24630 17780 24668
rect 17948 23266 18004 26350
rect 18284 26292 18340 26302
rect 18284 26198 18340 26236
rect 18060 25508 18116 25518
rect 18060 25414 18116 25452
rect 18396 25506 18452 25518
rect 18396 25454 18398 25506
rect 18450 25454 18452 25506
rect 18396 24052 18452 25454
rect 18508 25508 18564 25518
rect 18620 25508 18676 26852
rect 18508 25506 18676 25508
rect 18508 25454 18510 25506
rect 18562 25454 18676 25506
rect 18508 25452 18676 25454
rect 18732 25844 18788 25854
rect 18732 25506 18788 25788
rect 18732 25454 18734 25506
rect 18786 25454 18788 25506
rect 18508 25442 18564 25452
rect 18732 25442 18788 25454
rect 18956 25732 19012 25742
rect 18956 25506 19012 25676
rect 18956 25454 18958 25506
rect 19010 25454 19012 25506
rect 18956 25442 19012 25454
rect 18620 25284 18676 25294
rect 19180 25284 19236 30380
rect 19404 30322 19460 30716
rect 19404 30270 19406 30322
rect 19458 30270 19460 30322
rect 19404 30258 19460 30270
rect 19516 30324 19572 30334
rect 19292 30212 19348 30222
rect 19292 30118 19348 30156
rect 19516 29986 19572 30268
rect 19628 30212 19684 32508
rect 19740 32562 20356 32564
rect 19740 32510 19742 32562
rect 19794 32510 20356 32562
rect 19740 32508 20356 32510
rect 19740 32498 19796 32508
rect 20188 32340 20244 32350
rect 19852 31892 19908 31902
rect 19852 31798 19908 31836
rect 20188 31778 20244 32284
rect 20188 31726 20190 31778
rect 20242 31726 20244 31778
rect 20188 31714 20244 31726
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 30996 20356 32508
rect 20412 31892 20468 32620
rect 20748 32564 20804 33068
rect 20860 33058 20916 33068
rect 20412 31826 20468 31836
rect 20524 32450 20580 32462
rect 20524 32398 20526 32450
rect 20578 32398 20580 32450
rect 20300 30902 20356 30940
rect 20412 31666 20468 31678
rect 20412 31614 20414 31666
rect 20466 31614 20468 31666
rect 20412 31556 20468 31614
rect 20412 30436 20468 31500
rect 20524 31554 20580 32398
rect 20524 31502 20526 31554
rect 20578 31502 20580 31554
rect 20524 31490 20580 31502
rect 20412 30380 20580 30436
rect 20524 30324 20580 30380
rect 20524 30258 20580 30268
rect 19628 30146 19684 30156
rect 20412 30212 20468 30222
rect 20412 30118 20468 30156
rect 19516 29934 19518 29986
rect 19570 29934 19572 29986
rect 19404 28420 19460 28430
rect 19292 26740 19348 26750
rect 19292 26292 19348 26684
rect 19292 25618 19348 26236
rect 19404 25732 19460 28364
rect 19516 27972 19572 29934
rect 19628 29988 19684 29998
rect 19628 29894 19684 29932
rect 20076 29988 20132 30026
rect 20076 29922 20132 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20636 29540 20692 29550
rect 20748 29540 20804 32508
rect 20860 32788 20916 32798
rect 20860 31778 20916 32732
rect 20860 31726 20862 31778
rect 20914 31726 20916 31778
rect 20860 31714 20916 31726
rect 20692 29484 20804 29540
rect 20860 30882 20916 30894
rect 20860 30830 20862 30882
rect 20914 30830 20916 30882
rect 20636 29474 20692 29484
rect 20300 29204 20356 29214
rect 20188 28756 20244 28766
rect 20188 28662 20244 28700
rect 19628 28644 19684 28654
rect 19628 28550 19684 28588
rect 20076 28420 20132 28458
rect 20076 28354 20132 28364
rect 20188 28418 20244 28430
rect 20188 28366 20190 28418
rect 20242 28366 20244 28418
rect 20188 28308 20244 28366
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 27878 19572 27916
rect 20188 27972 20244 28252
rect 20300 28084 20356 29148
rect 20860 28868 20916 30830
rect 20972 30660 21028 36428
rect 21868 36482 21924 36542
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36418 21924 36430
rect 21308 36260 21364 36270
rect 21308 36166 21364 36204
rect 21532 36260 21588 36270
rect 21532 36258 21700 36260
rect 21532 36206 21534 36258
rect 21586 36206 21700 36258
rect 21532 36204 21700 36206
rect 21532 36194 21588 36204
rect 21420 34804 21476 34814
rect 21420 34354 21476 34748
rect 21532 34692 21588 34702
rect 21532 34598 21588 34636
rect 21420 34302 21422 34354
rect 21474 34302 21476 34354
rect 21420 34290 21476 34302
rect 21084 34132 21140 34142
rect 21308 34132 21364 34142
rect 21532 34132 21588 34142
rect 21644 34132 21700 36204
rect 21868 35588 21924 35598
rect 21980 35588 22036 37214
rect 22092 36594 22148 36606
rect 22092 36542 22094 36594
rect 22146 36542 22148 36594
rect 22092 36484 22148 36542
rect 22316 36484 22372 36494
rect 22092 36482 22372 36484
rect 22092 36430 22318 36482
rect 22370 36430 22372 36482
rect 22092 36428 22372 36430
rect 22316 36418 22372 36428
rect 21868 35586 22036 35588
rect 21868 35534 21870 35586
rect 21922 35534 22036 35586
rect 21868 35532 22036 35534
rect 21084 34130 21364 34132
rect 21084 34078 21086 34130
rect 21138 34078 21310 34130
rect 21362 34078 21364 34130
rect 21084 34076 21364 34078
rect 21084 34066 21140 34076
rect 21308 34066 21364 34076
rect 21420 34130 21700 34132
rect 21420 34078 21534 34130
rect 21586 34078 21700 34130
rect 21420 34076 21700 34078
rect 21756 35252 21812 35262
rect 21420 33908 21476 34076
rect 21532 34066 21588 34076
rect 21420 32788 21476 33852
rect 21644 33572 21700 33582
rect 21756 33572 21812 35196
rect 21868 34916 21924 35532
rect 21868 34822 21924 34860
rect 21420 32722 21476 32732
rect 21532 33570 21812 33572
rect 21532 33518 21646 33570
rect 21698 33518 21812 33570
rect 21532 33516 21812 33518
rect 21868 34692 21924 34702
rect 21420 31892 21476 31902
rect 21308 31780 21364 31790
rect 21308 31686 21364 31724
rect 21420 31218 21476 31836
rect 21420 31166 21422 31218
rect 21474 31166 21476 31218
rect 21084 31108 21140 31118
rect 21084 31014 21140 31052
rect 21420 30772 21476 31166
rect 21420 30706 21476 30716
rect 20972 30604 21364 30660
rect 21308 30210 21364 30604
rect 21308 30158 21310 30210
rect 21362 30158 21364 30210
rect 21308 29876 21364 30158
rect 21532 30212 21588 33516
rect 21644 33506 21700 33516
rect 21868 33348 21924 34636
rect 21980 34132 22036 34142
rect 21980 34038 22036 34076
rect 22316 34130 22372 34142
rect 22316 34078 22318 34130
rect 22370 34078 22372 34130
rect 22316 34020 22372 34078
rect 21980 33572 22036 33582
rect 21980 33478 22036 33516
rect 21980 33348 22036 33358
rect 21868 33346 22036 33348
rect 21868 33294 21982 33346
rect 22034 33294 22036 33346
rect 21868 33292 22036 33294
rect 21980 33012 22036 33292
rect 21980 32946 22036 32956
rect 21756 30996 21812 31006
rect 21532 30146 21588 30156
rect 21644 30940 21756 30996
rect 21308 29810 21364 29820
rect 21420 29986 21476 29998
rect 21420 29934 21422 29986
rect 21474 29934 21476 29986
rect 21420 29652 21476 29934
rect 20972 29596 21476 29652
rect 21532 29986 21588 29998
rect 21532 29934 21534 29986
rect 21586 29934 21588 29986
rect 20972 29538 21028 29596
rect 20972 29486 20974 29538
rect 21026 29486 21028 29538
rect 20972 29474 21028 29486
rect 20860 28802 20916 28812
rect 21532 29316 21588 29934
rect 21644 29426 21700 30940
rect 21756 30902 21812 30940
rect 22316 30884 22372 33964
rect 22428 33348 22484 40236
rect 22540 40226 22596 40236
rect 22540 39506 22596 39518
rect 22540 39454 22542 39506
rect 22594 39454 22596 39506
rect 22540 38276 22596 39454
rect 22876 39060 22932 39070
rect 22876 38946 22932 39004
rect 23100 39060 23156 42700
rect 23212 42690 23268 42700
rect 23324 42924 23436 42980
rect 23324 40740 23380 42924
rect 23436 42914 23492 42924
rect 23548 43652 23604 43662
rect 23660 43652 23940 43708
rect 23548 42754 23604 43596
rect 23884 43650 23940 43652
rect 23884 43598 23886 43650
rect 23938 43598 23940 43650
rect 23884 43586 23940 43598
rect 24556 43652 25060 43708
rect 25676 44210 25732 44222
rect 25676 44158 25678 44210
rect 25730 44158 25732 44210
rect 25676 43708 25732 44158
rect 27804 43764 27860 44382
rect 29148 44436 29204 44446
rect 29820 44436 29876 47200
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 31276 44548 31332 44558
rect 31276 44546 31780 44548
rect 31276 44494 31278 44546
rect 31330 44494 31780 44546
rect 31276 44492 31780 44494
rect 31276 44482 31332 44492
rect 29148 44434 29876 44436
rect 29148 44382 29150 44434
rect 29202 44382 29876 44434
rect 29148 44380 29876 44382
rect 29148 44370 29204 44380
rect 29820 44324 29876 44380
rect 30044 44324 30100 44334
rect 29820 44322 30100 44324
rect 29820 44270 30046 44322
rect 30098 44270 30100 44322
rect 29820 44268 30100 44270
rect 30044 44258 30100 44268
rect 30604 44324 30660 44334
rect 30604 44230 30660 44268
rect 29708 44212 29764 44222
rect 30940 44212 30996 44222
rect 29708 44210 29988 44212
rect 29708 44158 29710 44210
rect 29762 44158 29988 44210
rect 29708 44156 29988 44158
rect 29708 44146 29764 44156
rect 28700 44100 28756 44110
rect 28700 44098 28868 44100
rect 28700 44046 28702 44098
rect 28754 44046 28868 44098
rect 28700 44044 28868 44046
rect 28700 44034 28756 44044
rect 25676 43652 25844 43708
rect 27804 43698 27860 43708
rect 28476 43876 28532 43886
rect 24556 43538 24612 43652
rect 24556 43486 24558 43538
rect 24610 43486 24612 43538
rect 23548 42702 23550 42754
rect 23602 42702 23604 42754
rect 23548 42690 23604 42702
rect 24332 42754 24388 42766
rect 24332 42702 24334 42754
rect 24386 42702 24388 42754
rect 24220 42532 24276 42542
rect 24108 42476 24220 42532
rect 23436 41076 23492 41086
rect 23436 40982 23492 41020
rect 23324 40684 23492 40740
rect 23212 40516 23268 40526
rect 23212 40422 23268 40460
rect 23100 38966 23156 39004
rect 23212 39508 23268 39518
rect 23212 39058 23268 39452
rect 23212 39006 23214 39058
rect 23266 39006 23268 39058
rect 23212 38994 23268 39006
rect 23436 39058 23492 40684
rect 23548 40628 23604 40638
rect 23548 40534 23604 40572
rect 23660 40402 23716 40414
rect 23660 40350 23662 40402
rect 23714 40350 23716 40402
rect 23436 39006 23438 39058
rect 23490 39006 23492 39058
rect 22876 38894 22878 38946
rect 22930 38894 22932 38946
rect 22876 38882 22932 38894
rect 23324 38948 23380 38958
rect 23324 38854 23380 38892
rect 23436 38668 23492 39006
rect 22540 38210 22596 38220
rect 22988 38612 23492 38668
rect 23548 40292 23604 40302
rect 22540 38052 22596 38062
rect 22540 37958 22596 37996
rect 22876 37492 22932 37502
rect 22988 37492 23044 38612
rect 22876 37490 23044 37492
rect 22876 37438 22878 37490
rect 22930 37438 23044 37490
rect 22876 37436 23044 37438
rect 22876 37426 22932 37436
rect 22652 37268 22708 37278
rect 22652 37266 23044 37268
rect 22652 37214 22654 37266
rect 22706 37214 23044 37266
rect 22652 37212 23044 37214
rect 22652 37202 22708 37212
rect 22652 36372 22708 36382
rect 22652 36370 22820 36372
rect 22652 36318 22654 36370
rect 22706 36318 22820 36370
rect 22652 36316 22820 36318
rect 22652 36306 22708 36316
rect 22540 36258 22596 36270
rect 22540 36206 22542 36258
rect 22594 36206 22596 36258
rect 22540 35812 22596 36206
rect 22540 35746 22596 35756
rect 22764 35028 22820 36316
rect 22876 36260 22932 36270
rect 22876 36166 22932 36204
rect 22988 35252 23044 37212
rect 23324 37266 23380 37278
rect 23324 37214 23326 37266
rect 23378 37214 23380 37266
rect 23212 36932 23268 36942
rect 23212 36482 23268 36876
rect 23212 36430 23214 36482
rect 23266 36430 23268 36482
rect 23212 36418 23268 36430
rect 23100 36260 23156 36270
rect 23100 36258 23268 36260
rect 23100 36206 23102 36258
rect 23154 36206 23268 36258
rect 23100 36204 23268 36206
rect 23100 36194 23156 36204
rect 22988 35186 23044 35196
rect 23212 35924 23268 36204
rect 22764 34972 23156 35028
rect 22540 34804 22596 34814
rect 22540 34802 23044 34804
rect 22540 34750 22542 34802
rect 22594 34750 23044 34802
rect 22540 34748 23044 34750
rect 22540 34738 22596 34748
rect 22652 34356 22708 34366
rect 22652 34262 22708 34300
rect 22988 34354 23044 34748
rect 22988 34302 22990 34354
rect 23042 34302 23044 34354
rect 22988 34290 23044 34302
rect 23100 34244 23156 34972
rect 23212 34580 23268 35868
rect 23212 34514 23268 34524
rect 23324 34356 23380 37214
rect 23548 37268 23604 40236
rect 23660 40180 23716 40350
rect 24108 40402 24164 42476
rect 24220 42466 24276 42476
rect 24220 41188 24276 41198
rect 24220 41094 24276 41132
rect 24332 40740 24388 42702
rect 24444 41972 24500 41982
rect 24444 40964 24500 41916
rect 24556 41188 24612 43486
rect 25004 43540 25060 43652
rect 25004 43474 25060 43484
rect 25228 43540 25284 43550
rect 25676 43540 25732 43550
rect 25228 43538 25620 43540
rect 25228 43486 25230 43538
rect 25282 43486 25620 43538
rect 25228 43484 25620 43486
rect 25228 43474 25284 43484
rect 25340 43314 25396 43326
rect 25340 43262 25342 43314
rect 25394 43262 25396 43314
rect 24780 42866 24836 42878
rect 24780 42814 24782 42866
rect 24834 42814 24836 42866
rect 24668 42644 24724 42654
rect 24668 41300 24724 42588
rect 24780 42532 24836 42814
rect 24780 42466 24836 42476
rect 25340 41412 25396 43262
rect 25564 42980 25620 43484
rect 25676 43446 25732 43484
rect 25788 43204 25844 43652
rect 26460 43428 26516 43438
rect 26460 43334 26516 43372
rect 25788 43138 25844 43148
rect 26684 42980 26740 42990
rect 25564 42924 26516 42980
rect 26460 42866 26516 42924
rect 26460 42814 26462 42866
rect 26514 42814 26516 42866
rect 26460 42802 26516 42814
rect 26348 42756 26404 42766
rect 26348 42662 26404 42700
rect 26684 42754 26740 42924
rect 26684 42702 26686 42754
rect 26738 42702 26740 42754
rect 26684 42690 26740 42702
rect 26124 42644 26180 42654
rect 26124 42550 26180 42588
rect 28476 42644 28532 43820
rect 28700 43540 28756 43550
rect 28588 43484 28700 43540
rect 28588 43426 28644 43484
rect 28700 43474 28756 43484
rect 28588 43374 28590 43426
rect 28642 43374 28644 43426
rect 28588 43362 28644 43374
rect 28476 42578 28532 42588
rect 26572 42530 26628 42542
rect 27356 42532 27412 42542
rect 26572 42478 26574 42530
rect 26626 42478 26628 42530
rect 26572 42420 26628 42478
rect 26572 42354 26628 42364
rect 27244 42530 27412 42532
rect 27244 42478 27358 42530
rect 27410 42478 27412 42530
rect 27244 42476 27412 42478
rect 25340 41346 25396 41356
rect 27132 41412 27188 41422
rect 24668 41298 25060 41300
rect 24668 41246 24670 41298
rect 24722 41246 25060 41298
rect 24668 41244 25060 41246
rect 24668 41234 24724 41244
rect 24556 41122 24612 41132
rect 24556 40964 24612 40974
rect 24444 40962 24612 40964
rect 24444 40910 24558 40962
rect 24610 40910 24612 40962
rect 24444 40908 24612 40910
rect 24556 40898 24612 40908
rect 24332 40628 24388 40684
rect 24444 40628 24500 40638
rect 24332 40626 24500 40628
rect 24332 40574 24446 40626
rect 24498 40574 24500 40626
rect 24332 40572 24500 40574
rect 24444 40562 24500 40572
rect 24108 40350 24110 40402
rect 24162 40350 24164 40402
rect 24108 40338 24164 40350
rect 24332 40180 24388 40190
rect 23716 40124 23828 40180
rect 23660 40114 23716 40124
rect 23660 39060 23716 39070
rect 23660 37490 23716 39004
rect 23660 37438 23662 37490
rect 23714 37438 23716 37490
rect 23660 37426 23716 37438
rect 23548 37212 23716 37268
rect 23548 36932 23604 36942
rect 23548 36482 23604 36876
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 36418 23604 36430
rect 23660 36370 23716 37212
rect 23660 36318 23662 36370
rect 23714 36318 23716 36370
rect 23660 36306 23716 36318
rect 23772 35924 23828 40124
rect 24108 39060 24164 39070
rect 24108 38946 24164 39004
rect 24332 39058 24388 40124
rect 24668 39732 24724 39742
rect 24332 39006 24334 39058
rect 24386 39006 24388 39058
rect 24332 38994 24388 39006
rect 24556 39730 24724 39732
rect 24556 39678 24670 39730
rect 24722 39678 24724 39730
rect 24556 39676 24724 39678
rect 24108 38894 24110 38946
rect 24162 38894 24164 38946
rect 24108 38882 24164 38894
rect 24444 38836 24500 38846
rect 24556 38836 24612 39676
rect 24668 39666 24724 39676
rect 25004 39730 25060 41244
rect 25340 41188 25396 41198
rect 25340 41094 25396 41132
rect 26012 41074 26068 41086
rect 26012 41022 26014 41074
rect 26066 41022 26068 41074
rect 26012 40628 26068 41022
rect 26012 40562 26068 40572
rect 25228 40292 25284 40302
rect 25004 39678 25006 39730
rect 25058 39678 25060 39730
rect 25004 39666 25060 39678
rect 25116 40290 25284 40292
rect 25116 40238 25230 40290
rect 25282 40238 25284 40290
rect 25116 40236 25284 40238
rect 25116 39172 25172 40236
rect 25228 40226 25284 40236
rect 27132 39730 27188 41356
rect 27132 39678 27134 39730
rect 27186 39678 27188 39730
rect 27132 39666 27188 39678
rect 27244 39508 27300 42476
rect 27356 42466 27412 42476
rect 27804 42530 27860 42542
rect 27804 42478 27806 42530
rect 27858 42478 27860 42530
rect 27692 40964 27748 40974
rect 27580 40908 27692 40964
rect 27356 40404 27412 40414
rect 27356 40310 27412 40348
rect 27132 39452 27300 39508
rect 24668 39116 25116 39172
rect 24668 38946 24724 39116
rect 25116 39078 25172 39116
rect 26572 39284 26628 39294
rect 24668 38894 24670 38946
rect 24722 38894 24724 38946
rect 24668 38882 24724 38894
rect 26348 39060 26404 39070
rect 24500 38780 24612 38836
rect 25116 38836 25172 38846
rect 24444 38742 24500 38780
rect 24332 38724 24388 38734
rect 23884 38276 23940 38286
rect 23940 38220 24052 38276
rect 23884 38210 23940 38220
rect 23884 37938 23940 37950
rect 23884 37886 23886 37938
rect 23938 37886 23940 37938
rect 23884 36482 23940 37886
rect 23996 37044 24052 38220
rect 24108 37380 24164 37390
rect 24108 37286 24164 37324
rect 24220 37380 24276 37390
rect 24332 37380 24388 38668
rect 25116 38162 25172 38780
rect 25900 38834 25956 38846
rect 25900 38782 25902 38834
rect 25954 38782 25956 38834
rect 25228 38724 25284 38734
rect 25900 38668 25956 38782
rect 25228 38630 25284 38668
rect 25116 38110 25118 38162
rect 25170 38110 25172 38162
rect 25116 38098 25172 38110
rect 25452 38612 25956 38668
rect 26124 38724 26180 38734
rect 26124 38630 26180 38668
rect 25452 38162 25508 38612
rect 25452 38110 25454 38162
rect 25506 38110 25508 38162
rect 24220 37378 24388 37380
rect 24220 37326 24222 37378
rect 24274 37326 24388 37378
rect 24220 37324 24388 37326
rect 24444 38050 24500 38062
rect 24444 37998 24446 38050
rect 24498 37998 24500 38050
rect 24220 37314 24276 37324
rect 24444 37268 24500 37998
rect 25452 38052 25508 38110
rect 25452 37986 25508 37996
rect 25788 38050 25844 38062
rect 25788 37998 25790 38050
rect 25842 37998 25844 38050
rect 24668 37268 24724 37278
rect 24444 37212 24668 37268
rect 24668 37174 24724 37212
rect 25452 37156 25508 37166
rect 25788 37156 25844 37998
rect 26012 37826 26068 37838
rect 26012 37774 26014 37826
rect 26066 37774 26068 37826
rect 26012 37268 26068 37774
rect 26124 37268 26180 37278
rect 26012 37266 26292 37268
rect 26012 37214 26126 37266
rect 26178 37214 26292 37266
rect 26012 37212 26292 37214
rect 26124 37202 26180 37212
rect 25452 37154 25844 37156
rect 25452 37102 25454 37154
rect 25506 37102 25844 37154
rect 25452 37100 25844 37102
rect 24108 37044 24164 37054
rect 23996 37042 24164 37044
rect 23996 36990 24110 37042
rect 24162 36990 24164 37042
rect 23996 36988 24164 36990
rect 24108 36978 24164 36988
rect 25452 37044 25508 37100
rect 25452 36978 25508 36988
rect 23884 36430 23886 36482
rect 23938 36430 23940 36482
rect 23884 36418 23940 36430
rect 26012 36370 26068 36382
rect 26012 36318 26014 36370
rect 26066 36318 26068 36370
rect 23100 34132 23156 34188
rect 22988 34076 23156 34132
rect 23212 34300 23380 34356
rect 23548 35868 23772 35924
rect 22988 33348 23044 34076
rect 23100 33908 23156 33918
rect 23100 33814 23156 33852
rect 23212 33572 23268 34300
rect 23324 34132 23380 34142
rect 23548 34132 23604 35868
rect 23772 35858 23828 35868
rect 24444 36258 24500 36270
rect 24444 36206 24446 36258
rect 24498 36206 24500 36258
rect 24444 35308 24500 36206
rect 25228 36260 25284 36270
rect 26012 36260 26068 36318
rect 25228 36258 26068 36260
rect 25228 36206 25230 36258
rect 25282 36206 26068 36258
rect 25228 36204 26068 36206
rect 25228 36194 25284 36204
rect 25228 35924 25284 35934
rect 25228 35830 25284 35868
rect 25340 35700 25396 35710
rect 24220 35252 24500 35308
rect 24668 35698 25396 35700
rect 24668 35646 25342 35698
rect 25394 35646 25396 35698
rect 24668 35644 25396 35646
rect 23324 34130 23604 34132
rect 23324 34078 23326 34130
rect 23378 34078 23604 34130
rect 23324 34076 23604 34078
rect 23772 34356 23828 34366
rect 23772 34130 23828 34300
rect 23772 34078 23774 34130
rect 23826 34078 23828 34130
rect 23324 34066 23380 34076
rect 23772 34066 23828 34078
rect 24108 34132 24164 34142
rect 24108 34038 24164 34076
rect 23884 33908 23940 33918
rect 23884 33814 23940 33852
rect 23212 33506 23268 33516
rect 23996 33796 24052 33806
rect 22428 33346 22708 33348
rect 22428 33294 22430 33346
rect 22482 33294 22708 33346
rect 22428 33292 22708 33294
rect 22428 33282 22484 33292
rect 22540 33122 22596 33134
rect 22540 33070 22542 33122
rect 22594 33070 22596 33122
rect 22540 32900 22596 33070
rect 22428 32844 22596 32900
rect 22428 32340 22484 32844
rect 22652 32450 22708 33292
rect 22988 33346 23380 33348
rect 22988 33294 22990 33346
rect 23042 33294 23380 33346
rect 22988 33292 23380 33294
rect 22988 33282 23044 33292
rect 22764 33236 22820 33246
rect 22764 33142 22820 33180
rect 23324 33234 23380 33292
rect 23324 33182 23326 33234
rect 23378 33182 23380 33234
rect 23324 33170 23380 33182
rect 23436 33236 23492 33246
rect 23324 32788 23380 32798
rect 22652 32398 22654 32450
rect 22706 32398 22708 32450
rect 22652 32386 22708 32398
rect 22764 32786 23380 32788
rect 22764 32734 23326 32786
rect 23378 32734 23380 32786
rect 22764 32732 23380 32734
rect 22428 32274 22484 32284
rect 22540 31108 22596 31118
rect 22764 31108 22820 32732
rect 23324 32722 23380 32732
rect 22988 32564 23044 32574
rect 22988 32470 23044 32508
rect 23324 32564 23380 32574
rect 23324 32470 23380 32508
rect 23436 32340 23492 33180
rect 23660 33122 23716 33134
rect 23884 33124 23940 33134
rect 23660 33070 23662 33122
rect 23714 33070 23716 33122
rect 22540 31106 22820 31108
rect 22540 31054 22542 31106
rect 22594 31054 22820 31106
rect 22540 31052 22820 31054
rect 23212 31668 23268 31678
rect 22540 31042 22596 31052
rect 22316 30828 23156 30884
rect 22316 30324 22372 30334
rect 21980 30210 22036 30222
rect 21980 30158 21982 30210
rect 22034 30158 22036 30210
rect 21644 29374 21646 29426
rect 21698 29374 21700 29426
rect 21644 29362 21700 29374
rect 21756 29876 21812 29886
rect 20636 28642 20692 28654
rect 20636 28590 20638 28642
rect 20690 28590 20692 28642
rect 20300 28018 20356 28028
rect 20412 28418 20468 28430
rect 20412 28366 20414 28418
rect 20466 28366 20468 28418
rect 20188 27906 20244 27916
rect 19852 27746 19908 27758
rect 19852 27694 19854 27746
rect 19906 27694 19908 27746
rect 19740 27186 19796 27198
rect 19740 27134 19742 27186
rect 19794 27134 19796 27186
rect 19628 26962 19684 26974
rect 19628 26910 19630 26962
rect 19682 26910 19684 26962
rect 19628 26290 19684 26910
rect 19740 26852 19796 27134
rect 19852 27076 19908 27694
rect 20076 27076 20132 27086
rect 19852 27074 20132 27076
rect 19852 27022 20078 27074
rect 20130 27022 20132 27074
rect 19852 27020 20132 27022
rect 19740 26786 19796 26796
rect 20076 26852 20132 27020
rect 20412 26964 20468 28366
rect 20636 27636 20692 28590
rect 20636 27570 20692 27580
rect 20748 28644 20804 28654
rect 20412 26898 20468 26908
rect 20076 26786 20132 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26226 19684 26238
rect 19404 25666 19460 25676
rect 20412 26180 20468 26190
rect 20188 25620 20244 25630
rect 19292 25566 19294 25618
rect 19346 25566 19348 25618
rect 19292 25554 19348 25566
rect 20076 25564 20188 25620
rect 19404 25508 19460 25518
rect 19852 25508 19908 25518
rect 19404 25506 19908 25508
rect 19404 25454 19406 25506
rect 19458 25454 19854 25506
rect 19906 25454 19908 25506
rect 19404 25452 19908 25454
rect 19404 25442 19460 25452
rect 19852 25442 19908 25452
rect 20076 25506 20132 25564
rect 20188 25554 20244 25564
rect 20412 25618 20468 26124
rect 20412 25566 20414 25618
rect 20466 25566 20468 25618
rect 20412 25554 20468 25566
rect 20524 26178 20580 26190
rect 20524 26126 20526 26178
rect 20578 26126 20580 26178
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 20076 25442 20132 25454
rect 20300 25508 20356 25518
rect 20524 25508 20580 26126
rect 20524 25452 20692 25508
rect 19180 25228 19572 25284
rect 18620 25190 18676 25228
rect 18508 24052 18564 24062
rect 18396 24050 18676 24052
rect 18396 23998 18510 24050
rect 18562 23998 18676 24050
rect 18396 23996 18676 23998
rect 18508 23986 18564 23996
rect 17948 23214 17950 23266
rect 18002 23214 18004 23266
rect 17724 23042 17780 23054
rect 17724 22990 17726 23042
rect 17778 22990 17780 23042
rect 17724 22932 17780 22990
rect 17724 22866 17780 22876
rect 17948 22482 18004 23214
rect 18284 23156 18340 23166
rect 18284 23062 18340 23100
rect 17948 22430 17950 22482
rect 18002 22430 18004 22482
rect 17164 22306 17220 22316
rect 17724 22372 17780 22382
rect 17724 21812 17780 22316
rect 17612 21810 17780 21812
rect 17612 21758 17726 21810
rect 17778 21758 17780 21810
rect 17612 21756 17780 21758
rect 17388 21698 17444 21710
rect 17388 21646 17390 21698
rect 17442 21646 17444 21698
rect 17388 20356 17444 21646
rect 17388 20290 17444 20300
rect 17164 20244 17220 20254
rect 17052 20132 17108 20142
rect 17052 19234 17108 20076
rect 17052 19182 17054 19234
rect 17106 19182 17108 19234
rect 17052 19170 17108 19182
rect 17164 19122 17220 20188
rect 17612 20242 17668 21756
rect 17724 21746 17780 21756
rect 17948 21812 18004 22430
rect 18508 22482 18564 22494
rect 18508 22430 18510 22482
rect 18562 22430 18564 22482
rect 17948 21746 18004 21756
rect 18396 21812 18452 21822
rect 18396 21586 18452 21756
rect 18396 21534 18398 21586
rect 18450 21534 18452 21586
rect 18396 21522 18452 21534
rect 18508 21364 18564 22430
rect 18620 22370 18676 23996
rect 19180 23940 19236 23950
rect 19404 23940 19460 23950
rect 19180 23938 19460 23940
rect 19180 23886 19182 23938
rect 19234 23886 19406 23938
rect 19458 23886 19460 23938
rect 19180 23884 19460 23886
rect 19180 23874 19236 23884
rect 19404 23874 19460 23884
rect 19068 23826 19124 23838
rect 19068 23774 19070 23826
rect 19122 23774 19124 23826
rect 19068 23156 19124 23774
rect 19124 23100 19348 23156
rect 19068 23062 19124 23100
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22306 18676 22318
rect 19180 22484 19236 22494
rect 18844 21700 18900 21710
rect 19180 21700 19236 22428
rect 19292 22482 19348 23100
rect 19292 22430 19294 22482
rect 19346 22430 19348 22482
rect 19292 22418 19348 22430
rect 18844 21698 19236 21700
rect 18844 21646 18846 21698
rect 18898 21646 19236 21698
rect 18844 21644 19236 21646
rect 18844 21634 18900 21644
rect 19180 21474 19236 21644
rect 19180 21422 19182 21474
rect 19234 21422 19236 21474
rect 19180 21410 19236 21422
rect 18508 21298 18564 21308
rect 18732 21364 18788 21374
rect 18732 21362 19124 21364
rect 18732 21310 18734 21362
rect 18786 21310 19124 21362
rect 18732 21308 19124 21310
rect 18732 21298 18788 21308
rect 18172 20914 18228 20926
rect 18172 20862 18174 20914
rect 18226 20862 18228 20914
rect 18172 20804 18228 20862
rect 18228 20748 18340 20804
rect 18172 20738 18228 20748
rect 17612 20190 17614 20242
rect 17666 20190 17668 20242
rect 17612 20178 17668 20190
rect 18172 20244 18228 20254
rect 17836 20132 17892 20142
rect 17836 20038 17892 20076
rect 18172 20130 18228 20188
rect 18172 20078 18174 20130
rect 18226 20078 18228 20130
rect 17948 19908 18004 19918
rect 17948 19814 18004 19852
rect 18172 19796 18228 20078
rect 18284 20018 18340 20748
rect 19068 20802 19124 21308
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 18956 20690 19012 20702
rect 18956 20638 18958 20690
rect 19010 20638 19012 20690
rect 18508 20580 18564 20590
rect 18508 20486 18564 20524
rect 18956 20580 19012 20638
rect 18284 19966 18286 20018
rect 18338 19966 18340 20018
rect 18284 19954 18340 19966
rect 18620 20132 18676 20142
rect 18172 19740 18340 19796
rect 18172 19348 18228 19358
rect 17948 19292 18172 19348
rect 17388 19236 17444 19246
rect 17836 19236 17892 19246
rect 17388 19234 17892 19236
rect 17388 19182 17390 19234
rect 17442 19182 17838 19234
rect 17890 19182 17892 19234
rect 17388 19180 17892 19182
rect 17388 19170 17444 19180
rect 17836 19170 17892 19180
rect 17164 19070 17166 19122
rect 17218 19070 17220 19122
rect 17164 19058 17220 19070
rect 17948 19012 18004 19292
rect 18172 19254 18228 19292
rect 17724 18956 18004 19012
rect 17724 18674 17780 18956
rect 17724 18622 17726 18674
rect 17778 18622 17780 18674
rect 17724 18610 17780 18622
rect 17388 18562 17444 18574
rect 17388 18510 17390 18562
rect 17442 18510 17444 18562
rect 17388 18116 17444 18510
rect 17388 18050 17444 18060
rect 17500 18564 17556 18574
rect 17500 17106 17556 18508
rect 18284 18562 18340 19740
rect 18284 18510 18286 18562
rect 18338 18510 18340 18562
rect 18284 18498 18340 18510
rect 18620 18450 18676 20076
rect 18956 20132 19012 20524
rect 19068 20244 19124 20750
rect 19180 20804 19236 20814
rect 19180 20710 19236 20748
rect 19068 20178 19124 20188
rect 19292 20244 19348 20254
rect 18956 20066 19012 20076
rect 19292 20130 19348 20188
rect 19292 20078 19294 20130
rect 19346 20078 19348 20130
rect 18844 19906 18900 19918
rect 18844 19854 18846 19906
rect 18898 19854 18900 19906
rect 18844 18788 18900 19854
rect 19292 19012 19348 20078
rect 19516 20132 19572 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 23940 19684 23950
rect 19852 23940 19908 23950
rect 19628 23938 19908 23940
rect 19628 23886 19630 23938
rect 19682 23886 19854 23938
rect 19906 23886 19908 23938
rect 19628 23884 19908 23886
rect 19628 23874 19684 23884
rect 19852 23874 19908 23884
rect 20076 23938 20132 23950
rect 20076 23886 20078 23938
rect 20130 23886 20132 23938
rect 20076 23716 20132 23886
rect 20300 23938 20356 25452
rect 20524 25282 20580 25294
rect 20524 25230 20526 25282
rect 20578 25230 20580 25282
rect 20524 25172 20580 25230
rect 20524 25106 20580 25116
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 20300 23874 20356 23886
rect 20412 23716 20468 23726
rect 20076 23660 20244 23716
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23492 20244 23660
rect 20412 23622 20468 23660
rect 20524 23714 20580 23726
rect 20524 23662 20526 23714
rect 20578 23662 20580 23714
rect 20524 23604 20580 23662
rect 20524 23538 20580 23548
rect 20188 23436 20356 23492
rect 20188 23266 20244 23278
rect 20188 23214 20190 23266
rect 20242 23214 20244 23266
rect 19628 23154 19684 23166
rect 19628 23102 19630 23154
rect 19682 23102 19684 23154
rect 19628 22594 19684 23102
rect 19628 22542 19630 22594
rect 19682 22542 19684 22594
rect 19628 22530 19684 22542
rect 19740 22596 19796 22606
rect 19740 22370 19796 22540
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19740 22306 19796 22318
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19852 20804 19908 20814
rect 19852 20710 19908 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 23214
rect 20300 22820 20356 23436
rect 20636 23380 20692 25452
rect 20300 22754 20356 22764
rect 20412 23324 20692 23380
rect 20748 23828 20804 28588
rect 21532 28532 21588 29260
rect 21644 28868 21700 28878
rect 21644 28754 21700 28812
rect 21644 28702 21646 28754
rect 21698 28702 21700 28754
rect 21644 28690 21700 28702
rect 21532 28466 21588 28476
rect 21756 27972 21812 29820
rect 21980 28868 22036 30158
rect 22316 29204 22372 30268
rect 22764 30212 22820 30250
rect 22764 30146 22820 30156
rect 22988 30210 23044 30222
rect 22988 30158 22990 30210
rect 23042 30158 23044 30210
rect 22428 29988 22484 29998
rect 22428 29894 22484 29932
rect 22764 29988 22820 29998
rect 22428 29428 22484 29438
rect 22428 29334 22484 29372
rect 22652 29314 22708 29326
rect 22652 29262 22654 29314
rect 22706 29262 22708 29314
rect 22428 29204 22484 29214
rect 22316 29148 22428 29204
rect 22428 29138 22484 29148
rect 21980 28802 22036 28812
rect 21980 28644 22036 28654
rect 21756 27906 21812 27916
rect 21868 28642 22036 28644
rect 21868 28590 21982 28642
rect 22034 28590 22036 28642
rect 21868 28588 22036 28590
rect 21420 27074 21476 27086
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 21420 26908 21476 27022
rect 21308 26852 21364 26862
rect 21420 26852 21588 26908
rect 21196 26404 21252 26414
rect 21084 26402 21252 26404
rect 21084 26350 21198 26402
rect 21250 26350 21252 26402
rect 21084 26348 21252 26350
rect 20412 22484 20468 23324
rect 20636 23156 20692 23166
rect 20636 23062 20692 23100
rect 20748 22932 20804 23772
rect 20636 22876 20804 22932
rect 20972 25508 21028 25518
rect 20300 22428 20468 22484
rect 20524 22596 20580 22606
rect 20300 20804 20356 22428
rect 20524 22372 20580 22540
rect 20412 22316 20580 22372
rect 20412 22258 20468 22316
rect 20412 22206 20414 22258
rect 20466 22206 20468 22258
rect 20412 22194 20468 22206
rect 20524 22146 20580 22158
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20524 21026 20580 22094
rect 20524 20974 20526 21026
rect 20578 20974 20580 21026
rect 20524 20962 20580 20974
rect 20300 20748 20468 20804
rect 20300 20578 20356 20590
rect 20300 20526 20302 20578
rect 20354 20526 20356 20578
rect 20300 20468 20356 20526
rect 20300 20402 20356 20412
rect 20188 20178 20244 20188
rect 20076 20132 20132 20142
rect 19516 20130 20132 20132
rect 19516 20078 20078 20130
rect 20130 20078 20132 20130
rect 19516 20076 20132 20078
rect 20076 19460 20132 20076
rect 20076 19394 20132 19404
rect 20412 19348 20468 20748
rect 20524 20132 20580 20142
rect 20524 20018 20580 20076
rect 20524 19966 20526 20018
rect 20578 19966 20580 20018
rect 20524 19954 20580 19966
rect 20412 19282 20468 19292
rect 18844 18722 18900 18732
rect 19068 18956 19348 19012
rect 19516 19234 19572 19246
rect 19516 19182 19518 19234
rect 19570 19182 19572 19234
rect 18620 18398 18622 18450
rect 18674 18398 18676 18450
rect 18620 18386 18676 18398
rect 19068 18450 19124 18956
rect 19516 18788 19572 19182
rect 19964 19122 20020 19134
rect 19964 19070 19966 19122
rect 20018 19070 20020 19122
rect 19964 19012 20020 19070
rect 20412 19124 20468 19134
rect 20412 19030 20468 19068
rect 19516 18722 19572 18732
rect 19628 18956 20356 19012
rect 19404 18562 19460 18574
rect 19404 18510 19406 18562
rect 19458 18510 19460 18562
rect 19292 18452 19348 18462
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 18386 19124 18398
rect 19180 18396 19292 18452
rect 18732 18338 18788 18350
rect 18732 18286 18734 18338
rect 18786 18286 18788 18338
rect 17500 17054 17502 17106
rect 17554 17054 17556 17106
rect 17500 16996 17556 17054
rect 17500 16930 17556 16940
rect 18284 18116 18340 18126
rect 18284 16882 18340 18060
rect 18284 16830 18286 16882
rect 18338 16830 18340 16882
rect 18284 16818 18340 16830
rect 18396 16884 18452 16894
rect 17948 16772 18004 16782
rect 17724 16770 18004 16772
rect 17724 16718 17950 16770
rect 18002 16718 18004 16770
rect 17724 16716 18004 16718
rect 17724 16322 17780 16716
rect 17948 16706 18004 16716
rect 18172 16770 18228 16782
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 18172 16548 18228 16718
rect 17724 16270 17726 16322
rect 17778 16270 17780 16322
rect 16940 16046 16942 16098
rect 16994 16046 16996 16098
rect 15820 14868 15876 14878
rect 15820 14642 15876 14812
rect 15820 14590 15822 14642
rect 15874 14590 15876 14642
rect 15820 14578 15876 14590
rect 16268 14642 16324 15148
rect 16268 14590 16270 14642
rect 16322 14590 16324 14642
rect 16268 14578 16324 14590
rect 16492 15092 16772 15148
rect 16828 15540 16884 15550
rect 16940 15540 16996 16046
rect 17500 16098 17556 16110
rect 17500 16046 17502 16098
rect 17554 16046 17556 16098
rect 17500 15764 17556 16046
rect 17724 16100 17780 16270
rect 17724 16034 17780 16044
rect 17836 16492 18228 16548
rect 17836 15988 17892 16492
rect 18396 16322 18452 16828
rect 18396 16270 18398 16322
rect 18450 16270 18452 16322
rect 18396 16258 18452 16270
rect 17612 15764 17668 15774
rect 17500 15708 17612 15764
rect 16828 15538 16996 15540
rect 16828 15486 16830 15538
rect 16882 15486 16996 15538
rect 16828 15484 16996 15486
rect 17612 15538 17668 15708
rect 17836 15652 17892 15932
rect 17836 15586 17892 15596
rect 17948 16212 18004 16222
rect 17612 15486 17614 15538
rect 17666 15486 17668 15538
rect 14924 14478 14926 14530
rect 14978 14478 14980 14530
rect 14924 14466 14980 14478
rect 15484 14530 15540 14542
rect 15484 14478 15486 14530
rect 15538 14478 15540 14530
rect 14700 14308 14756 14318
rect 14700 14306 14980 14308
rect 14700 14254 14702 14306
rect 14754 14254 14980 14306
rect 14700 14252 14980 14254
rect 14700 14242 14756 14252
rect 14588 14018 14644 14028
rect 14924 14196 14980 14252
rect 15484 14196 15540 14478
rect 14924 14140 15540 14196
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13682 14084 13694
rect 14700 13858 14756 13870
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13748 14756 13806
rect 14700 13682 14756 13692
rect 14924 13746 14980 14140
rect 15484 13972 15540 14140
rect 15708 13972 15764 13982
rect 16156 13972 16212 13982
rect 15484 13970 16212 13972
rect 15484 13918 15710 13970
rect 15762 13918 16158 13970
rect 16210 13918 16212 13970
rect 15484 13916 16212 13918
rect 15708 13906 15764 13916
rect 16156 13906 16212 13916
rect 14924 13694 14926 13746
rect 14978 13694 14980 13746
rect 14924 13682 14980 13694
rect 15372 13858 15428 13870
rect 15372 13806 15374 13858
rect 15426 13806 15428 13858
rect 12908 13522 12964 13534
rect 12908 13470 12910 13522
rect 12962 13470 12964 13522
rect 12908 13188 12964 13470
rect 12908 13122 12964 13132
rect 13692 13188 13748 13198
rect 12908 12964 12964 12974
rect 12908 12870 12964 12908
rect 13692 12962 13748 13132
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 13468 12738 13524 12750
rect 13804 12740 13860 13580
rect 14252 12964 14308 12974
rect 14308 12908 14532 12964
rect 14252 12870 14308 12908
rect 13468 12686 13470 12738
rect 13522 12686 13524 12738
rect 13468 12290 13524 12686
rect 13468 12238 13470 12290
rect 13522 12238 13524 12290
rect 13468 12226 13524 12238
rect 13580 12684 13804 12740
rect 12908 11284 12964 11294
rect 12908 11190 12964 11228
rect 13356 11284 13412 11294
rect 13356 11190 13412 11228
rect 13580 11282 13636 12684
rect 13804 12674 13860 12684
rect 13580 11230 13582 11282
rect 13634 11230 13636 11282
rect 13580 11218 13636 11230
rect 13692 11284 13748 11294
rect 13692 11190 13748 11228
rect 12908 10500 12964 10510
rect 12964 10444 13188 10500
rect 12908 10434 12964 10444
rect 13020 9940 13076 9950
rect 13020 9266 13076 9884
rect 13020 9214 13022 9266
rect 13074 9214 13076 9266
rect 13020 8932 13076 9214
rect 13020 8866 13076 8876
rect 13132 8932 13188 10444
rect 14476 9938 14532 12908
rect 15372 12292 15428 13806
rect 16380 12962 16436 12974
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 15932 12404 15988 12414
rect 16156 12404 16212 12414
rect 15932 12402 16156 12404
rect 15932 12350 15934 12402
rect 15986 12350 16156 12402
rect 15932 12348 16156 12350
rect 15372 12236 15764 12292
rect 15596 12066 15652 12078
rect 15596 12014 15598 12066
rect 15650 12014 15652 12066
rect 15596 11732 15652 12014
rect 15708 11788 15764 12236
rect 15820 11788 15876 11798
rect 15708 11732 15820 11788
rect 15484 11676 15652 11732
rect 15820 11722 15876 11732
rect 15484 11620 15540 11676
rect 15484 11554 15540 11564
rect 15820 11620 15876 11630
rect 15484 11396 15540 11406
rect 15260 11284 15316 11294
rect 15260 11190 15316 11228
rect 15372 11284 15428 11294
rect 15484 11284 15540 11340
rect 15372 11282 15540 11284
rect 15372 11230 15374 11282
rect 15426 11230 15540 11282
rect 15372 11228 15540 11230
rect 15372 11218 15428 11228
rect 14924 11172 14980 11182
rect 15148 11172 15204 11182
rect 14924 11170 15092 11172
rect 14924 11118 14926 11170
rect 14978 11118 15092 11170
rect 14924 11116 15092 11118
rect 14924 11106 14980 11116
rect 15036 10836 15092 11116
rect 15148 10948 15204 11116
rect 15148 10892 15316 10948
rect 15036 10780 15204 10836
rect 14700 10500 14756 10510
rect 15036 10500 15092 10510
rect 14700 10498 15092 10500
rect 14700 10446 14702 10498
rect 14754 10446 15038 10498
rect 15090 10446 15092 10498
rect 14700 10444 15092 10446
rect 14700 10434 14756 10444
rect 15036 10434 15092 10444
rect 15148 10388 15204 10780
rect 15260 10612 15316 10892
rect 15484 10722 15540 11228
rect 15596 11394 15652 11406
rect 15596 11342 15598 11394
rect 15650 11342 15652 11394
rect 15596 11284 15652 11342
rect 15596 11218 15652 11228
rect 15820 10948 15876 11564
rect 15932 11508 15988 12348
rect 16156 12338 16212 12348
rect 16268 12292 16324 12302
rect 16268 11620 16324 12236
rect 16380 11956 16436 12910
rect 16492 12068 16548 15092
rect 16716 13748 16772 13758
rect 16828 13748 16884 15484
rect 17612 15474 17668 15486
rect 17948 15426 18004 16156
rect 18732 16212 18788 18286
rect 19180 16884 19236 18396
rect 19292 18386 19348 18396
rect 19404 18116 19460 18510
rect 19404 18050 19460 18060
rect 19516 18564 19572 18574
rect 19516 16996 19572 18508
rect 19180 16790 19236 16828
rect 19292 16994 19572 16996
rect 19292 16942 19518 16994
rect 19570 16942 19572 16994
rect 19292 16940 19572 16942
rect 19628 18228 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20300 18788 20356 18956
rect 20300 18732 20580 18788
rect 20076 18676 20132 18686
rect 19964 18452 20020 18462
rect 19964 18358 20020 18396
rect 20076 18340 20132 18620
rect 20188 18564 20244 18574
rect 20188 18470 20244 18508
rect 20412 18452 20468 18462
rect 20076 18284 20244 18340
rect 19628 16996 19684 18172
rect 19852 17780 19908 17790
rect 19852 17686 19908 17724
rect 20188 17444 20244 18284
rect 20188 17378 20244 17388
rect 20300 18338 20356 18350
rect 20300 18286 20302 18338
rect 20354 18286 20356 18338
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 17108 20356 18286
rect 20412 17890 20468 18396
rect 20524 18450 20580 18732
rect 20524 18398 20526 18450
rect 20578 18398 20580 18450
rect 20524 18386 20580 18398
rect 20636 18228 20692 22876
rect 20972 21700 21028 25452
rect 20748 21644 20972 21700
rect 20748 20804 20804 21644
rect 20972 21634 21028 21644
rect 21084 25396 21140 26348
rect 21196 26338 21252 26348
rect 21084 21252 21140 25340
rect 21196 25620 21252 25630
rect 21196 23938 21252 25564
rect 21308 25618 21364 26796
rect 21420 26068 21476 26078
rect 21420 25730 21476 26012
rect 21420 25678 21422 25730
rect 21474 25678 21476 25730
rect 21420 25666 21476 25678
rect 21308 25566 21310 25618
rect 21362 25566 21364 25618
rect 21308 25554 21364 25566
rect 21532 24612 21588 26852
rect 21868 26852 21924 28588
rect 21980 28578 22036 28588
rect 22652 28644 22708 29262
rect 22764 28754 22820 29932
rect 22876 29540 22932 29550
rect 22988 29540 23044 30158
rect 22932 29484 23044 29540
rect 22876 29426 22932 29484
rect 22876 29374 22878 29426
rect 22930 29374 22932 29426
rect 22876 29362 22932 29374
rect 22764 28702 22766 28754
rect 22818 28702 22820 28754
rect 22764 28690 22820 28702
rect 22876 29204 22932 29214
rect 22652 28578 22708 28588
rect 22652 27858 22708 27870
rect 22652 27806 22654 27858
rect 22706 27806 22708 27858
rect 21980 27748 22036 27758
rect 21980 27746 22260 27748
rect 21980 27694 21982 27746
rect 22034 27694 22260 27746
rect 21980 27692 22260 27694
rect 21980 27682 22036 27692
rect 22092 26962 22148 26974
rect 22092 26910 22094 26962
rect 22146 26910 22148 26962
rect 22092 26908 22148 26910
rect 21756 26292 21812 26302
rect 21756 26198 21812 26236
rect 21868 25506 21924 26796
rect 21868 25454 21870 25506
rect 21922 25454 21924 25506
rect 21868 25442 21924 25454
rect 21980 26852 22148 26908
rect 21532 24546 21588 24556
rect 21196 23886 21198 23938
rect 21250 23886 21252 23938
rect 21196 23874 21252 23886
rect 21532 23940 21588 23950
rect 21532 23846 21588 23884
rect 21420 23716 21476 23726
rect 21308 23714 21476 23716
rect 21308 23662 21422 23714
rect 21474 23662 21476 23714
rect 21308 23660 21476 23662
rect 21308 23268 21364 23660
rect 21420 23650 21476 23660
rect 21868 23716 21924 23726
rect 21868 23380 21924 23660
rect 21308 22932 21364 23212
rect 21308 22594 21364 22876
rect 21644 23324 21924 23380
rect 21532 22820 21588 22830
rect 21308 22542 21310 22594
rect 21362 22542 21364 22594
rect 21308 22530 21364 22542
rect 21420 22764 21532 22820
rect 21308 21476 21364 21486
rect 21308 21382 21364 21420
rect 21084 21186 21140 21196
rect 20860 21028 20916 21038
rect 21308 21028 21364 21038
rect 20860 21026 21364 21028
rect 20860 20974 20862 21026
rect 20914 20974 21310 21026
rect 21362 20974 21364 21026
rect 20860 20972 21364 20974
rect 20860 20962 20916 20972
rect 21308 20962 21364 20972
rect 21420 20916 21476 22764
rect 21532 22754 21588 22764
rect 21532 22594 21588 22606
rect 21532 22542 21534 22594
rect 21586 22542 21588 22594
rect 21532 22146 21588 22542
rect 21532 22094 21534 22146
rect 21586 22094 21588 22146
rect 21532 21588 21588 22094
rect 21644 21700 21700 23324
rect 21756 23154 21812 23166
rect 21756 23102 21758 23154
rect 21810 23102 21812 23154
rect 21756 23044 21812 23102
rect 21756 22978 21812 22988
rect 21980 22932 22036 26852
rect 22204 26628 22260 27692
rect 22652 26852 22708 27806
rect 22652 26786 22708 26796
rect 22204 26562 22260 26572
rect 22652 26404 22708 26414
rect 22540 26348 22652 26404
rect 22428 26068 22484 26078
rect 22428 25974 22484 26012
rect 22540 25844 22596 26348
rect 22652 26338 22708 26348
rect 22876 26290 22932 29148
rect 22988 27972 23044 27982
rect 22988 27858 23044 27916
rect 22988 27806 22990 27858
rect 23042 27806 23044 27858
rect 22988 27794 23044 27806
rect 23100 26908 23156 30828
rect 23212 29650 23268 31612
rect 23324 31666 23380 31678
rect 23324 31614 23326 31666
rect 23378 31614 23380 31666
rect 23324 30996 23380 31614
rect 23324 30930 23380 30940
rect 23212 29598 23214 29650
rect 23266 29598 23268 29650
rect 23212 29586 23268 29598
rect 23324 30772 23380 30782
rect 23324 30210 23380 30716
rect 23324 30158 23326 30210
rect 23378 30158 23380 30210
rect 23324 29316 23380 30158
rect 23324 29250 23380 29260
rect 23212 28868 23268 28878
rect 23212 28082 23268 28812
rect 23212 28030 23214 28082
rect 23266 28030 23268 28082
rect 23212 28018 23268 28030
rect 23324 28532 23380 28542
rect 23324 27858 23380 28476
rect 23324 27806 23326 27858
rect 23378 27806 23380 27858
rect 23324 27794 23380 27806
rect 23436 26908 23492 32284
rect 23548 32562 23604 32574
rect 23548 32510 23550 32562
rect 23602 32510 23604 32562
rect 23548 29204 23604 32510
rect 23660 31668 23716 33070
rect 23660 31602 23716 31612
rect 23772 33122 23940 33124
rect 23772 33070 23886 33122
rect 23938 33070 23940 33122
rect 23772 33068 23940 33070
rect 23660 31108 23716 31118
rect 23660 29650 23716 31052
rect 23660 29598 23662 29650
rect 23714 29598 23716 29650
rect 23660 29586 23716 29598
rect 23772 29538 23828 33068
rect 23884 33058 23940 33068
rect 23884 32788 23940 32798
rect 23996 32788 24052 33740
rect 24220 33236 24276 35252
rect 24668 35026 24724 35644
rect 25340 35634 25396 35644
rect 25452 35588 25508 36204
rect 26236 35698 26292 37212
rect 26236 35646 26238 35698
rect 26290 35646 26292 35698
rect 26236 35634 26292 35646
rect 26348 36372 26404 39004
rect 26572 38668 26628 39228
rect 26684 39060 26740 39070
rect 26684 38966 26740 39004
rect 26908 39060 26964 39070
rect 26908 38668 26964 39004
rect 27020 38836 27076 38846
rect 27020 38742 27076 38780
rect 27132 38668 27188 39452
rect 27356 39284 27412 39294
rect 27356 39058 27412 39228
rect 27356 39006 27358 39058
rect 27410 39006 27412 39058
rect 27356 38994 27412 39006
rect 27468 39172 27524 39182
rect 27468 39058 27524 39116
rect 27468 39006 27470 39058
rect 27522 39006 27524 39058
rect 27468 38994 27524 39006
rect 27580 39058 27636 40908
rect 27692 40898 27748 40908
rect 27804 39396 27860 42478
rect 28140 42532 28196 42542
rect 28140 42438 28196 42476
rect 28700 42530 28756 42542
rect 28700 42478 28702 42530
rect 28754 42478 28756 42530
rect 28700 42420 28756 42478
rect 28812 42532 28868 44044
rect 29484 44098 29540 44110
rect 29484 44046 29486 44098
rect 29538 44046 29540 44098
rect 29148 43764 29204 43774
rect 29148 43650 29204 43708
rect 29148 43598 29150 43650
rect 29202 43598 29204 43650
rect 28924 42532 28980 42542
rect 28812 42476 28924 42532
rect 29148 42532 29204 43598
rect 29484 43762 29540 44046
rect 29484 43710 29486 43762
rect 29538 43710 29540 43762
rect 29484 43652 29540 43710
rect 29596 44098 29652 44110
rect 29596 44046 29598 44098
rect 29650 44046 29652 44098
rect 29596 43764 29652 44046
rect 29932 43876 29988 44156
rect 30716 44210 30996 44212
rect 30716 44158 30942 44210
rect 30994 44158 30996 44210
rect 30716 44156 30996 44158
rect 29932 43820 30100 43876
rect 29596 43708 29988 43764
rect 29484 43586 29540 43596
rect 29596 43540 29652 43550
rect 29820 43540 29876 43550
rect 29652 43538 29876 43540
rect 29652 43486 29822 43538
rect 29874 43486 29876 43538
rect 29652 43484 29876 43486
rect 29596 43204 29652 43484
rect 29820 43474 29876 43484
rect 29484 43148 29652 43204
rect 29260 42868 29316 42878
rect 29260 42774 29316 42812
rect 29484 42754 29540 43148
rect 29484 42702 29486 42754
rect 29538 42702 29540 42754
rect 29484 42690 29540 42702
rect 29820 42756 29876 42766
rect 29596 42642 29652 42654
rect 29596 42590 29598 42642
rect 29650 42590 29652 42642
rect 29596 42532 29652 42590
rect 29148 42476 29652 42532
rect 28924 42466 28980 42476
rect 28028 41858 28084 41870
rect 28028 41806 28030 41858
rect 28082 41806 28084 41858
rect 28028 41188 28084 41806
rect 28028 40402 28084 41132
rect 28140 41300 28196 41310
rect 28140 41076 28196 41244
rect 28700 41188 28756 42364
rect 28700 41132 29092 41188
rect 28588 41076 28644 41086
rect 28140 41020 28308 41076
rect 28028 40350 28030 40402
rect 28082 40350 28084 40402
rect 27916 39620 27972 39630
rect 28028 39620 28084 40350
rect 27916 39618 28084 39620
rect 27916 39566 27918 39618
rect 27970 39566 28084 39618
rect 27916 39564 28084 39566
rect 28252 39618 28308 41020
rect 28588 41074 28868 41076
rect 28588 41022 28590 41074
rect 28642 41022 28868 41074
rect 28588 41020 28868 41022
rect 28588 41010 28644 41020
rect 28476 40964 28532 41002
rect 28476 40898 28532 40908
rect 28252 39566 28254 39618
rect 28306 39566 28308 39618
rect 27916 39554 27972 39564
rect 28252 39554 28308 39566
rect 28476 40740 28532 40750
rect 28476 40180 28532 40684
rect 28588 40626 28644 40638
rect 28588 40574 28590 40626
rect 28642 40574 28644 40626
rect 28588 40404 28644 40574
rect 28588 40338 28644 40348
rect 28588 40180 28644 40190
rect 28476 40178 28644 40180
rect 28476 40126 28590 40178
rect 28642 40126 28644 40178
rect 28476 40124 28644 40126
rect 27804 39340 27972 39396
rect 27580 39006 27582 39058
rect 27634 39006 27636 39058
rect 27580 38994 27636 39006
rect 27804 39060 27860 39070
rect 26572 38612 26740 38668
rect 26908 38612 27188 38668
rect 27244 38834 27300 38846
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 26684 38050 26740 38612
rect 26684 37998 26686 38050
rect 26738 37998 26740 38050
rect 26684 37716 26740 37998
rect 26796 38500 26852 38510
rect 26796 37940 26852 38444
rect 26796 37846 26852 37884
rect 26684 37660 26852 37716
rect 26348 35700 26404 36316
rect 26684 37378 26740 37390
rect 26684 37326 26686 37378
rect 26738 37326 26740 37378
rect 26684 36260 26740 37326
rect 26796 36484 26852 37660
rect 26908 36484 26964 36494
rect 26796 36482 26964 36484
rect 26796 36430 26910 36482
rect 26962 36430 26964 36482
rect 26796 36428 26964 36430
rect 26908 36418 26964 36428
rect 26908 36260 26964 36270
rect 26684 36258 26964 36260
rect 26684 36206 26910 36258
rect 26962 36206 26964 36258
rect 26684 36204 26964 36206
rect 26348 35644 26628 35700
rect 25900 35588 25956 35598
rect 25452 35522 25508 35532
rect 25676 35586 25956 35588
rect 25676 35534 25902 35586
rect 25954 35534 25956 35586
rect 25676 35532 25956 35534
rect 25676 35476 25732 35532
rect 25900 35522 25956 35532
rect 24668 34974 24670 35026
rect 24722 34974 24724 35026
rect 24668 34962 24724 34974
rect 25116 35364 25172 35374
rect 25116 34914 25172 35308
rect 25116 34862 25118 34914
rect 25170 34862 25172 34914
rect 25116 34850 25172 34862
rect 25340 34468 25396 34478
rect 25340 34354 25396 34412
rect 25340 34302 25342 34354
rect 25394 34302 25396 34354
rect 25340 34290 25396 34302
rect 24332 34242 24388 34254
rect 24332 34190 24334 34242
rect 24386 34190 24388 34242
rect 24332 33684 24388 34190
rect 24444 34244 24500 34254
rect 24444 34150 24500 34188
rect 25228 34244 25284 34254
rect 25228 34150 25284 34188
rect 25340 33908 25396 33918
rect 25564 33908 25620 33918
rect 25340 33814 25396 33852
rect 25452 33852 25564 33908
rect 24332 33618 24388 33628
rect 25452 33458 25508 33852
rect 25564 33842 25620 33852
rect 25676 33796 25732 35420
rect 26460 35476 26516 35486
rect 25788 34804 25844 34814
rect 25788 34802 26404 34804
rect 25788 34750 25790 34802
rect 25842 34750 26404 34802
rect 25788 34748 26404 34750
rect 25788 34738 25844 34748
rect 26348 34354 26404 34748
rect 26348 34302 26350 34354
rect 26402 34302 26404 34354
rect 26348 34290 26404 34302
rect 26460 34242 26516 35420
rect 26460 34190 26462 34242
rect 26514 34190 26516 34242
rect 26460 34178 26516 34190
rect 26012 34018 26068 34030
rect 26012 33966 26014 34018
rect 26066 33966 26068 34018
rect 25900 33908 25956 33918
rect 25900 33814 25956 33852
rect 25676 33730 25732 33740
rect 25452 33406 25454 33458
rect 25506 33406 25508 33458
rect 25452 33394 25508 33406
rect 26012 33460 26068 33966
rect 26012 33394 26068 33404
rect 26124 33684 26180 33694
rect 24780 33346 24836 33358
rect 24780 33294 24782 33346
rect 24834 33294 24836 33346
rect 24220 33234 24388 33236
rect 24220 33182 24222 33234
rect 24274 33182 24388 33234
rect 24220 33180 24388 33182
rect 24220 33170 24276 33180
rect 23884 32786 24052 32788
rect 23884 32734 23886 32786
rect 23938 32734 24052 32786
rect 23884 32732 24052 32734
rect 24108 33122 24164 33134
rect 24108 33070 24110 33122
rect 24162 33070 24164 33122
rect 23884 32722 23940 32732
rect 24108 32564 24164 33070
rect 24108 32498 24164 32508
rect 24220 32562 24276 32574
rect 24220 32510 24222 32562
rect 24274 32510 24276 32562
rect 24108 31668 24164 31678
rect 24220 31668 24276 32510
rect 24332 32452 24388 33180
rect 24556 32564 24612 32574
rect 24556 32470 24612 32508
rect 24444 32452 24500 32462
rect 24332 32396 24444 32452
rect 24444 32386 24500 32396
rect 24668 32338 24724 32350
rect 24668 32286 24670 32338
rect 24722 32286 24724 32338
rect 24164 31612 24276 31668
rect 24444 32116 24500 32126
rect 24108 31602 24164 31612
rect 23884 30210 23940 30222
rect 23884 30158 23886 30210
rect 23938 30158 23940 30210
rect 23884 29652 23940 30158
rect 24332 29764 24388 29774
rect 24332 29652 24388 29708
rect 23884 29596 24388 29652
rect 23772 29486 23774 29538
rect 23826 29486 23828 29538
rect 23772 29474 23828 29486
rect 23996 29426 24052 29438
rect 23996 29374 23998 29426
rect 24050 29374 24052 29426
rect 23660 29204 23716 29214
rect 23548 29202 23716 29204
rect 23548 29150 23662 29202
rect 23714 29150 23716 29202
rect 23548 29148 23716 29150
rect 23660 29138 23716 29148
rect 23996 28980 24052 29374
rect 23660 27860 23716 27870
rect 23660 27858 23828 27860
rect 23660 27806 23662 27858
rect 23714 27806 23828 27858
rect 23660 27804 23828 27806
rect 23660 27794 23716 27804
rect 23100 26852 23268 26908
rect 22988 26628 23044 26638
rect 22988 26514 23044 26572
rect 22988 26462 22990 26514
rect 23042 26462 23044 26514
rect 22988 26450 23044 26462
rect 23212 26516 23268 26852
rect 23212 26450 23268 26460
rect 23324 26852 23492 26908
rect 23660 27636 23716 27646
rect 22876 26238 22878 26290
rect 22930 26238 22932 26290
rect 22428 25788 22596 25844
rect 22652 26178 22708 26190
rect 22652 26126 22654 26178
rect 22706 26126 22708 26178
rect 22316 25172 22372 25182
rect 22204 25116 22316 25172
rect 22204 23940 22260 25116
rect 22316 25106 22372 25116
rect 22204 23874 22260 23884
rect 22316 24612 22372 24622
rect 22092 23714 22148 23726
rect 22092 23662 22094 23714
rect 22146 23662 22148 23714
rect 22092 23604 22148 23662
rect 22092 23538 22148 23548
rect 21868 22876 22036 22932
rect 21868 22596 21924 22876
rect 21756 22540 21924 22596
rect 21756 22148 21812 22540
rect 21980 22484 22036 22494
rect 21868 22372 21924 22382
rect 21980 22372 22036 22428
rect 21868 22370 22036 22372
rect 21868 22318 21870 22370
rect 21922 22318 22036 22370
rect 21868 22316 22036 22318
rect 22316 22370 22372 24556
rect 22428 23826 22484 25788
rect 22652 25620 22708 26126
rect 22652 25554 22708 25564
rect 22540 25394 22596 25406
rect 22540 25342 22542 25394
rect 22594 25342 22596 25394
rect 22540 24948 22596 25342
rect 22540 24882 22596 24892
rect 22652 25060 22708 25070
rect 22652 23940 22708 25004
rect 22876 24164 22932 26238
rect 23100 26290 23156 26302
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 23100 25284 23156 26238
rect 23100 25218 23156 25228
rect 23324 25060 23380 26852
rect 23324 24994 23380 25004
rect 23436 26516 23492 26526
rect 23324 24836 23380 24846
rect 23436 24836 23492 26460
rect 23660 26402 23716 27580
rect 23660 26350 23662 26402
rect 23714 26350 23716 26402
rect 23660 26338 23716 26350
rect 23772 26516 23828 27804
rect 23996 27858 24052 28924
rect 23996 27806 23998 27858
rect 24050 27806 24052 27858
rect 23996 27794 24052 27806
rect 24220 27186 24276 27198
rect 24220 27134 24222 27186
rect 24274 27134 24276 27186
rect 24108 26516 24164 26526
rect 23772 26514 24164 26516
rect 23772 26462 24110 26514
rect 24162 26462 24164 26514
rect 23772 26460 24164 26462
rect 23548 26292 23604 26302
rect 23548 26198 23604 26236
rect 23324 24834 23492 24836
rect 23324 24782 23326 24834
rect 23378 24782 23492 24834
rect 23324 24780 23492 24782
rect 23324 24770 23380 24780
rect 23660 24722 23716 24734
rect 23660 24670 23662 24722
rect 23714 24670 23716 24722
rect 23212 24500 23268 24510
rect 22876 24108 23044 24164
rect 22876 23940 22932 23950
rect 22652 23884 22820 23940
rect 22428 23774 22430 23826
rect 22482 23774 22484 23826
rect 22428 23762 22484 23774
rect 22540 23828 22596 23838
rect 22540 23826 22708 23828
rect 22540 23774 22542 23826
rect 22594 23774 22708 23826
rect 22540 23772 22708 23774
rect 22540 23762 22596 23772
rect 22540 23492 22596 23502
rect 22428 23380 22484 23390
rect 22428 22932 22484 23324
rect 22540 23378 22596 23436
rect 22540 23326 22542 23378
rect 22594 23326 22596 23378
rect 22540 23314 22596 23326
rect 22652 23154 22708 23772
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22540 22932 22596 22942
rect 22428 22930 22596 22932
rect 22428 22878 22542 22930
rect 22594 22878 22596 22930
rect 22428 22876 22596 22878
rect 22316 22318 22318 22370
rect 22370 22318 22372 22370
rect 21868 22306 21924 22316
rect 22316 22306 22372 22318
rect 21756 22092 21924 22148
rect 21644 21644 21812 21700
rect 21532 21532 21700 21588
rect 21532 20916 21588 20926
rect 21420 20914 21588 20916
rect 21420 20862 21534 20914
rect 21586 20862 21588 20914
rect 21420 20860 21588 20862
rect 21532 20850 21588 20860
rect 20748 20748 20916 20804
rect 20748 20578 20804 20590
rect 20748 20526 20750 20578
rect 20802 20526 20804 20578
rect 20748 20244 20804 20526
rect 20860 20468 20916 20748
rect 20860 20402 20916 20412
rect 21196 20692 21252 20702
rect 20748 20188 21140 20244
rect 21084 19908 21140 20188
rect 21196 20130 21252 20636
rect 21196 20078 21198 20130
rect 21250 20078 21252 20130
rect 21196 20066 21252 20078
rect 21644 19908 21700 21532
rect 21756 20804 21812 21644
rect 21868 20914 21924 22092
rect 21980 22146 22036 22158
rect 21980 22094 21982 22146
rect 22034 22094 22036 22146
rect 21980 22036 22036 22094
rect 22540 22148 22596 22876
rect 22652 22708 22708 23102
rect 22652 22642 22708 22652
rect 22540 22092 22708 22148
rect 21980 21980 22596 22036
rect 21868 20862 21870 20914
rect 21922 20862 21924 20914
rect 21868 20850 21924 20862
rect 21980 21812 22036 21822
rect 21756 20710 21812 20748
rect 21980 20802 22036 21756
rect 22428 21812 22484 21822
rect 21980 20750 21982 20802
rect 22034 20750 22036 20802
rect 21980 20738 22036 20750
rect 22092 21586 22148 21598
rect 22092 21534 22094 21586
rect 22146 21534 22148 21586
rect 22092 20132 22148 21534
rect 22092 20066 22148 20076
rect 21084 19852 21700 19908
rect 20748 19460 20804 19470
rect 20804 19404 20916 19460
rect 20748 19394 20804 19404
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 20412 17838 20414 17890
rect 20466 17838 20468 17890
rect 20412 17826 20468 17838
rect 20524 18172 20692 18228
rect 20524 17668 20580 18172
rect 20412 17612 20580 17668
rect 20636 17780 20692 17790
rect 20412 17220 20468 17612
rect 20524 17444 20580 17454
rect 20524 17350 20580 17388
rect 20412 17164 20580 17220
rect 20076 17052 20356 17108
rect 20524 17108 20580 17164
rect 19740 16996 19796 17006
rect 19628 16994 19796 16996
rect 19628 16942 19742 16994
rect 19794 16942 19796 16994
rect 19628 16940 19796 16942
rect 18956 16660 19012 16670
rect 18732 16146 18788 16156
rect 18844 16658 19012 16660
rect 18844 16606 18958 16658
rect 19010 16606 19012 16658
rect 18844 16604 19012 16606
rect 18284 16100 18340 16110
rect 18172 15876 18228 15886
rect 18060 15820 18172 15876
rect 18060 15538 18116 15820
rect 18172 15810 18228 15820
rect 18060 15486 18062 15538
rect 18114 15486 18116 15538
rect 18060 15474 18116 15486
rect 18172 15540 18228 15550
rect 18284 15540 18340 16044
rect 18172 15538 18340 15540
rect 18172 15486 18174 15538
rect 18226 15486 18340 15538
rect 18172 15484 18340 15486
rect 18732 15764 18788 15774
rect 18172 15474 18228 15484
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 15362 18004 15374
rect 18732 15314 18788 15708
rect 18732 15262 18734 15314
rect 18786 15262 18788 15314
rect 18732 15250 18788 15262
rect 18844 15316 18900 16604
rect 18956 16594 19012 16604
rect 18956 16100 19012 16138
rect 19012 16044 19124 16100
rect 18956 16034 19012 16044
rect 17500 15204 17556 15242
rect 17500 15138 17556 15148
rect 18396 15204 18452 15214
rect 18396 14642 18452 15148
rect 18396 14590 18398 14642
rect 18450 14590 18452 14642
rect 18396 14578 18452 14590
rect 16716 13746 16884 13748
rect 16716 13694 16718 13746
rect 16770 13694 16884 13746
rect 16716 13692 16884 13694
rect 16604 12404 16660 12414
rect 16604 12290 16660 12348
rect 16716 12404 16772 13692
rect 18396 13634 18452 13646
rect 18396 13582 18398 13634
rect 18450 13582 18452 13634
rect 18284 13524 18340 13534
rect 17724 13522 18340 13524
rect 17724 13470 18286 13522
rect 18338 13470 18340 13522
rect 17724 13468 18340 13470
rect 17052 12850 17108 12862
rect 17052 12798 17054 12850
rect 17106 12798 17108 12850
rect 17052 12404 17108 12798
rect 16716 12402 16884 12404
rect 16716 12350 16718 12402
rect 16770 12350 16884 12402
rect 16716 12348 16884 12350
rect 16716 12338 16772 12348
rect 16604 12238 16606 12290
rect 16658 12238 16660 12290
rect 16604 12226 16660 12238
rect 16492 12012 16772 12068
rect 16380 11900 16660 11956
rect 16268 11564 16548 11620
rect 15932 11452 16212 11508
rect 15932 11396 15988 11452
rect 16156 11396 16212 11452
rect 16268 11396 16324 11406
rect 16156 11394 16324 11396
rect 16156 11342 16270 11394
rect 16322 11342 16324 11394
rect 16156 11340 16324 11342
rect 15932 11330 15988 11340
rect 16268 11330 16324 11340
rect 16044 11172 16100 11182
rect 16044 11078 16100 11116
rect 16156 11170 16212 11182
rect 16156 11118 16158 11170
rect 16210 11118 16212 11170
rect 15820 10892 15988 10948
rect 15484 10670 15486 10722
rect 15538 10670 15540 10722
rect 15484 10658 15540 10670
rect 15372 10612 15428 10622
rect 15260 10556 15372 10612
rect 15372 10546 15428 10556
rect 15820 10612 15876 10622
rect 15596 10498 15652 10510
rect 15596 10446 15598 10498
rect 15650 10446 15652 10498
rect 15148 10386 15316 10388
rect 15148 10334 15150 10386
rect 15202 10334 15316 10386
rect 15148 10332 15316 10334
rect 15148 10322 15204 10332
rect 14476 9886 14478 9938
rect 14530 9886 14532 9938
rect 13468 9828 13524 9838
rect 13468 9714 13524 9772
rect 13468 9662 13470 9714
rect 13522 9662 13524 9714
rect 13468 9650 13524 9662
rect 13804 9714 13860 9726
rect 13804 9662 13806 9714
rect 13858 9662 13860 9714
rect 13804 9156 13860 9662
rect 14140 9268 14196 9278
rect 13804 9090 13860 9100
rect 14028 9154 14084 9166
rect 14028 9102 14030 9154
rect 14082 9102 14084 9154
rect 13692 9044 13748 9054
rect 13692 8950 13748 8988
rect 13244 8932 13300 8942
rect 13132 8876 13244 8932
rect 12908 8148 12964 8158
rect 12908 8054 12964 8092
rect 13132 7474 13188 8876
rect 13244 8866 13300 8876
rect 13804 8036 13860 8046
rect 13804 7942 13860 7980
rect 13916 7588 13972 7598
rect 14028 7588 14084 9102
rect 14140 8148 14196 9212
rect 14140 8054 14196 8092
rect 14364 9154 14420 9166
rect 14364 9102 14366 9154
rect 14418 9102 14420 9154
rect 13916 7586 14084 7588
rect 13916 7534 13918 7586
rect 13970 7534 14084 7586
rect 13916 7532 14084 7534
rect 13916 7522 13972 7532
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 12908 7028 12964 7038
rect 12908 6914 12964 6972
rect 12908 6862 12910 6914
rect 12962 6862 12964 6914
rect 12908 6850 12964 6862
rect 13132 6804 13188 7422
rect 13132 6738 13188 6748
rect 14028 6804 14084 6814
rect 13244 6692 13300 6702
rect 12796 5954 12852 5964
rect 13020 6580 13076 6590
rect 12908 5908 12964 5918
rect 12572 5460 12628 5470
rect 11564 3378 11620 3388
rect 12124 4452 12180 4462
rect 12124 800 12180 4396
rect 12572 3666 12628 5404
rect 12908 5234 12964 5852
rect 12908 5182 12910 5234
rect 12962 5182 12964 5234
rect 12908 5170 12964 5182
rect 12908 4228 12964 4238
rect 13020 4228 13076 6524
rect 12908 4226 13076 4228
rect 12908 4174 12910 4226
rect 12962 4174 13076 4226
rect 12908 4172 13076 4174
rect 13132 5794 13188 5806
rect 13132 5742 13134 5794
rect 13186 5742 13188 5794
rect 13132 5124 13188 5742
rect 12908 4162 12964 4172
rect 12572 3614 12574 3666
rect 12626 3614 12628 3666
rect 12572 3602 12628 3614
rect 13132 3554 13188 5068
rect 13244 4338 13300 6636
rect 13580 6466 13636 6478
rect 13580 6414 13582 6466
rect 13634 6414 13636 6466
rect 13580 6132 13636 6414
rect 13916 6468 13972 6478
rect 13916 6374 13972 6412
rect 13580 6066 13636 6076
rect 13916 4564 13972 4574
rect 13580 4452 13636 4462
rect 13580 4358 13636 4396
rect 13244 4286 13246 4338
rect 13298 4286 13300 4338
rect 13244 4274 13300 4286
rect 13356 4228 13412 4238
rect 13356 4134 13412 4172
rect 13916 3666 13972 4508
rect 14028 4338 14084 6748
rect 14364 6692 14420 9102
rect 14476 8820 14532 9886
rect 14812 9826 14868 9838
rect 14812 9774 14814 9826
rect 14866 9774 14868 9826
rect 14700 9268 14756 9278
rect 14700 9174 14756 9212
rect 14476 8754 14532 8764
rect 14588 8932 14644 8942
rect 14588 8428 14644 8876
rect 14812 8428 14868 9774
rect 15148 9156 15204 9166
rect 15148 9062 15204 9100
rect 15260 9044 15316 10332
rect 15596 9938 15652 10446
rect 15596 9886 15598 9938
rect 15650 9886 15652 9938
rect 15596 9874 15652 9886
rect 15708 9154 15764 9166
rect 15708 9102 15710 9154
rect 15762 9102 15764 9154
rect 15484 9044 15540 9054
rect 15260 9042 15540 9044
rect 15260 8990 15486 9042
rect 15538 8990 15540 9042
rect 15260 8988 15540 8990
rect 15484 8978 15540 8988
rect 15708 9042 15764 9102
rect 15708 8990 15710 9042
rect 15762 8990 15764 9042
rect 15708 8978 15764 8990
rect 15260 8820 15316 8830
rect 15260 8818 15540 8820
rect 15260 8766 15262 8818
rect 15314 8766 15540 8818
rect 15260 8764 15540 8766
rect 15260 8754 15316 8764
rect 15484 8596 15540 8764
rect 15820 8596 15876 10556
rect 15484 8540 15876 8596
rect 14588 8372 14868 8428
rect 14812 8278 14868 8316
rect 14364 6626 14420 6636
rect 15148 7028 15204 7038
rect 14252 6580 14308 6590
rect 14252 6486 14308 6524
rect 14476 6468 14532 6478
rect 14476 6374 14532 6412
rect 14588 6466 14644 6478
rect 14588 6414 14590 6466
rect 14642 6414 14644 6466
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 14588 3780 14644 6414
rect 14700 6466 14756 6478
rect 14700 6414 14702 6466
rect 14754 6414 14756 6466
rect 14700 5460 14756 6414
rect 14812 6468 14868 6478
rect 14812 6374 14868 6412
rect 15148 5796 15204 6972
rect 15596 6804 15652 6814
rect 15596 6710 15652 6748
rect 15372 6690 15428 6702
rect 15372 6638 15374 6690
rect 15426 6638 15428 6690
rect 15260 6468 15316 6478
rect 15260 6130 15316 6412
rect 15260 6078 15262 6130
rect 15314 6078 15316 6130
rect 15260 6066 15316 6078
rect 15372 6132 15428 6638
rect 15708 6580 15764 6590
rect 15708 6486 15764 6524
rect 15484 6466 15540 6478
rect 15484 6414 15486 6466
rect 15538 6414 15540 6466
rect 15484 6356 15540 6414
rect 15820 6468 15876 6478
rect 15820 6374 15876 6412
rect 15484 6132 15540 6300
rect 15596 6132 15652 6142
rect 15484 6130 15652 6132
rect 15484 6078 15598 6130
rect 15650 6078 15652 6130
rect 15484 6076 15652 6078
rect 15372 6038 15428 6076
rect 15596 6066 15652 6076
rect 15820 6020 15876 6030
rect 15820 5926 15876 5964
rect 15372 5796 15428 5806
rect 15148 5794 15428 5796
rect 15148 5742 15374 5794
rect 15426 5742 15428 5794
rect 15148 5740 15428 5742
rect 15372 5730 15428 5740
rect 14700 5394 14756 5404
rect 14700 5236 14756 5246
rect 14700 4450 14756 5180
rect 15932 5122 15988 10892
rect 16044 10724 16100 10734
rect 16156 10724 16212 11118
rect 16044 10722 16212 10724
rect 16044 10670 16046 10722
rect 16098 10670 16212 10722
rect 16044 10668 16212 10670
rect 16044 10658 16100 10668
rect 16044 9268 16100 9278
rect 16492 9268 16548 11564
rect 16604 10612 16660 11900
rect 16604 10546 16660 10556
rect 16044 9266 16548 9268
rect 16044 9214 16046 9266
rect 16098 9214 16548 9266
rect 16044 9212 16548 9214
rect 16604 9604 16660 9614
rect 16604 9266 16660 9548
rect 16604 9214 16606 9266
rect 16658 9214 16660 9266
rect 16044 9202 16100 9212
rect 16156 8932 16212 8942
rect 16156 8838 16212 8876
rect 16492 8932 16548 8942
rect 16380 8372 16436 8382
rect 16380 8036 16436 8316
rect 16044 7362 16100 7374
rect 16044 7310 16046 7362
rect 16098 7310 16100 7362
rect 16044 6804 16100 7310
rect 16044 6738 16100 6748
rect 16380 6690 16436 7980
rect 16492 7362 16548 8876
rect 16604 7924 16660 9214
rect 16716 9156 16772 12012
rect 16828 11956 16884 12348
rect 17052 12338 17108 12348
rect 16940 12180 16996 12190
rect 17388 12180 17444 12190
rect 16940 12178 17444 12180
rect 16940 12126 16942 12178
rect 16994 12126 17390 12178
rect 17442 12126 17444 12178
rect 16940 12124 17444 12126
rect 16940 12114 16996 12124
rect 17388 12114 17444 12124
rect 17724 12178 17780 13468
rect 18284 13458 18340 13468
rect 18396 13076 18452 13582
rect 18396 13010 18452 13020
rect 18172 12852 18228 12862
rect 17836 12404 17892 12414
rect 17836 12310 17892 12348
rect 18172 12402 18228 12796
rect 18172 12350 18174 12402
rect 18226 12350 18228 12402
rect 17724 12126 17726 12178
rect 17778 12126 17780 12178
rect 17724 12114 17780 12126
rect 18060 12180 18116 12190
rect 18172 12180 18228 12350
rect 18732 12740 18788 12750
rect 18060 12178 18228 12180
rect 18060 12126 18062 12178
rect 18114 12126 18228 12178
rect 18060 12124 18228 12126
rect 18396 12290 18452 12302
rect 18396 12238 18398 12290
rect 18450 12238 18452 12290
rect 18060 12114 18116 12124
rect 16828 11900 17220 11956
rect 17164 11506 17220 11900
rect 18396 11844 18452 12238
rect 18508 12180 18564 12190
rect 18508 12178 18676 12180
rect 18508 12126 18510 12178
rect 18562 12126 18676 12178
rect 18508 12124 18676 12126
rect 18508 12114 18564 12124
rect 18396 11778 18452 11788
rect 17164 11454 17166 11506
rect 17218 11454 17220 11506
rect 17164 11442 17220 11454
rect 18396 11508 18452 11518
rect 18396 11394 18452 11452
rect 18396 11342 18398 11394
rect 18450 11342 18452 11394
rect 18396 11330 18452 11342
rect 18620 11396 18676 12124
rect 18732 11618 18788 12684
rect 18844 12292 18900 15260
rect 18956 15874 19012 15886
rect 18956 15822 18958 15874
rect 19010 15822 19012 15874
rect 18956 15148 19012 15822
rect 19068 15540 19124 16044
rect 19180 16098 19236 16110
rect 19180 16046 19182 16098
rect 19234 16046 19236 16098
rect 19180 15764 19236 16046
rect 19180 15698 19236 15708
rect 19180 15540 19236 15550
rect 19068 15538 19236 15540
rect 19068 15486 19182 15538
rect 19234 15486 19236 15538
rect 19068 15484 19236 15486
rect 19180 15474 19236 15484
rect 19292 15538 19348 16940
rect 19516 16930 19572 16940
rect 19740 16930 19796 16940
rect 19964 16772 20020 16782
rect 19964 16678 20020 16716
rect 19292 15486 19294 15538
rect 19346 15486 19348 15538
rect 19292 15474 19348 15486
rect 19404 16212 19460 16222
rect 19404 15538 19460 16156
rect 20076 15876 20132 17052
rect 20524 17042 20580 17052
rect 20412 16996 20468 17006
rect 20412 16884 20468 16940
rect 20412 16828 20580 16884
rect 20300 16660 20356 16670
rect 20300 15988 20356 16604
rect 20300 15894 20356 15932
rect 20076 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 15820
rect 19404 15486 19406 15538
rect 19458 15486 19460 15538
rect 19404 15474 19460 15486
rect 19964 15484 20244 15540
rect 20524 15540 20580 16828
rect 19516 15316 19572 15326
rect 19740 15316 19796 15326
rect 19572 15314 19796 15316
rect 19572 15262 19742 15314
rect 19794 15262 19796 15314
rect 19572 15260 19796 15262
rect 19516 15250 19572 15260
rect 19740 15250 19796 15260
rect 19964 15314 20020 15484
rect 19964 15262 19966 15314
rect 20018 15262 20020 15314
rect 19964 15250 20020 15262
rect 20300 15204 20356 15242
rect 18956 15092 19124 15148
rect 20300 15138 20356 15148
rect 18844 12290 19012 12292
rect 18844 12238 18846 12290
rect 18898 12238 19012 12290
rect 18844 12236 19012 12238
rect 18844 12226 18900 12236
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11554 18788 11566
rect 18620 11340 18900 11396
rect 17388 11172 17444 11182
rect 17388 10834 17444 11116
rect 17388 10782 17390 10834
rect 17442 10782 17444 10834
rect 17388 10770 17444 10782
rect 18620 11170 18676 11182
rect 18620 11118 18622 11170
rect 18674 11118 18676 11170
rect 18620 10836 18676 11118
rect 18844 11172 18900 11340
rect 18956 11284 19012 12236
rect 19068 12178 19124 15092
rect 20188 15090 20244 15102
rect 20188 15038 20190 15090
rect 20242 15038 20244 15090
rect 20188 14980 20244 15038
rect 20524 14980 20580 15484
rect 20636 15148 20692 17724
rect 20748 17778 20804 17790
rect 20748 17726 20750 17778
rect 20802 17726 20804 17778
rect 20748 16772 20804 17726
rect 20748 16678 20804 16716
rect 20748 16212 20804 16222
rect 20860 16212 20916 19404
rect 20972 19124 21028 19134
rect 20972 16436 21028 19068
rect 21084 17892 21140 19852
rect 21532 19460 21588 19470
rect 21532 19346 21588 19404
rect 21532 19294 21534 19346
rect 21586 19294 21588 19346
rect 21532 19282 21588 19294
rect 22428 19348 22484 21756
rect 22540 21586 22596 21980
rect 22652 21924 22708 22092
rect 22652 21858 22708 21868
rect 22540 21534 22542 21586
rect 22594 21534 22596 21586
rect 22540 20802 22596 21534
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 22540 20738 22596 20750
rect 22764 20804 22820 23884
rect 22876 21812 22932 23884
rect 22988 23716 23044 24108
rect 22988 23622 23044 23660
rect 22988 23380 23044 23390
rect 22988 23266 23044 23324
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22988 23202 23044 23214
rect 23100 23268 23156 23278
rect 23100 23174 23156 23212
rect 23100 22930 23156 22942
rect 23100 22878 23102 22930
rect 23154 22878 23156 22930
rect 23100 22820 23156 22878
rect 23100 22754 23156 22764
rect 23100 22484 23156 22494
rect 23212 22484 23268 24444
rect 23548 24388 23604 24398
rect 23548 23940 23604 24332
rect 23100 22482 23268 22484
rect 23100 22430 23102 22482
rect 23154 22430 23268 22482
rect 23100 22428 23268 22430
rect 23324 23938 23604 23940
rect 23324 23886 23550 23938
rect 23602 23886 23604 23938
rect 23324 23884 23604 23886
rect 23100 22418 23156 22428
rect 22876 21746 22932 21756
rect 23212 21812 23268 21822
rect 23212 21718 23268 21756
rect 22988 21700 23044 21710
rect 22876 21588 22932 21598
rect 22876 21494 22932 21532
rect 22764 20748 22932 20804
rect 22764 20580 22820 20590
rect 22764 20486 22820 20524
rect 22876 20020 22932 20748
rect 22988 20244 23044 21644
rect 23100 21476 23156 21486
rect 23100 21382 23156 21420
rect 23324 21252 23380 23884
rect 23548 23874 23604 23884
rect 22988 20178 23044 20188
rect 23100 21196 23380 21252
rect 23436 23604 23492 23614
rect 23660 23604 23716 24670
rect 23492 23548 23716 23604
rect 22764 19964 22932 20020
rect 22428 19346 22596 19348
rect 22428 19294 22430 19346
rect 22482 19294 22596 19346
rect 22428 19292 22596 19294
rect 22428 19282 22484 19292
rect 21980 19234 22036 19246
rect 21980 19182 21982 19234
rect 22034 19182 22036 19234
rect 21420 19012 21476 19022
rect 21420 18918 21476 18956
rect 21980 19012 22036 19182
rect 21980 18946 22036 18956
rect 21308 18452 21364 18462
rect 21532 18452 21588 18462
rect 21308 18450 21588 18452
rect 21308 18398 21310 18450
rect 21362 18398 21534 18450
rect 21586 18398 21588 18450
rect 21308 18396 21588 18398
rect 21308 18386 21364 18396
rect 21532 18116 21588 18396
rect 21756 18452 21812 18462
rect 21756 18358 21812 18396
rect 22092 18450 22148 18462
rect 22092 18398 22094 18450
rect 22146 18398 22148 18450
rect 21644 18340 21700 18350
rect 21644 18246 21700 18284
rect 21084 17836 21364 17892
rect 20972 16380 21252 16436
rect 21196 16322 21252 16380
rect 21196 16270 21198 16322
rect 21250 16270 21252 16322
rect 21196 16258 21252 16270
rect 20748 16210 21140 16212
rect 20748 16158 20750 16210
rect 20802 16158 21140 16210
rect 20748 16156 21140 16158
rect 20748 16146 20804 16156
rect 20860 15428 20916 15438
rect 20636 15092 20804 15148
rect 20188 14924 20580 14980
rect 20076 14756 20132 14766
rect 20132 14700 20244 14756
rect 20076 14690 20132 14700
rect 19180 14530 19236 14542
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 13748 19236 14478
rect 19852 14420 19908 14430
rect 20076 14420 20132 14430
rect 19852 14418 20076 14420
rect 19852 14366 19854 14418
rect 19906 14366 20076 14418
rect 19852 14364 20076 14366
rect 19852 14354 19908 14364
rect 20076 14326 20132 14364
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19180 13682 19236 13692
rect 20076 13636 20132 13646
rect 20188 13636 20244 14700
rect 20076 13634 20244 13636
rect 20076 13582 20078 13634
rect 20130 13582 20244 13634
rect 20076 13580 20244 13582
rect 20076 13570 20132 13580
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 11506 19124 12126
rect 19180 13076 19236 13086
rect 19180 12180 19236 13020
rect 19516 12852 19572 12862
rect 19516 12758 19572 12796
rect 19628 12738 19684 12750
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19628 12628 19684 12686
rect 19852 12740 19908 12778
rect 19852 12674 19908 12684
rect 19628 12562 19684 12572
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20188 12516 20244 13580
rect 20188 12450 20244 12460
rect 20524 14642 20580 14924
rect 20524 14590 20526 14642
rect 20578 14590 20580 14642
rect 19292 12292 19348 12302
rect 20412 12292 20468 12302
rect 19292 12198 19348 12236
rect 20300 12290 20468 12292
rect 20300 12238 20414 12290
rect 20466 12238 20468 12290
rect 20300 12236 20468 12238
rect 19180 12114 19236 12124
rect 20076 12180 20132 12190
rect 20076 12086 20132 12124
rect 20300 11844 20356 12236
rect 20412 12226 20468 12236
rect 19068 11454 19070 11506
rect 19122 11454 19124 11506
rect 19068 11442 19124 11454
rect 20188 11508 20244 11518
rect 20188 11414 20244 11452
rect 19292 11394 19348 11406
rect 19292 11342 19294 11394
rect 19346 11342 19348 11394
rect 19292 11284 19348 11342
rect 20300 11394 20356 11788
rect 20300 11342 20302 11394
rect 20354 11342 20356 11394
rect 20300 11330 20356 11342
rect 18956 11228 19348 11284
rect 19964 11282 20020 11294
rect 19964 11230 19966 11282
rect 20018 11230 20020 11282
rect 19628 11172 19684 11182
rect 19964 11172 20020 11230
rect 18844 11170 20020 11172
rect 18844 11118 19630 11170
rect 19682 11118 20020 11170
rect 18844 11116 20020 11118
rect 19628 11106 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 18620 10780 19124 10836
rect 19068 10722 19124 10780
rect 19068 10670 19070 10722
rect 19122 10670 19124 10722
rect 19068 10658 19124 10670
rect 20524 10724 20580 14590
rect 20748 12740 20804 15092
rect 20860 14532 20916 15372
rect 21084 15314 21140 16156
rect 21084 15262 21086 15314
rect 21138 15262 21140 15314
rect 21084 15250 21140 15262
rect 21308 15148 21364 17836
rect 21532 17444 21588 18060
rect 22092 17780 22148 18398
rect 22316 18452 22372 18462
rect 22204 17780 22260 17790
rect 22092 17778 22260 17780
rect 22092 17726 22206 17778
rect 22258 17726 22260 17778
rect 22092 17724 22260 17726
rect 22204 17714 22260 17724
rect 22316 17666 22372 18396
rect 22428 18450 22484 18462
rect 22428 18398 22430 18450
rect 22482 18398 22484 18450
rect 22428 18228 22484 18398
rect 22428 18162 22484 18172
rect 22540 18004 22596 19292
rect 22540 17938 22596 17948
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 22316 17602 22372 17614
rect 22764 17666 22820 19964
rect 23100 19346 23156 21196
rect 23436 21140 23492 23548
rect 23772 23380 23828 26460
rect 24108 26450 24164 26460
rect 24220 26292 24276 27134
rect 23548 23324 23828 23380
rect 23884 26236 24276 26292
rect 23548 22932 23604 23324
rect 23660 23156 23716 23166
rect 23660 23062 23716 23100
rect 23660 22932 23716 22942
rect 23548 22876 23660 22932
rect 23660 22866 23716 22876
rect 23772 22930 23828 22942
rect 23772 22878 23774 22930
rect 23826 22878 23828 22930
rect 23772 21476 23828 22878
rect 23884 22596 23940 26236
rect 24108 25284 24164 25294
rect 23996 24948 24052 24958
rect 23996 24854 24052 24892
rect 24108 24834 24164 25228
rect 24108 24782 24110 24834
rect 24162 24782 24164 24834
rect 24108 24770 24164 24782
rect 24332 23380 24388 29596
rect 24444 29428 24500 32060
rect 24556 32004 24612 32014
rect 24556 30210 24612 31948
rect 24668 31668 24724 32286
rect 24780 31892 24836 33294
rect 25452 33124 25508 33134
rect 25228 32676 25284 32686
rect 25284 32620 25396 32676
rect 25228 32610 25284 32620
rect 24780 31826 24836 31836
rect 24668 31612 24948 31668
rect 24668 31108 24724 31118
rect 24668 30882 24724 31052
rect 24892 30996 24948 31612
rect 25228 30996 25284 31006
rect 24892 30994 25284 30996
rect 24892 30942 25230 30994
rect 25282 30942 25284 30994
rect 24892 30940 25284 30942
rect 25228 30930 25284 30940
rect 24668 30830 24670 30882
rect 24722 30830 24724 30882
rect 24668 30818 24724 30830
rect 24556 30158 24558 30210
rect 24610 30158 24612 30210
rect 24556 30146 24612 30158
rect 24668 30212 24724 30222
rect 24556 29652 24612 29662
rect 24556 29558 24612 29596
rect 24668 29650 24724 30156
rect 25340 30212 25396 32620
rect 25452 32562 25508 33068
rect 25452 32510 25454 32562
rect 25506 32510 25508 32562
rect 25452 32116 25508 32510
rect 25900 32452 25956 32462
rect 25452 32050 25508 32060
rect 25788 32450 25956 32452
rect 25788 32398 25902 32450
rect 25954 32398 25956 32450
rect 25788 32396 25956 32398
rect 24892 30100 24948 30110
rect 24892 30006 24948 30044
rect 25228 30098 25284 30110
rect 25228 30046 25230 30098
rect 25282 30046 25284 30098
rect 24668 29598 24670 29650
rect 24722 29598 24724 29650
rect 24444 29334 24500 29372
rect 24556 28532 24612 28542
rect 24556 28082 24612 28476
rect 24556 28030 24558 28082
rect 24610 28030 24612 28082
rect 24556 28018 24612 28030
rect 24668 28082 24724 29598
rect 25228 29652 25284 30046
rect 25340 29876 25396 30156
rect 25564 31892 25620 31902
rect 25340 29810 25396 29820
rect 25452 30098 25508 30110
rect 25452 30046 25454 30098
rect 25506 30046 25508 30098
rect 25228 29586 25284 29596
rect 25452 28868 25508 30046
rect 25452 28774 25508 28812
rect 25564 29314 25620 31836
rect 25676 29988 25732 29998
rect 25676 29894 25732 29932
rect 25564 29262 25566 29314
rect 25618 29262 25620 29314
rect 25564 29204 25620 29262
rect 24892 28756 24948 28766
rect 24668 28030 24670 28082
rect 24722 28030 24724 28082
rect 24668 28018 24724 28030
rect 24780 28700 24892 28756
rect 24444 27860 24500 27870
rect 24444 27858 24612 27860
rect 24444 27806 24446 27858
rect 24498 27806 24612 27858
rect 24444 27804 24612 27806
rect 24444 27794 24500 27804
rect 24556 27412 24612 27804
rect 24668 27412 24724 27422
rect 24556 27356 24668 27412
rect 24556 27188 24612 27198
rect 24556 25396 24612 27132
rect 24668 26516 24724 27356
rect 24780 27074 24836 28700
rect 24892 28662 24948 28700
rect 25340 28756 25396 28766
rect 25340 28662 25396 28700
rect 25564 28644 25620 29148
rect 25788 29092 25844 32396
rect 25900 32386 25956 32396
rect 26124 30772 26180 33628
rect 26572 32788 26628 35644
rect 26684 35698 26740 36204
rect 26908 36194 26964 36204
rect 26684 35646 26686 35698
rect 26738 35646 26740 35698
rect 26684 35634 26740 35646
rect 27020 35700 27076 38612
rect 27244 38274 27300 38782
rect 27580 38724 27636 38734
rect 27244 38222 27246 38274
rect 27298 38222 27300 38274
rect 27244 38210 27300 38222
rect 27356 38612 27636 38668
rect 27356 38164 27412 38612
rect 27356 38162 27636 38164
rect 27356 38110 27358 38162
rect 27410 38110 27636 38162
rect 27356 38108 27636 38110
rect 27356 38098 27412 38108
rect 27244 37940 27300 37950
rect 27244 36594 27300 37884
rect 27244 36542 27246 36594
rect 27298 36542 27300 36594
rect 27244 36530 27300 36542
rect 27132 36036 27188 36046
rect 27132 35922 27188 35980
rect 27132 35870 27134 35922
rect 27186 35870 27188 35922
rect 27132 35858 27188 35870
rect 27244 35812 27300 35822
rect 27020 35644 27188 35700
rect 26572 32722 26628 32732
rect 26908 34692 26964 34702
rect 26908 34354 26964 34636
rect 26908 34302 26910 34354
rect 26962 34302 26964 34354
rect 26348 32676 26404 32686
rect 26348 32582 26404 32620
rect 26572 32562 26628 32574
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 26572 32004 26628 32510
rect 26908 32564 26964 34302
rect 26908 32498 26964 32508
rect 26572 31938 26628 31948
rect 27020 31780 27076 31790
rect 27020 31668 27076 31724
rect 26908 31666 27076 31668
rect 26908 31614 27022 31666
rect 27074 31614 27076 31666
rect 26908 31612 27076 31614
rect 26908 31332 26964 31612
rect 27020 31602 27076 31612
rect 27132 31332 27188 35644
rect 27244 33012 27300 35756
rect 27468 35698 27524 35710
rect 27468 35646 27470 35698
rect 27522 35646 27524 35698
rect 27468 35364 27524 35646
rect 27468 35298 27524 35308
rect 27356 34692 27412 34702
rect 27356 34354 27412 34636
rect 27356 34302 27358 34354
rect 27410 34302 27412 34354
rect 27356 34290 27412 34302
rect 27580 33460 27636 38108
rect 27692 38052 27748 38062
rect 27692 37604 27748 37996
rect 27692 37538 27748 37548
rect 27804 37490 27860 39004
rect 27804 37438 27806 37490
rect 27858 37438 27860 37490
rect 27804 37426 27860 37438
rect 27916 38948 27972 39340
rect 27916 35252 27972 38892
rect 28028 39172 28084 39182
rect 28028 38946 28084 39116
rect 28476 39060 28532 40124
rect 28588 40114 28644 40124
rect 28700 40180 28756 40190
rect 28700 40086 28756 40124
rect 28476 38994 28532 39004
rect 28588 39394 28644 39406
rect 28588 39342 28590 39394
rect 28642 39342 28644 39394
rect 28028 38894 28030 38946
rect 28082 38894 28084 38946
rect 28028 38882 28084 38894
rect 28588 38948 28644 39342
rect 28588 38882 28644 38892
rect 28364 38834 28420 38846
rect 28364 38782 28366 38834
rect 28418 38782 28420 38834
rect 28028 38724 28084 38734
rect 28028 38050 28084 38668
rect 28028 37998 28030 38050
rect 28082 37998 28084 38050
rect 28028 37986 28084 37998
rect 28140 38610 28196 38622
rect 28140 38558 28142 38610
rect 28194 38558 28196 38610
rect 28140 37828 28196 38558
rect 28364 38052 28420 38782
rect 28700 38834 28756 38846
rect 28700 38782 28702 38834
rect 28754 38782 28756 38834
rect 28700 38724 28756 38782
rect 28700 38658 28756 38668
rect 28364 37986 28420 37996
rect 28812 38164 28868 41020
rect 28924 40178 28980 40190
rect 28924 40126 28926 40178
rect 28978 40126 28980 40178
rect 28924 40068 28980 40126
rect 28924 40002 28980 40012
rect 28924 39508 28980 39518
rect 28924 38834 28980 39452
rect 28924 38782 28926 38834
rect 28978 38782 28980 38834
rect 28924 38770 28980 38782
rect 28252 37940 28308 37950
rect 28252 37846 28308 37884
rect 28140 37734 28196 37772
rect 28364 37828 28420 37838
rect 28812 37828 28868 38108
rect 28364 37826 28868 37828
rect 28364 37774 28366 37826
rect 28418 37774 28868 37826
rect 28364 37772 28868 37774
rect 28140 37604 28196 37614
rect 28140 37266 28196 37548
rect 28140 37214 28142 37266
rect 28194 37214 28196 37266
rect 28140 37202 28196 37214
rect 28252 36260 28308 36270
rect 28252 35810 28308 36204
rect 28252 35758 28254 35810
rect 28306 35758 28308 35810
rect 28252 35746 28308 35758
rect 28364 36148 28420 37772
rect 27804 35196 27972 35252
rect 27804 34692 27860 35196
rect 27916 35028 27972 35038
rect 28364 35028 28420 36092
rect 27916 35026 28420 35028
rect 27916 34974 27918 35026
rect 27970 34974 28420 35026
rect 27916 34972 28420 34974
rect 28700 36258 28756 36270
rect 28700 36206 28702 36258
rect 28754 36206 28756 36258
rect 27916 34962 27972 34972
rect 28588 34692 28644 34702
rect 27804 34636 28084 34692
rect 27804 34468 27860 34478
rect 27804 34354 27860 34412
rect 27804 34302 27806 34354
rect 27858 34302 27860 34354
rect 27804 34290 27860 34302
rect 27580 33458 27972 33460
rect 27580 33406 27582 33458
rect 27634 33406 27972 33458
rect 27580 33404 27972 33406
rect 27580 33394 27636 33404
rect 27916 33346 27972 33404
rect 27916 33294 27918 33346
rect 27970 33294 27972 33346
rect 27916 33282 27972 33294
rect 27244 31778 27300 32956
rect 28028 32788 28084 34636
rect 28588 34598 28644 34636
rect 28364 34020 28420 34030
rect 28364 33926 28420 33964
rect 28700 33572 28756 36206
rect 28364 33516 28700 33572
rect 28252 33460 28308 33470
rect 28252 33366 28308 33404
rect 28364 33346 28420 33516
rect 28700 33478 28756 33516
rect 28364 33294 28366 33346
rect 28418 33294 28420 33346
rect 28140 33236 28196 33246
rect 28140 33142 28196 33180
rect 28364 33124 28420 33294
rect 28588 33348 28644 33358
rect 28588 33254 28644 33292
rect 28364 33058 28420 33068
rect 28028 32732 28532 32788
rect 27356 32562 27412 32574
rect 27356 32510 27358 32562
rect 27410 32510 27412 32562
rect 27356 31890 27412 32510
rect 27580 32562 27636 32574
rect 27580 32510 27582 32562
rect 27634 32510 27636 32562
rect 27356 31838 27358 31890
rect 27410 31838 27412 31890
rect 27356 31826 27412 31838
rect 27468 32004 27524 32014
rect 27244 31726 27246 31778
rect 27298 31726 27300 31778
rect 27244 31714 27300 31726
rect 27468 31778 27524 31948
rect 27580 31892 27636 32510
rect 27804 32562 27860 32574
rect 27804 32510 27806 32562
rect 27858 32510 27860 32562
rect 27692 32452 27748 32462
rect 27692 32358 27748 32396
rect 27580 31826 27636 31836
rect 27468 31726 27470 31778
rect 27522 31726 27524 31778
rect 27468 31714 27524 31726
rect 26572 31276 26964 31332
rect 27020 31276 27188 31332
rect 26572 31220 26628 31276
rect 26124 30706 26180 30716
rect 26460 31164 26628 31220
rect 25900 30210 25956 30222
rect 25900 30158 25902 30210
rect 25954 30158 25956 30210
rect 25900 30100 25956 30158
rect 25900 30034 25956 30044
rect 26348 30100 26404 30110
rect 25788 29026 25844 29036
rect 26012 29092 26068 29102
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24780 27010 24836 27022
rect 25452 28588 25620 28644
rect 25228 26964 25284 26974
rect 24780 26516 24836 26526
rect 24668 26514 24836 26516
rect 24668 26462 24782 26514
rect 24834 26462 24836 26514
rect 24668 26460 24836 26462
rect 24780 26450 24836 26460
rect 24668 25618 24724 25630
rect 24668 25566 24670 25618
rect 24722 25566 24724 25618
rect 24668 25508 24724 25566
rect 25116 25508 25172 25518
rect 24668 25506 25172 25508
rect 24668 25454 25118 25506
rect 25170 25454 25172 25506
rect 24668 25452 25172 25454
rect 24556 25330 24612 25340
rect 24556 24610 24612 24622
rect 24556 24558 24558 24610
rect 24610 24558 24612 24610
rect 24444 24500 24500 24510
rect 24444 24406 24500 24444
rect 24556 23380 24612 24558
rect 24332 23324 24500 23380
rect 24220 23268 24276 23278
rect 24220 23174 24276 23212
rect 23884 22530 23940 22540
rect 23996 23154 24052 23166
rect 23996 23102 23998 23154
rect 24050 23102 24052 23154
rect 23996 21588 24052 23102
rect 24332 23154 24388 23166
rect 24332 23102 24334 23154
rect 24386 23102 24388 23154
rect 24332 22148 24388 23102
rect 24332 21812 24388 22092
rect 24332 21718 24388 21756
rect 24108 21700 24164 21710
rect 24108 21606 24164 21644
rect 23996 21494 24052 21532
rect 23772 21410 23828 21420
rect 24220 21474 24276 21486
rect 24220 21422 24222 21474
rect 24274 21422 24276 21474
rect 23100 19294 23102 19346
rect 23154 19294 23156 19346
rect 23100 19282 23156 19294
rect 23212 21084 23492 21140
rect 23660 21362 23716 21374
rect 23660 21310 23662 21362
rect 23714 21310 23716 21362
rect 23100 19012 23156 19022
rect 22764 17614 22766 17666
rect 22818 17614 22820 17666
rect 21756 17444 21812 17454
rect 22092 17444 22148 17454
rect 21532 17442 22148 17444
rect 21532 17390 21758 17442
rect 21810 17390 22094 17442
rect 22146 17390 22148 17442
rect 21532 17388 22148 17390
rect 21756 17378 21812 17388
rect 21420 16322 21476 16334
rect 21420 16270 21422 16322
rect 21474 16270 21476 16322
rect 21420 16212 21476 16270
rect 21420 16210 21588 16212
rect 21420 16158 21422 16210
rect 21474 16158 21588 16210
rect 21420 16156 21588 16158
rect 21420 16146 21476 16156
rect 21532 15538 21588 16156
rect 21868 15876 21924 15886
rect 21868 15782 21924 15820
rect 21532 15486 21534 15538
rect 21586 15486 21588 15538
rect 21532 15474 21588 15486
rect 21980 15148 22036 17388
rect 22092 17378 22148 17388
rect 22764 16772 22820 17614
rect 22876 18340 22932 18350
rect 22876 16994 22932 18284
rect 22988 18338 23044 18350
rect 22988 18286 22990 18338
rect 23042 18286 23044 18338
rect 22988 18116 23044 18286
rect 22988 18050 23044 18060
rect 23100 17666 23156 18956
rect 23100 17614 23102 17666
rect 23154 17614 23156 17666
rect 23100 17602 23156 17614
rect 23212 17556 23268 21084
rect 23660 20804 23716 21310
rect 23996 20804 24052 20814
rect 23660 20802 24052 20804
rect 23660 20750 23998 20802
rect 24050 20750 24052 20802
rect 23660 20748 24052 20750
rect 23660 20242 23716 20748
rect 23996 20738 24052 20748
rect 24220 20692 24276 21422
rect 24220 20626 24276 20636
rect 23660 20190 23662 20242
rect 23714 20190 23716 20242
rect 23660 20178 23716 20190
rect 24332 20244 24388 20254
rect 23436 20132 23492 20142
rect 23324 20020 23380 20030
rect 23324 19906 23380 19964
rect 23324 19854 23326 19906
rect 23378 19854 23380 19906
rect 23324 19842 23380 19854
rect 23324 18452 23380 18462
rect 23436 18452 23492 20076
rect 24332 20130 24388 20188
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 20066 24388 20078
rect 23772 20020 23828 20030
rect 23772 19926 23828 19964
rect 24332 18452 24388 18462
rect 24444 18452 24500 23324
rect 24556 23314 24612 23324
rect 25116 21700 25172 25452
rect 25228 25506 25284 26908
rect 25452 26852 25508 28588
rect 25788 28532 25844 28542
rect 25788 28438 25844 28476
rect 26012 27748 26068 29036
rect 26348 28868 26404 30044
rect 26460 29986 26516 31164
rect 26684 31108 26740 31118
rect 26684 31014 26740 31052
rect 26460 29934 26462 29986
rect 26514 29934 26516 29986
rect 26460 29764 26516 29934
rect 26460 29698 26516 29708
rect 26572 30882 26628 30894
rect 26572 30830 26574 30882
rect 26626 30830 26628 30882
rect 26572 29092 26628 30830
rect 26684 30772 26740 30782
rect 26684 30210 26740 30716
rect 26796 30324 26852 30334
rect 26796 30230 26852 30268
rect 26684 30158 26686 30210
rect 26738 30158 26740 30210
rect 26684 30146 26740 30158
rect 26908 29988 26964 29998
rect 26908 29894 26964 29932
rect 26628 29036 26964 29092
rect 26572 29026 26628 29036
rect 26572 28868 26628 28878
rect 26796 28868 26852 28878
rect 26348 28812 26516 28868
rect 26236 28756 26292 28766
rect 26292 28700 26404 28756
rect 26236 28690 26292 28700
rect 26124 28642 26180 28654
rect 26124 28590 26126 28642
rect 26178 28590 26180 28642
rect 26124 27972 26180 28590
rect 26236 28420 26292 28430
rect 26236 28326 26292 28364
rect 26124 27858 26180 27916
rect 26124 27806 26126 27858
rect 26178 27806 26180 27858
rect 26124 27794 26180 27806
rect 26348 27858 26404 28700
rect 26460 28642 26516 28812
rect 26628 28812 26740 28868
rect 26572 28802 26628 28812
rect 26460 28590 26462 28642
rect 26514 28590 26516 28642
rect 26460 28578 26516 28590
rect 26684 28642 26740 28812
rect 26684 28590 26686 28642
rect 26738 28590 26740 28642
rect 26684 28578 26740 28590
rect 26572 28420 26628 28430
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26348 27794 26404 27806
rect 26460 28364 26572 28420
rect 25676 27746 26068 27748
rect 25676 27694 26014 27746
rect 26066 27694 26068 27746
rect 25676 27692 26068 27694
rect 25676 26962 25732 27692
rect 26012 27682 26068 27692
rect 26460 27636 26516 28364
rect 26572 28354 26628 28364
rect 26796 28084 26852 28812
rect 26908 28866 26964 29036
rect 26908 28814 26910 28866
rect 26962 28814 26964 28866
rect 26908 28802 26964 28814
rect 25676 26910 25678 26962
rect 25730 26910 25732 26962
rect 25676 26898 25732 26910
rect 26348 27580 26516 27636
rect 26572 28082 26852 28084
rect 26572 28030 26798 28082
rect 26850 28030 26852 28082
rect 26572 28028 26852 28030
rect 26124 26852 26180 26862
rect 25452 26290 25508 26796
rect 26012 26796 26124 26852
rect 26012 26404 26068 26796
rect 26124 26758 26180 26796
rect 26012 26338 26068 26348
rect 26236 26404 26292 26414
rect 26236 26310 26292 26348
rect 25452 26238 25454 26290
rect 25506 26238 25508 26290
rect 25452 26226 25508 26238
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 25228 24946 25284 25454
rect 25564 25732 25620 25742
rect 25452 25396 25508 25434
rect 25452 25330 25508 25340
rect 25564 25396 25620 25676
rect 26236 25508 26292 25518
rect 26124 25506 26292 25508
rect 26124 25454 26238 25506
rect 26290 25454 26292 25506
rect 26124 25452 26292 25454
rect 26012 25396 26068 25406
rect 25564 25394 26068 25396
rect 25564 25342 25566 25394
rect 25618 25342 26014 25394
rect 26066 25342 26068 25394
rect 25564 25340 26068 25342
rect 25564 25330 25620 25340
rect 26012 25330 26068 25340
rect 25340 25284 25396 25294
rect 25340 25190 25396 25228
rect 26124 25284 26180 25452
rect 26236 25442 26292 25452
rect 25228 24894 25230 24946
rect 25282 24894 25284 24946
rect 25228 24882 25284 24894
rect 25564 24724 25620 24734
rect 25564 24722 25844 24724
rect 25564 24670 25566 24722
rect 25618 24670 25844 24722
rect 25564 24668 25844 24670
rect 25564 24658 25620 24668
rect 25676 24164 25732 24174
rect 25340 23828 25396 23838
rect 25340 23734 25396 23772
rect 25228 23156 25284 23166
rect 25228 22482 25284 23100
rect 25564 23156 25620 23166
rect 25564 23062 25620 23100
rect 25228 22430 25230 22482
rect 25282 22430 25284 22482
rect 25228 22418 25284 22430
rect 25676 22258 25732 24108
rect 25788 23378 25844 24668
rect 25788 23326 25790 23378
rect 25842 23326 25844 23378
rect 25788 23156 25844 23326
rect 25900 23380 25956 23390
rect 25900 23286 25956 23324
rect 26124 23380 26180 25228
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 23492 26292 24558
rect 26236 23426 26292 23436
rect 26124 23286 26180 23324
rect 26012 23268 26068 23278
rect 26012 23174 26068 23212
rect 25788 23090 25844 23100
rect 26348 22932 26404 27580
rect 26460 27076 26516 27086
rect 26460 26982 26516 27020
rect 25788 22876 26404 22932
rect 26460 26740 26516 26750
rect 25788 22708 25844 22876
rect 25788 22370 25844 22652
rect 25788 22318 25790 22370
rect 25842 22318 25844 22370
rect 25788 22306 25844 22318
rect 25676 22206 25678 22258
rect 25730 22206 25732 22258
rect 25676 22194 25732 22206
rect 25452 22148 25508 22158
rect 26348 22148 26404 22158
rect 25452 22054 25508 22092
rect 26124 22146 26404 22148
rect 26124 22094 26350 22146
rect 26402 22094 26404 22146
rect 26124 22092 26404 22094
rect 26124 21810 26180 22092
rect 26348 22082 26404 22092
rect 26124 21758 26126 21810
rect 26178 21758 26180 21810
rect 25228 21700 25284 21710
rect 25116 21698 25284 21700
rect 25116 21646 25230 21698
rect 25282 21646 25284 21698
rect 25116 21644 25284 21646
rect 25228 21634 25284 21644
rect 26124 21700 26180 21758
rect 26460 21812 26516 26684
rect 26572 24164 26628 28028
rect 26796 28018 26852 28028
rect 26796 25396 26852 25406
rect 26796 25302 26852 25340
rect 26572 24098 26628 24108
rect 26796 24836 26852 24846
rect 26796 23716 26852 24780
rect 26684 23492 26740 23502
rect 26684 23266 26740 23436
rect 26684 23214 26686 23266
rect 26738 23214 26740 23266
rect 26684 23202 26740 23214
rect 26572 23044 26628 23054
rect 26572 22950 26628 22988
rect 26796 22482 26852 23660
rect 27020 23548 27076 31276
rect 27244 30324 27300 30334
rect 27244 30210 27300 30268
rect 27244 30158 27246 30210
rect 27298 30158 27300 30210
rect 27244 30146 27300 30158
rect 27580 30210 27636 30222
rect 27580 30158 27582 30210
rect 27634 30158 27636 30210
rect 27580 29876 27636 30158
rect 27804 30210 27860 32510
rect 28140 32564 28196 32574
rect 28028 32004 28084 32014
rect 28028 31910 28084 31948
rect 28140 31666 28196 32508
rect 28140 31614 28142 31666
rect 28194 31614 28196 31666
rect 28140 31602 28196 31614
rect 28252 32450 28308 32462
rect 28252 32398 28254 32450
rect 28306 32398 28308 32450
rect 27916 31108 27972 31118
rect 28252 31108 28308 32398
rect 27972 31052 28308 31108
rect 28364 32228 28420 32238
rect 28364 31554 28420 32172
rect 28364 31502 28366 31554
rect 28418 31502 28420 31554
rect 28364 31444 28420 31502
rect 27916 31014 27972 31052
rect 28364 30994 28420 31388
rect 28476 31332 28532 32732
rect 29036 32676 29092 41132
rect 29372 40964 29428 40974
rect 29260 40962 29428 40964
rect 29260 40910 29374 40962
rect 29426 40910 29428 40962
rect 29260 40908 29428 40910
rect 29148 39396 29204 39406
rect 29260 39396 29316 40908
rect 29372 40898 29428 40908
rect 29484 40962 29540 40974
rect 29484 40910 29486 40962
rect 29538 40910 29540 40962
rect 29484 40628 29540 40910
rect 29484 40562 29540 40572
rect 29596 40962 29652 40974
rect 29596 40910 29598 40962
rect 29650 40910 29652 40962
rect 29372 40516 29428 40526
rect 29372 40422 29428 40460
rect 29484 40178 29540 40190
rect 29484 40126 29486 40178
rect 29538 40126 29540 40178
rect 29484 40068 29540 40126
rect 29484 40002 29540 40012
rect 29596 39732 29652 40910
rect 29708 40964 29764 40974
rect 29708 40290 29764 40908
rect 29708 40238 29710 40290
rect 29762 40238 29764 40290
rect 29708 40226 29764 40238
rect 29820 40290 29876 42700
rect 29932 41972 29988 43708
rect 30044 42756 30100 43820
rect 30156 43650 30212 43662
rect 30156 43598 30158 43650
rect 30210 43598 30212 43650
rect 30156 43316 30212 43598
rect 30268 43652 30324 43662
rect 30324 43596 30436 43652
rect 30268 43586 30324 43596
rect 30156 43250 30212 43260
rect 30044 42662 30100 42700
rect 30380 42868 30436 43596
rect 30716 43538 30772 44156
rect 30716 43486 30718 43538
rect 30770 43486 30772 43538
rect 30716 43474 30772 43486
rect 30492 43426 30548 43438
rect 30492 43374 30494 43426
rect 30546 43374 30548 43426
rect 30492 43316 30548 43374
rect 30492 43250 30548 43260
rect 30940 42980 30996 44156
rect 31164 44098 31220 44110
rect 31164 44046 31166 44098
rect 31218 44046 31220 44098
rect 31052 43764 31108 43774
rect 31052 43650 31108 43708
rect 31052 43598 31054 43650
rect 31106 43598 31108 43650
rect 31052 43586 31108 43598
rect 31164 43316 31220 44046
rect 31724 43538 31780 44492
rect 32508 44434 32564 44446
rect 32508 44382 32510 44434
rect 32562 44382 32564 44434
rect 32172 44212 32228 44222
rect 31724 43486 31726 43538
rect 31778 43486 31780 43538
rect 31724 43474 31780 43486
rect 31836 44210 32228 44212
rect 31836 44158 32174 44210
rect 32226 44158 32228 44210
rect 31836 44156 32228 44158
rect 31836 43764 31892 44156
rect 32172 44146 32228 44156
rect 32396 44100 32452 44110
rect 31836 43538 31892 43708
rect 31836 43486 31838 43538
rect 31890 43486 31892 43538
rect 31836 43474 31892 43486
rect 32284 44098 32452 44100
rect 32284 44046 32398 44098
rect 32450 44046 32452 44098
rect 32284 44044 32452 44046
rect 31388 43428 31444 43438
rect 31388 43334 31444 43372
rect 31276 43316 31332 43326
rect 31164 43260 31276 43316
rect 31276 43250 31332 43260
rect 31500 43314 31556 43326
rect 31500 43262 31502 43314
rect 31554 43262 31556 43314
rect 31052 43204 31108 43214
rect 31108 43148 31220 43204
rect 31052 43138 31108 43148
rect 31052 42980 31108 42990
rect 30940 42978 31108 42980
rect 30940 42926 31054 42978
rect 31106 42926 31108 42978
rect 30940 42924 31108 42926
rect 30492 42868 30548 42878
rect 30380 42866 30548 42868
rect 30380 42814 30494 42866
rect 30546 42814 30548 42866
rect 30380 42812 30548 42814
rect 29932 41906 29988 41916
rect 30156 42532 30212 42542
rect 30156 41970 30212 42476
rect 30268 42530 30324 42542
rect 30268 42478 30270 42530
rect 30322 42478 30324 42530
rect 30268 42308 30324 42478
rect 30268 42242 30324 42252
rect 30156 41918 30158 41970
rect 30210 41918 30212 41970
rect 30156 41906 30212 41918
rect 30044 41412 30100 41422
rect 30044 41186 30100 41356
rect 30268 41300 30324 41310
rect 30268 41206 30324 41244
rect 30044 41134 30046 41186
rect 30098 41134 30100 41186
rect 30044 41122 30100 41134
rect 29820 40238 29822 40290
rect 29874 40238 29876 40290
rect 29820 40226 29876 40238
rect 30380 40402 30436 42812
rect 30492 42802 30548 42812
rect 30716 42756 30772 42766
rect 30772 42700 30884 42756
rect 30716 42662 30772 42700
rect 30716 41412 30772 41422
rect 30492 41186 30548 41198
rect 30492 41134 30494 41186
rect 30546 41134 30548 41186
rect 30492 40740 30548 41134
rect 30716 40740 30772 41356
rect 30828 41410 30884 42700
rect 30940 41970 30996 42924
rect 31052 42914 31108 42924
rect 31052 42196 31108 42206
rect 31164 42196 31220 43148
rect 31500 42756 31556 43262
rect 31052 42194 31220 42196
rect 31052 42142 31054 42194
rect 31106 42142 31220 42194
rect 31052 42140 31220 42142
rect 31388 42700 31556 42756
rect 32284 42868 32340 44044
rect 32396 44034 32452 44044
rect 32508 42978 32564 44382
rect 39228 44436 39284 44446
rect 39228 44342 39284 44380
rect 34524 44324 34580 44334
rect 33852 44322 34580 44324
rect 33852 44270 34526 44322
rect 34578 44270 34580 44322
rect 33852 44268 34580 44270
rect 33404 44210 33460 44222
rect 33404 44158 33406 44210
rect 33458 44158 33460 44210
rect 33180 44098 33236 44110
rect 33180 44046 33182 44098
rect 33234 44046 33236 44098
rect 32620 43652 32676 43662
rect 32620 43558 32676 43596
rect 32508 42926 32510 42978
rect 32562 42926 32564 42978
rect 32508 42914 32564 42926
rect 32844 43428 32900 43438
rect 33068 43428 33124 43438
rect 32844 42978 32900 43372
rect 32844 42926 32846 42978
rect 32898 42926 32900 42978
rect 32844 42914 32900 42926
rect 32956 43426 33124 43428
rect 32956 43374 33070 43426
rect 33122 43374 33124 43426
rect 32956 43372 33124 43374
rect 31052 42130 31108 42140
rect 30940 41918 30942 41970
rect 30994 41918 30996 41970
rect 30940 41906 30996 41918
rect 31164 41972 31220 41982
rect 31164 41878 31220 41916
rect 30828 41358 30830 41410
rect 30882 41358 30884 41410
rect 30828 41346 30884 41358
rect 31388 41746 31444 42700
rect 31500 42532 31556 42542
rect 31500 42438 31556 42476
rect 31948 42532 32004 42542
rect 31948 42438 32004 42476
rect 32172 42082 32228 42094
rect 32172 42030 32174 42082
rect 32226 42030 32228 42082
rect 31836 41972 31892 41982
rect 31388 41694 31390 41746
rect 31442 41694 31444 41746
rect 31388 41412 31444 41694
rect 31388 41346 31444 41356
rect 31724 41970 31892 41972
rect 31724 41918 31838 41970
rect 31890 41918 31892 41970
rect 31724 41916 31892 41918
rect 31164 41074 31220 41086
rect 31164 41022 31166 41074
rect 31218 41022 31220 41074
rect 31164 40852 31220 41022
rect 31276 40964 31332 40974
rect 31276 40870 31332 40908
rect 31388 40962 31444 40974
rect 31388 40910 31390 40962
rect 31442 40910 31444 40962
rect 31164 40786 31220 40796
rect 30492 40674 30548 40684
rect 30604 40684 30716 40740
rect 30604 40626 30660 40684
rect 30716 40674 30772 40684
rect 31388 40628 31444 40910
rect 30604 40574 30606 40626
rect 30658 40574 30660 40626
rect 30604 40562 30660 40574
rect 30828 40572 31444 40628
rect 30492 40516 30548 40526
rect 30492 40422 30548 40460
rect 30716 40516 30772 40554
rect 30716 40450 30772 40460
rect 30380 40350 30382 40402
rect 30434 40350 30436 40402
rect 30268 39956 30324 39966
rect 30268 39842 30324 39900
rect 30268 39790 30270 39842
rect 30322 39790 30324 39842
rect 29708 39732 29764 39742
rect 29596 39676 29708 39732
rect 29708 39638 29764 39676
rect 29820 39620 29876 39630
rect 29820 39526 29876 39564
rect 29932 39618 29988 39630
rect 29932 39566 29934 39618
rect 29986 39566 29988 39618
rect 29596 39396 29652 39406
rect 29708 39396 29764 39406
rect 29260 39340 29540 39396
rect 29148 39172 29204 39340
rect 29148 39106 29204 39116
rect 29372 38948 29428 38958
rect 29372 38854 29428 38892
rect 29260 38836 29316 38846
rect 29260 38742 29316 38780
rect 29148 38722 29204 38734
rect 29148 38670 29150 38722
rect 29202 38670 29204 38722
rect 29148 38612 29204 38670
rect 29148 38546 29204 38556
rect 29484 38162 29540 39340
rect 29596 39394 29708 39396
rect 29596 39342 29598 39394
rect 29650 39342 29708 39394
rect 29596 39340 29708 39342
rect 29596 39330 29652 39340
rect 29484 38110 29486 38162
rect 29538 38110 29540 38162
rect 29484 38098 29540 38110
rect 29596 38948 29652 38958
rect 29372 38052 29428 38062
rect 29372 37958 29428 37996
rect 29596 38050 29652 38892
rect 29596 37998 29598 38050
rect 29650 37998 29652 38050
rect 29596 37986 29652 37998
rect 29148 37940 29204 37950
rect 29148 37846 29204 37884
rect 29260 36596 29316 36606
rect 29148 36594 29316 36596
rect 29148 36542 29262 36594
rect 29314 36542 29316 36594
rect 29148 36540 29316 36542
rect 29148 35476 29204 36540
rect 29260 36530 29316 36540
rect 29372 36484 29428 36494
rect 29260 36258 29316 36270
rect 29260 36206 29262 36258
rect 29314 36206 29316 36258
rect 29260 35924 29316 36206
rect 29260 35858 29316 35868
rect 29372 36258 29428 36428
rect 29596 36372 29652 36382
rect 29596 36278 29652 36316
rect 29372 36206 29374 36258
rect 29426 36206 29428 36258
rect 29148 35410 29204 35420
rect 29372 35364 29428 36206
rect 29260 35308 29428 35364
rect 29708 35308 29764 39340
rect 29820 39172 29876 39182
rect 29820 39058 29876 39116
rect 29820 39006 29822 39058
rect 29874 39006 29876 39058
rect 29820 38994 29876 39006
rect 29932 38612 29988 39566
rect 30268 38948 30324 39790
rect 30380 39620 30436 40350
rect 30828 39956 30884 40572
rect 31724 40516 31780 41916
rect 31836 41906 31892 41916
rect 32172 41412 32228 42030
rect 32172 41346 32228 41356
rect 32284 41300 32340 42812
rect 32956 42868 33012 43372
rect 33068 43362 33124 43372
rect 33180 42868 33236 44046
rect 33404 43988 33460 44158
rect 33516 44212 33572 44222
rect 33516 44118 33572 44156
rect 33852 44210 33908 44268
rect 34524 44258 34580 44268
rect 34860 44322 34916 44334
rect 34860 44270 34862 44322
rect 34914 44270 34916 44322
rect 33852 44158 33854 44210
rect 33906 44158 33908 44210
rect 33404 43922 33460 43932
rect 32956 42802 33012 42812
rect 33068 42812 33236 42868
rect 33516 42866 33572 42878
rect 33516 42814 33518 42866
rect 33570 42814 33572 42866
rect 32396 42754 32452 42766
rect 32396 42702 32398 42754
rect 32450 42702 32452 42754
rect 32396 42308 32452 42702
rect 32732 42754 32788 42766
rect 32732 42702 32734 42754
rect 32786 42702 32788 42754
rect 32396 42242 32452 42252
rect 32508 42644 32564 42654
rect 32396 41300 32452 41310
rect 32284 41298 32452 41300
rect 32284 41246 32398 41298
rect 32450 41246 32452 41298
rect 32284 41244 32452 41246
rect 32396 41234 32452 41244
rect 31948 41076 32004 41086
rect 31948 40982 32004 41020
rect 30940 40404 30996 40414
rect 31276 40404 31332 40414
rect 30940 40402 31332 40404
rect 30940 40350 30942 40402
rect 30994 40350 31278 40402
rect 31330 40350 31332 40402
rect 30940 40348 31332 40350
rect 30940 40338 30996 40348
rect 31276 40338 31332 40348
rect 31388 40292 31444 40302
rect 30828 39890 30884 39900
rect 31276 40068 31332 40078
rect 31164 39844 31220 39854
rect 30940 39842 31220 39844
rect 30940 39790 31166 39842
rect 31218 39790 31220 39842
rect 30940 39788 31220 39790
rect 30380 39554 30436 39564
rect 30492 39732 30548 39742
rect 30268 38882 30324 38892
rect 30492 38834 30548 39676
rect 30492 38782 30494 38834
rect 30546 38782 30548 38834
rect 30492 38770 30548 38782
rect 30604 39506 30660 39518
rect 30604 39454 30606 39506
rect 30658 39454 30660 39506
rect 30604 38668 30660 39454
rect 30716 39396 30772 39406
rect 30716 38834 30772 39340
rect 30828 39394 30884 39406
rect 30828 39342 30830 39394
rect 30882 39342 30884 39394
rect 30828 39284 30884 39342
rect 30828 39218 30884 39228
rect 30716 38782 30718 38834
rect 30770 38782 30772 38834
rect 30716 38770 30772 38782
rect 30940 38834 30996 39788
rect 31164 39778 31220 39788
rect 31164 39618 31220 39630
rect 31164 39566 31166 39618
rect 31218 39566 31220 39618
rect 30940 38782 30942 38834
rect 30994 38782 30996 38834
rect 30940 38770 30996 38782
rect 31052 39394 31108 39406
rect 31052 39342 31054 39394
rect 31106 39342 31108 39394
rect 29820 38052 29876 38062
rect 29932 38052 29988 38556
rect 30492 38612 30660 38668
rect 29820 38050 29988 38052
rect 29820 37998 29822 38050
rect 29874 37998 29988 38050
rect 29820 37996 29988 37998
rect 29820 37986 29876 37996
rect 29932 37716 29988 37996
rect 30156 38164 30212 38174
rect 30156 38050 30212 38108
rect 30156 37998 30158 38050
rect 30210 37998 30212 38050
rect 30156 37986 30212 37998
rect 30492 38052 30548 38612
rect 30492 37958 30548 37996
rect 30604 38500 30660 38510
rect 29820 37660 29988 37716
rect 30268 37828 30324 37838
rect 29820 37156 29876 37660
rect 29932 37380 29988 37390
rect 30268 37380 30324 37772
rect 30604 37604 30660 38444
rect 31052 38388 31108 39342
rect 31164 39060 31220 39566
rect 31164 38994 31220 39004
rect 31276 38836 31332 40012
rect 31388 39172 31444 40236
rect 31724 40068 31780 40460
rect 31836 40962 31892 40974
rect 31836 40910 31838 40962
rect 31890 40910 31892 40962
rect 31836 40402 31892 40910
rect 32284 40962 32340 40974
rect 32284 40910 32286 40962
rect 32338 40910 32340 40962
rect 31948 40628 32004 40638
rect 32172 40628 32228 40638
rect 32284 40628 32340 40910
rect 32004 40572 32116 40628
rect 31948 40562 32004 40572
rect 31836 40350 31838 40402
rect 31890 40350 31892 40402
rect 31836 40338 31892 40350
rect 31948 40402 32004 40414
rect 31948 40350 31950 40402
rect 32002 40350 32004 40402
rect 31948 40292 32004 40350
rect 31948 40226 32004 40236
rect 31724 40002 31780 40012
rect 31724 39732 31780 39742
rect 31612 39620 31668 39630
rect 31612 39526 31668 39564
rect 31724 39506 31780 39676
rect 32060 39620 32116 40572
rect 32172 40626 32284 40628
rect 32172 40574 32174 40626
rect 32226 40574 32284 40626
rect 32172 40572 32284 40574
rect 32172 40562 32228 40572
rect 32284 40562 32340 40572
rect 32396 40404 32452 40414
rect 32396 40310 32452 40348
rect 32284 40290 32340 40302
rect 32284 40238 32286 40290
rect 32338 40238 32340 40290
rect 32284 39844 32340 40238
rect 32508 40180 32564 42588
rect 32732 41412 32788 42702
rect 33068 42532 33124 42812
rect 33404 42756 33460 42766
rect 33068 42466 33124 42476
rect 33180 42642 33236 42654
rect 33180 42590 33182 42642
rect 33234 42590 33236 42642
rect 33180 42308 33236 42590
rect 33404 42642 33460 42700
rect 33404 42590 33406 42642
rect 33458 42590 33460 42642
rect 33404 42578 33460 42590
rect 33180 42242 33236 42252
rect 33404 42420 33460 42430
rect 33068 41858 33124 41870
rect 33068 41806 33070 41858
rect 33122 41806 33124 41858
rect 33068 41748 33124 41806
rect 33068 41682 33124 41692
rect 33180 41860 33236 41870
rect 32732 41346 32788 41356
rect 33180 41410 33236 41804
rect 33180 41358 33182 41410
rect 33234 41358 33236 41410
rect 33180 41346 33236 41358
rect 33292 41412 33348 41422
rect 33292 41318 33348 41356
rect 33404 41188 33460 42364
rect 33516 41412 33572 42814
rect 33852 42420 33908 44158
rect 34860 44212 34916 44270
rect 36428 44322 36484 44334
rect 36428 44270 36430 44322
rect 36482 44270 36484 44322
rect 33964 44098 34020 44110
rect 33964 44046 33966 44098
rect 34018 44046 34020 44098
rect 33964 43988 34020 44046
rect 34188 44100 34244 44110
rect 34188 44006 34244 44044
rect 33964 43922 34020 43932
rect 34860 42980 34916 44156
rect 35420 44212 35476 44222
rect 35420 44210 35588 44212
rect 35420 44158 35422 44210
rect 35474 44158 35588 44210
rect 35420 44156 35588 44158
rect 35420 44146 35476 44156
rect 35196 43428 35252 43438
rect 35196 43334 35252 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34188 42756 34244 42766
rect 34636 42756 34692 42766
rect 34244 42700 34356 42756
rect 34188 42690 34244 42700
rect 33852 42354 33908 42364
rect 33628 41412 33684 41422
rect 33516 41410 33684 41412
rect 33516 41358 33630 41410
rect 33682 41358 33684 41410
rect 33516 41356 33684 41358
rect 33628 41346 33684 41356
rect 33516 41188 33572 41198
rect 33404 41186 33572 41188
rect 33404 41134 33518 41186
rect 33570 41134 33572 41186
rect 33404 41132 33572 41134
rect 33516 41122 33572 41132
rect 33852 41188 33908 41198
rect 32844 40964 32900 40974
rect 32284 39778 32340 39788
rect 32396 40124 32564 40180
rect 32620 40962 32900 40964
rect 32620 40910 32846 40962
rect 32898 40910 32900 40962
rect 32620 40908 32900 40910
rect 32060 39564 32340 39620
rect 31724 39454 31726 39506
rect 31778 39454 31780 39506
rect 31724 39442 31780 39454
rect 32284 39506 32340 39564
rect 32284 39454 32286 39506
rect 32338 39454 32340 39506
rect 32284 39442 32340 39454
rect 31948 39396 32004 39406
rect 31948 39302 32004 39340
rect 32172 39172 32228 39182
rect 31388 39116 31668 39172
rect 31052 38322 31108 38332
rect 31164 38780 31332 38836
rect 30716 38276 30772 38286
rect 30716 38050 30772 38220
rect 30716 37998 30718 38050
rect 30770 37998 30772 38050
rect 30716 37986 30772 37998
rect 31052 38052 31108 38062
rect 31164 38052 31220 38780
rect 31388 38612 31444 38622
rect 31388 38610 31556 38612
rect 31388 38558 31390 38610
rect 31442 38558 31556 38610
rect 31388 38556 31556 38558
rect 31388 38546 31444 38556
rect 31052 38050 31220 38052
rect 31052 37998 31054 38050
rect 31106 37998 31220 38050
rect 31052 37996 31220 37998
rect 31388 38050 31444 38062
rect 31388 37998 31390 38050
rect 31442 37998 31444 38050
rect 31052 37986 31108 37996
rect 30828 37828 30884 37838
rect 30828 37826 30996 37828
rect 30828 37774 30830 37826
rect 30882 37774 30996 37826
rect 30828 37772 30996 37774
rect 30828 37762 30884 37772
rect 30604 37548 30884 37604
rect 30828 37490 30884 37548
rect 30828 37438 30830 37490
rect 30882 37438 30884 37490
rect 30828 37426 30884 37438
rect 30940 37492 30996 37772
rect 30940 37426 30996 37436
rect 31388 37490 31444 37998
rect 31388 37438 31390 37490
rect 31442 37438 31444 37490
rect 31388 37426 31444 37438
rect 29932 37378 30324 37380
rect 29932 37326 29934 37378
rect 29986 37326 30324 37378
rect 29932 37324 30324 37326
rect 29932 37314 29988 37324
rect 31276 37268 31332 37278
rect 31500 37268 31556 38556
rect 31276 37266 31556 37268
rect 31276 37214 31278 37266
rect 31330 37214 31556 37266
rect 31276 37212 31556 37214
rect 31276 37202 31332 37212
rect 30268 37156 30324 37166
rect 29820 37154 30324 37156
rect 29820 37102 30270 37154
rect 30322 37102 30324 37154
rect 29820 37100 30324 37102
rect 30268 37090 30324 37100
rect 30380 37154 30436 37166
rect 30380 37102 30382 37154
rect 30434 37102 30436 37154
rect 29820 36370 29876 36382
rect 29820 36318 29822 36370
rect 29874 36318 29876 36370
rect 29820 36148 29876 36318
rect 29820 36082 29876 36092
rect 29932 36372 29988 36382
rect 29932 35700 29988 36316
rect 30268 36372 30324 36382
rect 30268 36278 30324 36316
rect 30156 36260 30212 36270
rect 30156 36166 30212 36204
rect 30044 35924 30100 35934
rect 30100 35868 30212 35924
rect 30044 35858 30100 35868
rect 29932 35634 29988 35644
rect 29260 35252 29316 35308
rect 29148 35196 29316 35252
rect 29484 35252 29764 35308
rect 29148 34468 29204 35196
rect 29372 35140 29428 35150
rect 29484 35140 29540 35252
rect 29372 35138 29540 35140
rect 29372 35086 29374 35138
rect 29426 35086 29540 35138
rect 29372 35084 29540 35086
rect 29372 35074 29428 35084
rect 29148 34402 29204 34412
rect 29260 34802 29316 34814
rect 29260 34750 29262 34802
rect 29314 34750 29316 34802
rect 29260 34020 29316 34750
rect 30156 34804 30212 35868
rect 30380 35812 30436 37102
rect 31612 37044 31668 39116
rect 32172 39058 32228 39116
rect 32172 39006 32174 39058
rect 32226 39006 32228 39058
rect 32172 38994 32228 39006
rect 31724 38948 31780 38958
rect 31724 38724 31780 38892
rect 31724 38658 31780 38668
rect 31948 38164 32004 38174
rect 31836 38052 31892 38062
rect 31836 37958 31892 37996
rect 31948 37268 32004 38108
rect 32396 37828 32452 40124
rect 32508 39732 32564 39742
rect 32508 39618 32564 39676
rect 32508 39566 32510 39618
rect 32562 39566 32564 39618
rect 32508 39554 32564 39566
rect 32508 38276 32564 38286
rect 32508 38182 32564 38220
rect 32396 37716 32452 37772
rect 31836 37154 31892 37166
rect 31836 37102 31838 37154
rect 31890 37102 31892 37154
rect 31388 36988 31668 37044
rect 31724 37042 31780 37054
rect 31724 36990 31726 37042
rect 31778 36990 31780 37042
rect 30828 36482 30884 36494
rect 30828 36430 30830 36482
rect 30882 36430 30884 36482
rect 30716 35812 30772 35822
rect 30380 35810 30772 35812
rect 30380 35758 30718 35810
rect 30770 35758 30772 35810
rect 30380 35756 30772 35758
rect 30380 35586 30436 35756
rect 30716 35746 30772 35756
rect 30380 35534 30382 35586
rect 30434 35534 30436 35586
rect 30380 35522 30436 35534
rect 30268 35364 30324 35374
rect 30268 35026 30324 35308
rect 30716 35364 30772 35374
rect 30828 35364 30884 36430
rect 30940 36372 30996 36382
rect 31388 36372 31444 36988
rect 31724 36932 31780 36990
rect 31500 36876 31780 36932
rect 31836 36932 31892 37102
rect 31500 36594 31556 36876
rect 31836 36866 31892 36876
rect 31948 36708 32004 37212
rect 32284 37660 32452 37716
rect 31500 36542 31502 36594
rect 31554 36542 31556 36594
rect 31500 36530 31556 36542
rect 31724 36652 32004 36708
rect 32172 36932 32228 36942
rect 30996 36316 31108 36372
rect 31388 36316 31556 36372
rect 30940 36306 30996 36316
rect 31052 35922 31108 36316
rect 31388 36036 31444 36046
rect 31052 35870 31054 35922
rect 31106 35870 31108 35922
rect 31052 35858 31108 35870
rect 31276 35924 31332 35934
rect 31276 35830 31332 35868
rect 31164 35812 31220 35822
rect 31164 35718 31220 35756
rect 30940 35700 30996 35710
rect 30940 35476 30996 35644
rect 30940 35420 31332 35476
rect 30772 35308 31220 35364
rect 30716 35298 30772 35308
rect 30268 34974 30270 35026
rect 30322 34974 30324 35026
rect 30268 34962 30324 34974
rect 30156 34748 30324 34804
rect 29148 33572 29204 33582
rect 29148 32786 29204 33516
rect 29260 33348 29316 33964
rect 30044 33460 30100 33470
rect 30044 33366 30100 33404
rect 29484 33348 29540 33358
rect 29260 33346 29540 33348
rect 29260 33294 29486 33346
rect 29538 33294 29540 33346
rect 29260 33292 29540 33294
rect 29484 33282 29540 33292
rect 30156 33348 30212 33358
rect 30268 33348 30324 34748
rect 31164 34130 31220 35308
rect 31164 34078 31166 34130
rect 31218 34078 31220 34130
rect 30492 34018 30548 34030
rect 30492 33966 30494 34018
rect 30546 33966 30548 34018
rect 30492 33796 30548 33966
rect 30492 33730 30548 33740
rect 30604 33684 30660 33694
rect 30212 33292 30548 33348
rect 30156 33254 30212 33292
rect 29708 33236 29764 33246
rect 29708 33142 29764 33180
rect 30492 33234 30548 33292
rect 30492 33182 30494 33234
rect 30546 33182 30548 33234
rect 30492 33170 30548 33182
rect 29932 33124 29988 33134
rect 29932 33030 29988 33068
rect 30492 32900 30548 32910
rect 29148 32734 29150 32786
rect 29202 32734 29204 32786
rect 29148 32722 29204 32734
rect 30380 32844 30492 32900
rect 30380 32786 30436 32844
rect 30492 32834 30548 32844
rect 30380 32734 30382 32786
rect 30434 32734 30436 32786
rect 30380 32722 30436 32734
rect 28700 32620 29092 32676
rect 29596 32676 29652 32686
rect 29652 32620 29764 32676
rect 28700 32228 28756 32620
rect 29596 32582 29652 32620
rect 28812 32452 28868 32462
rect 29484 32452 29540 32462
rect 28812 32450 29092 32452
rect 28812 32398 28814 32450
rect 28866 32398 29092 32450
rect 28812 32396 29092 32398
rect 28812 32386 28868 32396
rect 28700 32172 28868 32228
rect 28588 31668 28644 31678
rect 28588 31574 28644 31612
rect 28476 31266 28532 31276
rect 28364 30942 28366 30994
rect 28418 30942 28420 30994
rect 28364 30930 28420 30942
rect 28812 31108 28868 32172
rect 29036 32004 29092 32396
rect 29036 31948 29316 32004
rect 29036 31780 29092 31948
rect 29260 31890 29316 31948
rect 29260 31838 29262 31890
rect 29314 31838 29316 31890
rect 29260 31826 29316 31838
rect 29036 31714 29092 31724
rect 29484 31108 29540 32396
rect 29708 31890 29764 32620
rect 30492 32452 30548 32462
rect 30604 32452 30660 33628
rect 31164 33572 31220 34078
rect 31164 33506 31220 33516
rect 31052 33348 31108 33358
rect 30828 33122 30884 33134
rect 30828 33070 30830 33122
rect 30882 33070 30884 33122
rect 30828 32564 30884 33070
rect 30940 32564 30996 32574
rect 30828 32562 30996 32564
rect 30828 32510 30942 32562
rect 30994 32510 30996 32562
rect 30828 32508 30996 32510
rect 30492 32450 30660 32452
rect 30492 32398 30494 32450
rect 30546 32398 30660 32450
rect 30492 32396 30660 32398
rect 30492 32386 30548 32396
rect 30156 32340 30212 32350
rect 29708 31838 29710 31890
rect 29762 31838 29764 31890
rect 29708 31444 29764 31838
rect 29708 31378 29764 31388
rect 30044 32284 30156 32340
rect 29596 31108 29652 31118
rect 29484 31106 29652 31108
rect 29484 31054 29598 31106
rect 29650 31054 29652 31106
rect 29484 31052 29652 31054
rect 27804 30158 27806 30210
rect 27858 30158 27860 30210
rect 27804 30100 27860 30158
rect 28476 30210 28532 30222
rect 28476 30158 28478 30210
rect 28530 30158 28532 30210
rect 27804 30034 27860 30044
rect 28140 30098 28196 30110
rect 28140 30046 28142 30098
rect 28194 30046 28196 30098
rect 27692 29988 27748 29998
rect 27692 29894 27748 29932
rect 27580 29810 27636 29820
rect 27132 29428 27188 29438
rect 27132 27860 27188 29372
rect 28140 28980 28196 30046
rect 28252 29986 28308 29998
rect 28252 29934 28254 29986
rect 28306 29934 28308 29986
rect 28252 29092 28308 29934
rect 28252 29036 28420 29092
rect 28140 28924 28308 28980
rect 28140 28756 28196 28766
rect 27804 28644 27860 28654
rect 27804 28550 27860 28588
rect 28140 28642 28196 28700
rect 28140 28590 28142 28642
rect 28194 28590 28196 28642
rect 28140 28578 28196 28590
rect 27244 28420 27300 28430
rect 28252 28420 28308 28924
rect 27244 28418 28308 28420
rect 27244 28366 27246 28418
rect 27298 28366 28308 28418
rect 27244 28364 28308 28366
rect 27244 28354 27300 28364
rect 27244 28084 27300 28094
rect 27244 27990 27300 28028
rect 27132 27804 27860 27860
rect 27580 27300 27636 27310
rect 27580 27206 27636 27244
rect 27692 27076 27748 27086
rect 27692 26962 27748 27020
rect 27692 26910 27694 26962
rect 27746 26910 27748 26962
rect 27692 26898 27748 26910
rect 27132 25394 27188 25406
rect 27132 25342 27134 25394
rect 27186 25342 27188 25394
rect 27132 24052 27188 25342
rect 27244 25282 27300 25294
rect 27244 25230 27246 25282
rect 27298 25230 27300 25282
rect 27244 24948 27300 25230
rect 27244 24882 27300 24892
rect 27132 23996 27412 24052
rect 26908 23492 26964 23502
rect 27020 23492 27188 23548
rect 26908 23156 26964 23436
rect 27020 23156 27076 23166
rect 26908 23154 27076 23156
rect 26908 23102 27022 23154
rect 27074 23102 27076 23154
rect 26908 23100 27076 23102
rect 27020 23090 27076 23100
rect 26796 22430 26798 22482
rect 26850 22430 26852 22482
rect 26796 22418 26852 22430
rect 26460 21746 26516 21756
rect 26124 21634 26180 21644
rect 25564 21588 25620 21626
rect 25564 21522 25620 21532
rect 26908 21588 26964 21598
rect 25340 21474 25396 21486
rect 25340 21422 25342 21474
rect 25394 21422 25396 21474
rect 25340 21028 25396 21422
rect 25004 20972 25396 21028
rect 25788 21476 25844 21486
rect 25004 20802 25060 20972
rect 25004 20750 25006 20802
rect 25058 20750 25060 20802
rect 25004 20738 25060 20750
rect 25788 20690 25844 21420
rect 26236 21476 26292 21486
rect 26236 21382 26292 21420
rect 26572 21474 26628 21486
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 21364 26628 21422
rect 26572 21298 26628 21308
rect 26348 21252 26404 21262
rect 26348 20802 26404 21196
rect 26908 20804 26964 21532
rect 27020 20804 27076 20814
rect 26348 20750 26350 20802
rect 26402 20750 26404 20802
rect 26348 20738 26404 20750
rect 26572 20802 27076 20804
rect 26572 20750 27022 20802
rect 27074 20750 27076 20802
rect 26572 20748 27076 20750
rect 25788 20638 25790 20690
rect 25842 20638 25844 20690
rect 25788 20626 25844 20638
rect 25340 20132 25396 20142
rect 23436 18396 23828 18452
rect 23324 18340 23380 18396
rect 23324 18284 23492 18340
rect 23324 17556 23380 17566
rect 23212 17500 23324 17556
rect 23324 17462 23380 17500
rect 22876 16942 22878 16994
rect 22930 16942 22932 16994
rect 22876 16930 22932 16942
rect 22764 16716 23044 16772
rect 22988 16210 23044 16716
rect 22988 16158 22990 16210
rect 23042 16158 23044 16210
rect 22988 16146 23044 16158
rect 22428 16100 22484 16110
rect 23100 16100 23156 16110
rect 22428 16098 22708 16100
rect 22428 16046 22430 16098
rect 22482 16046 22708 16098
rect 22428 16044 22708 16046
rect 22428 16034 22484 16044
rect 22540 15540 22596 15550
rect 22540 15446 22596 15484
rect 21308 15092 21700 15148
rect 21420 14532 21476 14542
rect 20860 14530 21476 14532
rect 20860 14478 21422 14530
rect 21474 14478 21476 14530
rect 20860 14476 21476 14478
rect 21308 12962 21364 12974
rect 21308 12910 21310 12962
rect 21362 12910 21364 12962
rect 21308 12740 21364 12910
rect 20748 12738 21364 12740
rect 20748 12686 20750 12738
rect 20802 12686 21364 12738
rect 20748 12684 21364 12686
rect 20748 12674 20804 12684
rect 20524 10658 20580 10668
rect 17500 10612 17556 10622
rect 18396 10612 18452 10622
rect 17500 10610 17780 10612
rect 17500 10558 17502 10610
rect 17554 10558 17780 10610
rect 17500 10556 17780 10558
rect 17500 10546 17556 10556
rect 17724 9938 17780 10556
rect 18396 10518 18452 10556
rect 17724 9886 17726 9938
rect 17778 9886 17780 9938
rect 17724 9874 17780 9886
rect 18396 9714 18452 9726
rect 18396 9662 18398 9714
rect 18450 9662 18452 9714
rect 18172 9604 18228 9614
rect 18172 9510 18228 9548
rect 18284 9602 18340 9614
rect 18284 9550 18286 9602
rect 18338 9550 18340 9602
rect 16716 9090 16772 9100
rect 17388 9042 17444 9054
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 16604 7698 16660 7868
rect 16716 8930 16772 8942
rect 16716 8878 16718 8930
rect 16770 8878 16772 8930
rect 16716 7812 16772 8878
rect 16828 8818 16884 8830
rect 16828 8766 16830 8818
rect 16882 8766 16884 8818
rect 16828 8148 16884 8766
rect 16828 8082 16884 8092
rect 17388 8036 17444 8990
rect 18172 8932 18228 8942
rect 18172 8838 18228 8876
rect 17948 8260 18004 8270
rect 17388 7970 17444 7980
rect 17836 8204 17948 8260
rect 16716 7756 17108 7812
rect 16604 7646 16606 7698
rect 16658 7646 16660 7698
rect 16604 7634 16660 7646
rect 16828 7588 16884 7598
rect 16828 7494 16884 7532
rect 16492 7310 16494 7362
rect 16546 7310 16548 7362
rect 16492 7298 16548 7310
rect 16380 6638 16382 6690
rect 16434 6638 16436 6690
rect 16380 6626 16436 6638
rect 17052 6690 17108 7756
rect 17388 7476 17444 7486
rect 17388 7382 17444 7420
rect 17052 6638 17054 6690
rect 17106 6638 17108 6690
rect 17052 6626 17108 6638
rect 16716 6468 16772 6478
rect 16380 6356 16436 6366
rect 16380 6130 16436 6300
rect 16380 6078 16382 6130
rect 16434 6078 16436 6130
rect 16380 6066 16436 6078
rect 16156 5906 16212 5918
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 16156 5460 16212 5854
rect 16604 5908 16660 5918
rect 16492 5796 16548 5806
rect 16492 5702 16548 5740
rect 16156 5394 16212 5404
rect 16604 5348 16660 5852
rect 16716 5906 16772 6412
rect 16716 5854 16718 5906
rect 16770 5854 16772 5906
rect 16716 5572 16772 5854
rect 16940 6468 16996 6478
rect 16940 6020 16996 6412
rect 17724 6244 17780 6254
rect 17724 6130 17780 6188
rect 17724 6078 17726 6130
rect 17778 6078 17780 6130
rect 17724 6066 17780 6078
rect 16828 5572 16884 5582
rect 16716 5516 16828 5572
rect 16828 5506 16884 5516
rect 16604 5292 16884 5348
rect 15932 5070 15934 5122
rect 15986 5070 15988 5122
rect 15932 5058 15988 5070
rect 14700 4398 14702 4450
rect 14754 4398 14756 4450
rect 14700 4386 14756 4398
rect 15372 4898 15428 4910
rect 15372 4846 15374 4898
rect 15426 4846 15428 4898
rect 14588 3714 14644 3724
rect 13916 3614 13918 3666
rect 13970 3614 13972 3666
rect 13916 3602 13972 3614
rect 13132 3502 13134 3554
rect 13186 3502 13188 3554
rect 13132 3490 13188 3502
rect 13692 3444 13748 3454
rect 15372 3388 15428 4846
rect 16828 4226 16884 5292
rect 16940 5234 16996 5964
rect 16940 5182 16942 5234
rect 16994 5182 16996 5234
rect 16940 5170 16996 5182
rect 17052 5572 17108 5582
rect 16828 4174 16830 4226
rect 16882 4174 16884 4226
rect 16828 4162 16884 4174
rect 16044 3666 16100 3678
rect 16044 3614 16046 3666
rect 16098 3614 16100 3666
rect 16044 3556 16100 3614
rect 16044 3490 16100 3500
rect 13692 800 13748 3388
rect 15260 3332 15428 3388
rect 16940 3444 16996 3454
rect 17052 3444 17108 5516
rect 17276 5572 17332 5582
rect 16940 3442 17108 3444
rect 16940 3390 16942 3442
rect 16994 3390 17108 3442
rect 16940 3388 17108 3390
rect 17164 5348 17220 5358
rect 16940 3378 16996 3388
rect 15260 800 15316 3332
rect 17164 980 17220 5292
rect 17276 3554 17332 5516
rect 17724 4564 17780 4574
rect 17836 4564 17892 8204
rect 17948 8194 18004 8204
rect 18284 7252 18340 9550
rect 18396 7700 18452 9662
rect 20636 9714 20692 9726
rect 20636 9662 20638 9714
rect 20690 9662 20692 9714
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20300 8930 20356 8942
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 19740 8260 19796 8270
rect 19740 8166 19796 8204
rect 20300 8258 20356 8878
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 20188 8036 20244 8046
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 18396 7634 18452 7644
rect 19852 7700 19908 7710
rect 19628 7476 19684 7486
rect 18284 7186 18340 7196
rect 18508 7362 18564 7374
rect 18508 7310 18510 7362
rect 18562 7310 18564 7362
rect 18060 6132 18116 6142
rect 18060 6038 18116 6076
rect 18396 5908 18452 5918
rect 18396 5814 18452 5852
rect 18508 5348 18564 7310
rect 19068 7252 19124 7262
rect 18620 6244 18676 6254
rect 18620 6130 18676 6188
rect 18620 6078 18622 6130
rect 18674 6078 18676 6130
rect 18620 5460 18676 6078
rect 18844 5906 18900 5918
rect 18844 5854 18846 5906
rect 18898 5854 18900 5906
rect 18620 5394 18676 5404
rect 18732 5794 18788 5806
rect 18732 5742 18734 5794
rect 18786 5742 18788 5794
rect 18508 5282 18564 5292
rect 17724 4562 17892 4564
rect 17724 4510 17726 4562
rect 17778 4510 17892 4562
rect 17724 4508 17892 4510
rect 18060 5124 18116 5134
rect 17724 4498 17780 4508
rect 18060 4338 18116 5068
rect 18732 4452 18788 5742
rect 18844 5348 18900 5854
rect 18956 5906 19012 5918
rect 18956 5854 18958 5906
rect 19010 5854 19012 5906
rect 18956 5572 19012 5854
rect 18956 5506 19012 5516
rect 18844 5282 18900 5292
rect 19068 5234 19124 7196
rect 19180 6804 19236 6814
rect 19628 6804 19684 7420
rect 19180 6802 19684 6804
rect 19180 6750 19182 6802
rect 19234 6750 19684 6802
rect 19180 6748 19684 6750
rect 19180 6738 19236 6748
rect 19628 6690 19684 6748
rect 19852 6802 19908 7644
rect 19852 6750 19854 6802
rect 19906 6750 19908 6802
rect 19852 6738 19908 6750
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19628 6626 19684 6638
rect 20188 6692 20244 7980
rect 20300 7586 20356 8206
rect 20636 8930 20692 9662
rect 20636 8878 20638 8930
rect 20690 8878 20692 8930
rect 20636 8258 20692 8878
rect 20748 9602 20804 9614
rect 20748 9550 20750 9602
rect 20802 9550 20804 9602
rect 20748 8372 20804 9550
rect 20748 8306 20804 8316
rect 20636 8206 20638 8258
rect 20690 8206 20692 8258
rect 20636 8194 20692 8206
rect 20860 8260 20916 12684
rect 21084 12516 21140 12526
rect 21084 12402 21140 12460
rect 21084 12350 21086 12402
rect 21138 12350 21140 12402
rect 21084 12338 21140 12350
rect 21420 12178 21476 14476
rect 21644 14420 21700 15092
rect 21420 12126 21422 12178
rect 21474 12126 21476 12178
rect 21420 12114 21476 12126
rect 21532 14418 21700 14420
rect 21532 14366 21646 14418
rect 21698 14366 21700 14418
rect 21532 14364 21700 14366
rect 21196 11844 21252 11854
rect 21196 10498 21252 11788
rect 21532 11508 21588 14364
rect 21644 14354 21700 14364
rect 21868 15092 22036 15148
rect 22092 15202 22148 15214
rect 22092 15150 22094 15202
rect 22146 15150 22148 15202
rect 21420 11452 21588 11508
rect 21644 13860 21700 13870
rect 21644 12402 21700 13804
rect 21644 12350 21646 12402
rect 21698 12350 21700 12402
rect 21196 10446 21198 10498
rect 21250 10446 21252 10498
rect 21196 10434 21252 10446
rect 21308 11170 21364 11182
rect 21308 11118 21310 11170
rect 21362 11118 21364 11170
rect 21308 9940 21364 11118
rect 21308 9874 21364 9884
rect 21420 9268 21476 11452
rect 21644 11396 21700 12350
rect 21868 11844 21924 15092
rect 22092 14420 22148 15150
rect 22540 14756 22596 14766
rect 22092 13524 22148 14364
rect 22316 14754 22596 14756
rect 22316 14702 22542 14754
rect 22594 14702 22596 14754
rect 22316 14700 22596 14702
rect 22204 14308 22260 14318
rect 22204 14214 22260 14252
rect 22204 13860 22260 13870
rect 22316 13860 22372 14700
rect 22540 14690 22596 14700
rect 22204 13858 22372 13860
rect 22204 13806 22206 13858
rect 22258 13806 22372 13858
rect 22204 13804 22372 13806
rect 22428 14418 22484 14430
rect 22428 14366 22430 14418
rect 22482 14366 22484 14418
rect 22204 13794 22260 13804
rect 22092 13458 22148 13468
rect 22428 13076 22484 14366
rect 22540 14308 22596 14318
rect 22540 14214 22596 14252
rect 21980 13020 22484 13076
rect 22540 13524 22596 13534
rect 21980 12290 22036 13020
rect 21980 12238 21982 12290
rect 22034 12238 22036 12290
rect 21980 12226 22036 12238
rect 22428 12516 22484 12526
rect 22428 12178 22484 12460
rect 22428 12126 22430 12178
rect 22482 12126 22484 12178
rect 22428 12114 22484 12126
rect 21868 11778 21924 11788
rect 21420 9202 21476 9212
rect 21532 11394 21700 11396
rect 21532 11342 21646 11394
rect 21698 11342 21700 11394
rect 21532 11340 21700 11342
rect 20860 8194 20916 8204
rect 21420 8260 21476 8270
rect 20748 8148 20804 8158
rect 20300 7534 20302 7586
rect 20354 7534 20356 7586
rect 20300 7522 20356 7534
rect 20412 8034 20468 8046
rect 20412 7982 20414 8034
rect 20466 7982 20468 8034
rect 20412 7588 20468 7982
rect 20412 7522 20468 7532
rect 20524 8034 20580 8046
rect 20524 7982 20526 8034
rect 20578 7982 20580 8034
rect 20524 7474 20580 7982
rect 20636 7700 20692 7710
rect 20748 7700 20804 8092
rect 20636 7698 20804 7700
rect 20636 7646 20638 7698
rect 20690 7646 20804 7698
rect 20636 7644 20804 7646
rect 20972 8148 21028 8158
rect 20636 7634 20692 7644
rect 20524 7422 20526 7474
rect 20578 7422 20580 7474
rect 20188 6690 20468 6692
rect 20188 6638 20190 6690
rect 20242 6638 20468 6690
rect 20188 6636 20468 6638
rect 20188 6626 20244 6636
rect 19740 6468 19796 6478
rect 19628 6466 19796 6468
rect 19628 6414 19742 6466
rect 19794 6414 19796 6466
rect 19628 6412 19796 6414
rect 19628 6132 19684 6412
rect 19740 6402 19796 6412
rect 19964 6468 20020 6506
rect 19964 6402 20020 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19628 6066 19684 6076
rect 19068 5182 19070 5234
rect 19122 5182 19124 5234
rect 19068 5170 19124 5182
rect 19852 5124 19908 5134
rect 19852 5030 19908 5068
rect 20412 5010 20468 6636
rect 20524 6132 20580 7422
rect 20748 7476 20804 7486
rect 20748 7382 20804 7420
rect 20972 7474 21028 8092
rect 20972 7422 20974 7474
rect 21026 7422 21028 7474
rect 20972 7410 21028 7422
rect 21420 8034 21476 8204
rect 21420 7982 21422 8034
rect 21474 7982 21476 8034
rect 21420 7140 21476 7982
rect 21532 7924 21588 11340
rect 21644 11330 21700 11340
rect 21756 11396 21812 11406
rect 21644 10612 21700 10622
rect 21756 10612 21812 11340
rect 22428 11172 22484 11182
rect 22540 11172 22596 13468
rect 22428 11170 22596 11172
rect 22428 11118 22430 11170
rect 22482 11118 22596 11170
rect 22428 11116 22596 11118
rect 22428 11060 22484 11116
rect 21700 10556 21812 10612
rect 22204 11004 22484 11060
rect 21644 10518 21700 10556
rect 21532 7858 21588 7868
rect 21644 9826 21700 9838
rect 21644 9774 21646 9826
rect 21698 9774 21700 9826
rect 21644 7588 21700 9774
rect 22204 9602 22260 11004
rect 22652 10612 22708 16044
rect 23100 14530 23156 16044
rect 23436 15092 23492 18284
rect 23772 17666 23828 18396
rect 24388 18396 24500 18452
rect 24556 19908 24612 19918
rect 24332 18358 24388 18396
rect 23884 18338 23940 18350
rect 23884 18286 23886 18338
rect 23938 18286 23940 18338
rect 23884 18228 23940 18286
rect 24220 18228 24276 18238
rect 23884 18172 24220 18228
rect 23772 17614 23774 17666
rect 23826 17614 23828 17666
rect 23660 16884 23716 16894
rect 23772 16884 23828 17614
rect 23660 16882 23940 16884
rect 23660 16830 23662 16882
rect 23714 16830 23940 16882
rect 23660 16828 23940 16830
rect 23660 16818 23716 16828
rect 23884 16100 23940 16828
rect 23884 16006 23940 16044
rect 24108 16770 24164 16782
rect 24108 16718 24110 16770
rect 24162 16718 24164 16770
rect 24108 15316 24164 16718
rect 23436 15026 23492 15036
rect 23772 15204 23828 15214
rect 24108 15148 24164 15260
rect 23772 14642 23828 15148
rect 23772 14590 23774 14642
rect 23826 14590 23828 14642
rect 23772 14578 23828 14590
rect 23884 15092 24164 15148
rect 24220 15148 24276 18172
rect 24556 17778 24612 19852
rect 24556 17726 24558 17778
rect 24610 17726 24612 17778
rect 24556 17714 24612 17726
rect 24668 19906 24724 19918
rect 24668 19854 24670 19906
rect 24722 19854 24724 19906
rect 24668 19234 24724 19854
rect 25340 19348 25396 20076
rect 25340 19254 25396 19292
rect 26012 20132 26068 20142
rect 26012 19906 26068 20076
rect 26012 19854 26014 19906
rect 26066 19854 26068 19906
rect 24668 19182 24670 19234
rect 24722 19182 24724 19234
rect 24668 17780 24724 19182
rect 24668 17714 24724 17724
rect 25228 18562 25284 18574
rect 25228 18510 25230 18562
rect 25282 18510 25284 18562
rect 24668 17108 24724 17118
rect 24668 17014 24724 17052
rect 25228 16996 25284 18510
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 25452 17108 25508 18398
rect 26012 18228 26068 19854
rect 26460 20020 26516 20030
rect 26572 20020 26628 20748
rect 27020 20738 27076 20748
rect 27132 20244 27188 23492
rect 27356 23378 27412 23996
rect 27580 23604 27636 23614
rect 27636 23548 27748 23604
rect 27580 23538 27636 23548
rect 27356 23326 27358 23378
rect 27410 23326 27412 23378
rect 27356 23314 27412 23326
rect 27468 23492 27524 23502
rect 27468 23378 27524 23436
rect 27468 23326 27470 23378
rect 27522 23326 27524 23378
rect 27468 23314 27524 23326
rect 27580 23380 27636 23390
rect 27244 23156 27300 23166
rect 27244 22594 27300 23100
rect 27244 22542 27246 22594
rect 27298 22542 27300 22594
rect 27244 22530 27300 22542
rect 27580 22594 27636 23324
rect 27580 22542 27582 22594
rect 27634 22542 27636 22594
rect 27580 22530 27636 22542
rect 27692 22372 27748 23548
rect 27804 22596 27860 27804
rect 27916 27298 27972 28364
rect 27916 27246 27918 27298
rect 27970 27246 27972 27298
rect 27916 27234 27972 27246
rect 28140 28196 28196 28206
rect 28140 27300 28196 28140
rect 28252 27970 28308 28364
rect 28364 28084 28420 29036
rect 28476 28980 28532 30158
rect 28476 28924 28644 28980
rect 28476 28756 28532 28766
rect 28476 28662 28532 28700
rect 28588 28532 28644 28924
rect 28476 28476 28644 28532
rect 28476 28196 28532 28476
rect 28476 28130 28532 28140
rect 28364 28018 28420 28028
rect 28252 27918 28254 27970
rect 28306 27918 28308 27970
rect 28252 27906 28308 27918
rect 28700 27860 28756 27870
rect 28364 27858 28756 27860
rect 28364 27806 28702 27858
rect 28754 27806 28756 27858
rect 28364 27804 28756 27806
rect 28252 27300 28308 27310
rect 28140 27298 28308 27300
rect 28140 27246 28254 27298
rect 28306 27246 28308 27298
rect 28140 27244 28308 27246
rect 28252 27234 28308 27244
rect 28364 27076 28420 27804
rect 28700 27794 28756 27804
rect 28700 27524 28756 27534
rect 28364 26516 28420 27020
rect 28476 27300 28532 27310
rect 28476 26740 28532 27244
rect 28476 26684 28644 26740
rect 28476 26516 28532 26526
rect 28364 26514 28532 26516
rect 28364 26462 28478 26514
rect 28530 26462 28532 26514
rect 28364 26460 28532 26462
rect 28476 26450 28532 26460
rect 28588 26292 28644 26684
rect 28476 26236 28644 26292
rect 28364 24948 28420 24958
rect 28364 24834 28420 24892
rect 28364 24782 28366 24834
rect 28418 24782 28420 24834
rect 28364 24770 28420 24782
rect 28140 23380 28196 23390
rect 28140 23286 28196 23324
rect 28476 23156 28532 26236
rect 28700 23716 28756 27468
rect 28588 23660 28756 23716
rect 28588 23268 28644 23660
rect 28700 23492 28756 23502
rect 28700 23378 28756 23436
rect 28700 23326 28702 23378
rect 28754 23326 28756 23378
rect 28700 23314 28756 23326
rect 28812 23380 28868 31052
rect 29596 31042 29652 31052
rect 28924 30994 28980 31006
rect 28924 30942 28926 30994
rect 28978 30942 28980 30994
rect 28924 29204 28980 30942
rect 29260 30324 29316 30334
rect 29148 29204 29204 29214
rect 28924 29148 29148 29204
rect 29148 28642 29204 29148
rect 29148 28590 29150 28642
rect 29202 28590 29204 28642
rect 29148 28578 29204 28590
rect 29260 28644 29316 30268
rect 29596 30100 29652 30110
rect 29260 28532 29316 28588
rect 29484 29986 29540 29998
rect 29484 29934 29486 29986
rect 29538 29934 29540 29986
rect 29484 29876 29540 29934
rect 29484 28644 29540 29820
rect 29596 28756 29652 30044
rect 29596 28690 29652 28700
rect 29932 29988 29988 29998
rect 29932 28754 29988 29932
rect 29932 28702 29934 28754
rect 29986 28702 29988 28754
rect 29932 28690 29988 28702
rect 29484 28578 29540 28588
rect 29260 28476 29428 28532
rect 29148 28420 29204 28430
rect 28924 27972 28980 27982
rect 28924 25620 28980 27916
rect 29148 27748 29204 28364
rect 29148 27682 29204 27692
rect 29260 28084 29316 28094
rect 29260 27300 29316 28028
rect 29372 27972 29428 28476
rect 29932 28420 29988 28430
rect 29820 28364 29932 28420
rect 29708 27972 29764 27982
rect 29372 27970 29764 27972
rect 29372 27918 29710 27970
rect 29762 27918 29764 27970
rect 29372 27916 29764 27918
rect 29708 27906 29764 27916
rect 29260 27186 29316 27244
rect 29484 27748 29540 27758
rect 29820 27748 29876 28364
rect 29932 28354 29988 28364
rect 29484 27298 29540 27692
rect 29484 27246 29486 27298
rect 29538 27246 29540 27298
rect 29484 27234 29540 27246
rect 29708 27692 29876 27748
rect 29260 27134 29262 27186
rect 29314 27134 29316 27186
rect 29260 26908 29316 27134
rect 29260 26852 29428 26908
rect 29372 25732 29428 26852
rect 29596 26290 29652 26302
rect 29596 26238 29598 26290
rect 29650 26238 29652 26290
rect 29484 25732 29540 25742
rect 29372 25730 29540 25732
rect 29372 25678 29486 25730
rect 29538 25678 29540 25730
rect 29372 25676 29540 25678
rect 29484 25666 29540 25676
rect 28924 25554 28980 25564
rect 29148 25284 29204 25294
rect 29148 25190 29204 25228
rect 29148 24724 29204 24734
rect 29596 24724 29652 26238
rect 29708 25620 29764 27692
rect 29820 27300 29876 27310
rect 30044 27300 30100 32284
rect 30156 32246 30212 32284
rect 30940 32340 30996 32508
rect 30940 32274 30996 32284
rect 31052 32564 31108 33292
rect 31164 33236 31220 33246
rect 31276 33236 31332 35420
rect 31220 33180 31332 33236
rect 31164 33142 31220 33180
rect 31388 33012 31444 35980
rect 31500 35308 31556 36316
rect 31500 35252 31668 35308
rect 31500 33684 31556 33694
rect 31500 33346 31556 33628
rect 31500 33294 31502 33346
rect 31554 33294 31556 33346
rect 31500 33282 31556 33294
rect 31612 33348 31668 35252
rect 31612 33282 31668 33292
rect 31164 32956 31444 33012
rect 31164 32676 31220 32956
rect 31276 32788 31332 32798
rect 31724 32788 31780 36652
rect 32060 36148 32116 36158
rect 31836 35698 31892 35710
rect 31836 35646 31838 35698
rect 31890 35646 31892 35698
rect 31836 34132 31892 35646
rect 32060 35698 32116 36092
rect 32172 35922 32228 36876
rect 32172 35870 32174 35922
rect 32226 35870 32228 35922
rect 32172 35858 32228 35870
rect 32284 35924 32340 37660
rect 32620 37492 32676 40908
rect 32844 40898 32900 40908
rect 33180 40628 33236 40638
rect 33852 40628 33908 41132
rect 34188 40964 34244 40974
rect 34188 40870 34244 40908
rect 34300 40740 34356 42700
rect 34412 42644 34468 42654
rect 34412 42550 34468 42588
rect 34636 42642 34692 42700
rect 34636 42590 34638 42642
rect 34690 42590 34692 42642
rect 34636 42578 34692 42590
rect 33180 40534 33236 40572
rect 33740 40626 33908 40628
rect 33740 40574 33854 40626
rect 33906 40574 33908 40626
rect 33740 40572 33908 40574
rect 33180 40404 33236 40414
rect 33404 40404 33460 40414
rect 33236 40402 33460 40404
rect 33236 40350 33406 40402
rect 33458 40350 33460 40402
rect 33236 40348 33460 40350
rect 33180 40338 33236 40348
rect 33068 40180 33124 40190
rect 32844 40178 33124 40180
rect 32844 40126 33070 40178
rect 33122 40126 33124 40178
rect 32844 40124 33124 40126
rect 32732 39620 32788 39630
rect 32844 39620 32900 40124
rect 33068 40114 33124 40124
rect 32732 39618 32900 39620
rect 32732 39566 32734 39618
rect 32786 39566 32900 39618
rect 32732 39564 32900 39566
rect 32956 39732 33012 39742
rect 32732 39508 32788 39564
rect 32732 39442 32788 39452
rect 32956 39060 33012 39676
rect 33068 39620 33124 39630
rect 33068 39526 33124 39564
rect 33180 39508 33236 39518
rect 33180 39414 33236 39452
rect 33068 39060 33124 39070
rect 32956 39058 33124 39060
rect 32956 39006 33070 39058
rect 33122 39006 33124 39058
rect 32956 39004 33124 39006
rect 33068 38994 33124 39004
rect 33180 38722 33236 38734
rect 33180 38670 33182 38722
rect 33234 38670 33236 38722
rect 33180 38668 33236 38670
rect 33180 38612 33348 38668
rect 32732 38164 32788 38174
rect 32732 38050 32788 38108
rect 32732 37998 32734 38050
rect 32786 37998 32788 38050
rect 32732 37986 32788 37998
rect 33180 37828 33236 37838
rect 32620 37426 32676 37436
rect 33068 37826 33236 37828
rect 33068 37774 33182 37826
rect 33234 37774 33236 37826
rect 33068 37772 33236 37774
rect 32396 37156 32452 37166
rect 32396 37062 32452 37100
rect 32508 37044 32564 37054
rect 32956 37044 33012 37054
rect 32508 37042 32788 37044
rect 32508 36990 32510 37042
rect 32562 36990 32788 37042
rect 32508 36988 32788 36990
rect 32508 36978 32564 36988
rect 32508 36596 32564 36606
rect 32284 35868 32452 35924
rect 32060 35646 32062 35698
rect 32114 35646 32116 35698
rect 32060 35634 32116 35646
rect 32284 35698 32340 35710
rect 32284 35646 32286 35698
rect 32338 35646 32340 35698
rect 32172 35588 32228 35598
rect 31836 34038 31892 34076
rect 32060 35252 32116 35262
rect 32060 34130 32116 35196
rect 32172 34354 32228 35532
rect 32172 34302 32174 34354
rect 32226 34302 32228 34354
rect 32172 34290 32228 34302
rect 32060 34078 32062 34130
rect 32114 34078 32116 34130
rect 32060 33908 32116 34078
rect 32060 33842 32116 33852
rect 32284 34244 32340 35646
rect 32396 35252 32452 35868
rect 32508 35810 32564 36540
rect 32508 35758 32510 35810
rect 32562 35758 32564 35810
rect 32508 35746 32564 35758
rect 32620 36036 32676 36046
rect 32396 35186 32452 35196
rect 32508 35476 32564 35486
rect 32284 34130 32340 34188
rect 32508 34242 32564 35420
rect 32508 34190 32510 34242
rect 32562 34190 32564 34242
rect 32508 34178 32564 34190
rect 32284 34078 32286 34130
rect 32338 34078 32340 34130
rect 31948 33572 32004 33582
rect 31948 33346 32004 33516
rect 31948 33294 31950 33346
rect 32002 33294 32004 33346
rect 31948 33282 32004 33294
rect 31276 32694 31332 32732
rect 31500 32732 31780 32788
rect 31948 32788 32004 32798
rect 32284 32788 32340 34078
rect 31948 32786 32340 32788
rect 31948 32734 31950 32786
rect 32002 32734 32340 32786
rect 31948 32732 32340 32734
rect 32396 34132 32452 34142
rect 32396 32788 32452 34076
rect 31164 32610 31220 32620
rect 30380 31892 30436 31902
rect 30380 31666 30436 31836
rect 31052 31890 31108 32508
rect 31052 31838 31054 31890
rect 31106 31838 31108 31890
rect 31052 31826 31108 31838
rect 30380 31614 30382 31666
rect 30434 31614 30436 31666
rect 30156 30884 30212 30894
rect 30156 30210 30212 30828
rect 30380 30324 30436 31614
rect 30716 31666 30772 31678
rect 30716 31614 30718 31666
rect 30770 31614 30772 31666
rect 30716 30884 30772 31614
rect 30716 30818 30772 30828
rect 30828 31444 30884 31454
rect 30828 30434 30884 31388
rect 30828 30382 30830 30434
rect 30882 30382 30884 30434
rect 30828 30370 30884 30382
rect 30380 30258 30436 30268
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 30156 30146 30212 30158
rect 31388 30212 31444 30222
rect 30268 30100 30324 30110
rect 30268 30006 30324 30044
rect 30380 30098 30436 30110
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 29820 27298 30100 27300
rect 29820 27246 29822 27298
rect 29874 27246 30100 27298
rect 29820 27244 30100 27246
rect 30156 29876 30212 29886
rect 30156 29540 30212 29820
rect 29820 27234 29876 27244
rect 30156 27186 30212 29484
rect 30380 28532 30436 30046
rect 31276 29988 31332 29998
rect 31052 29876 31108 29886
rect 30716 29652 30772 29662
rect 30604 29596 30716 29652
rect 30492 29540 30548 29550
rect 30492 29426 30548 29484
rect 30492 29374 30494 29426
rect 30546 29374 30548 29426
rect 30492 29362 30548 29374
rect 30156 27134 30158 27186
rect 30210 27134 30212 27186
rect 30156 27122 30212 27134
rect 30268 28476 30436 28532
rect 30268 26852 30324 28476
rect 30380 27300 30436 27310
rect 30380 27206 30436 27244
rect 30604 26908 30660 29596
rect 30716 29586 30772 29596
rect 31052 29426 31108 29820
rect 31276 29652 31332 29932
rect 31276 29586 31332 29596
rect 31388 29650 31444 30156
rect 31500 29764 31556 32732
rect 31948 32722 32004 32732
rect 31836 32676 31892 32686
rect 31612 32564 31668 32574
rect 31612 32452 31668 32508
rect 31724 32562 31780 32574
rect 31724 32510 31726 32562
rect 31778 32510 31780 32562
rect 31724 32452 31780 32510
rect 31612 32396 31780 32452
rect 31724 32116 31780 32126
rect 31836 32116 31892 32620
rect 32172 32562 32228 32574
rect 32172 32510 32174 32562
rect 32226 32510 32228 32562
rect 32172 32452 32228 32510
rect 32172 32386 32228 32396
rect 32284 32564 32340 32574
rect 32284 32450 32340 32508
rect 32396 32562 32452 32732
rect 32396 32510 32398 32562
rect 32450 32510 32452 32562
rect 32396 32498 32452 32510
rect 32284 32398 32286 32450
rect 32338 32398 32340 32450
rect 32284 32386 32340 32398
rect 32620 32452 32676 35980
rect 32732 33458 32788 36988
rect 32956 34356 33012 36988
rect 33068 36484 33124 37772
rect 33180 37762 33236 37772
rect 33292 37604 33348 38612
rect 33292 37538 33348 37548
rect 33068 36418 33124 36428
rect 33180 37156 33236 37166
rect 33068 35698 33124 35710
rect 33068 35646 33070 35698
rect 33122 35646 33124 35698
rect 33068 35364 33124 35646
rect 33180 35588 33236 37100
rect 33292 37154 33348 37166
rect 33292 37102 33294 37154
rect 33346 37102 33348 37154
rect 33292 36036 33348 37102
rect 33292 35970 33348 35980
rect 33404 35700 33460 40348
rect 33628 40178 33684 40190
rect 33628 40126 33630 40178
rect 33682 40126 33684 40178
rect 33516 39732 33572 39742
rect 33516 39618 33572 39676
rect 33516 39566 33518 39618
rect 33570 39566 33572 39618
rect 33516 39554 33572 39566
rect 33628 39508 33684 40126
rect 33628 39414 33684 39452
rect 33628 39060 33684 39070
rect 33628 38966 33684 39004
rect 33516 37828 33572 37838
rect 33516 37734 33572 37772
rect 33740 37380 33796 40572
rect 33852 40562 33908 40572
rect 34188 40684 34356 40740
rect 34748 42532 34804 42542
rect 34748 40962 34804 42476
rect 34860 41188 34916 42924
rect 35308 42980 35364 42990
rect 35532 42980 35588 44156
rect 35868 44100 35924 44110
rect 35308 42978 35588 42980
rect 35308 42926 35310 42978
rect 35362 42926 35588 42978
rect 35308 42924 35588 42926
rect 35644 43428 35700 43438
rect 35644 42978 35700 43372
rect 35644 42926 35646 42978
rect 35698 42926 35700 42978
rect 35308 42914 35364 42924
rect 35644 42914 35700 42926
rect 35868 42868 35924 44044
rect 36428 43876 36484 44270
rect 40124 44322 40180 44334
rect 40124 44270 40126 44322
rect 40178 44270 40180 44322
rect 37100 44212 37156 44222
rect 37100 44118 37156 44156
rect 39228 43988 39284 43998
rect 36428 43810 36484 43820
rect 37324 43876 37380 43886
rect 35980 43596 36148 43652
rect 35980 43538 36036 43596
rect 35980 43486 35982 43538
rect 36034 43486 36036 43538
rect 35980 43474 36036 43486
rect 36092 43540 36148 43596
rect 36428 43540 36484 43550
rect 36092 43538 36596 43540
rect 36092 43486 36430 43538
rect 36482 43486 36596 43538
rect 36092 43484 36596 43486
rect 36428 43474 36484 43484
rect 36316 43092 36372 43102
rect 35868 42812 36036 42868
rect 35644 42756 35700 42766
rect 35644 42754 35812 42756
rect 35644 42702 35646 42754
rect 35698 42702 35812 42754
rect 35644 42700 35812 42702
rect 35644 42690 35700 42700
rect 34972 42530 35028 42542
rect 34972 42478 34974 42530
rect 35026 42478 35028 42530
rect 34972 41748 35028 42478
rect 35532 42308 35588 42318
rect 35196 41860 35252 41870
rect 35196 41766 35252 41804
rect 34972 41300 35028 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35308 41412 35364 41422
rect 35532 41412 35588 42252
rect 35308 41410 35588 41412
rect 35308 41358 35310 41410
rect 35362 41358 35588 41410
rect 35308 41356 35588 41358
rect 35644 42084 35700 42094
rect 35644 41410 35700 42028
rect 35644 41358 35646 41410
rect 35698 41358 35700 41410
rect 35308 41346 35364 41356
rect 35644 41346 35700 41358
rect 35084 41300 35140 41310
rect 34972 41298 35140 41300
rect 34972 41246 35086 41298
rect 35138 41246 35140 41298
rect 34972 41244 35140 41246
rect 35084 41234 35140 41244
rect 34860 41132 35028 41188
rect 34748 40910 34750 40962
rect 34802 40910 34804 40962
rect 34188 40178 34244 40684
rect 34300 40404 34356 40414
rect 34300 40310 34356 40348
rect 34188 40126 34190 40178
rect 34242 40126 34244 40178
rect 33964 39956 34020 39966
rect 33964 39844 34020 39900
rect 34076 39844 34132 39854
rect 33964 39842 34132 39844
rect 33964 39790 34078 39842
rect 34130 39790 34132 39842
rect 33964 39788 34132 39790
rect 34076 39778 34132 39788
rect 34188 39730 34244 40126
rect 34188 39678 34190 39730
rect 34242 39678 34244 39730
rect 34188 39666 34244 39678
rect 33852 39394 33908 39406
rect 34636 39396 34692 39406
rect 33852 39342 33854 39394
rect 33906 39342 33908 39394
rect 33852 39284 33908 39342
rect 33852 39218 33908 39228
rect 34300 39394 34692 39396
rect 34300 39342 34638 39394
rect 34690 39342 34692 39394
rect 34300 39340 34692 39342
rect 34188 39172 34244 39182
rect 33852 38836 33908 38846
rect 33852 38742 33908 38780
rect 34188 38276 34244 39116
rect 34300 38946 34356 39340
rect 34636 39330 34692 39340
rect 34300 38894 34302 38946
rect 34354 38894 34356 38946
rect 34300 38724 34356 38894
rect 34412 38836 34468 38846
rect 34636 38836 34692 38874
rect 34412 38742 34468 38780
rect 34524 38780 34636 38836
rect 34300 38658 34356 38668
rect 34188 38220 34468 38276
rect 34412 38050 34468 38220
rect 34524 38162 34580 38780
rect 34636 38770 34692 38780
rect 34524 38110 34526 38162
rect 34578 38110 34580 38162
rect 34524 38098 34580 38110
rect 34636 38500 34692 38510
rect 34412 37998 34414 38050
rect 34466 37998 34468 38050
rect 34412 37986 34468 37998
rect 33964 37940 34020 37950
rect 33964 37846 34020 37884
rect 34188 37826 34244 37838
rect 34188 37774 34190 37826
rect 34242 37774 34244 37826
rect 33628 37324 33796 37380
rect 33852 37604 33908 37614
rect 34188 37604 34244 37774
rect 33908 37548 34244 37604
rect 34524 37828 34580 37838
rect 34636 37828 34692 38444
rect 34524 37826 34692 37828
rect 34524 37774 34526 37826
rect 34578 37774 34692 37826
rect 34524 37772 34692 37774
rect 33628 36932 33684 37324
rect 33516 36876 33684 36932
rect 33740 37154 33796 37166
rect 33740 37102 33742 37154
rect 33794 37102 33796 37154
rect 33516 36148 33572 36876
rect 33628 36596 33684 36606
rect 33628 36502 33684 36540
rect 33516 36082 33572 36092
rect 33404 35644 33572 35700
rect 33180 35532 33460 35588
rect 33068 35298 33124 35308
rect 33292 34356 33348 34366
rect 32956 34354 33348 34356
rect 32956 34302 33294 34354
rect 33346 34302 33348 34354
rect 32956 34300 33348 34302
rect 33292 34290 33348 34300
rect 33404 34354 33460 35532
rect 33516 35252 33572 35644
rect 33516 35196 33684 35252
rect 33404 34302 33406 34354
rect 33458 34302 33460 34354
rect 33404 34290 33460 34302
rect 33516 34244 33572 34254
rect 33516 34150 33572 34188
rect 32844 34132 32900 34142
rect 33068 34132 33124 34142
rect 32900 34130 33124 34132
rect 32900 34078 33070 34130
rect 33122 34078 33124 34130
rect 32900 34076 33124 34078
rect 32844 34066 32900 34076
rect 33068 34066 33124 34076
rect 33628 34132 33684 35196
rect 33628 34038 33684 34076
rect 32732 33406 32734 33458
rect 32786 33406 32788 33458
rect 32732 33394 32788 33406
rect 33180 33572 33236 33582
rect 32620 32386 32676 32396
rect 31780 32060 31892 32116
rect 31724 32050 31780 32060
rect 31724 30884 31780 30894
rect 31724 30790 31780 30828
rect 31836 30210 31892 32060
rect 33068 32338 33124 32350
rect 33068 32286 33070 32338
rect 33122 32286 33124 32338
rect 33068 31332 33124 32286
rect 33180 31890 33236 33516
rect 33740 33236 33796 37102
rect 33852 36596 33908 37548
rect 34524 37380 34580 37772
rect 34188 37324 34580 37380
rect 34076 37154 34132 37166
rect 34076 37102 34078 37154
rect 34130 37102 34132 37154
rect 33852 36530 33908 36540
rect 33964 37042 34020 37054
rect 33964 36990 33966 37042
rect 34018 36990 34020 37042
rect 33852 35812 33908 35822
rect 33964 35812 34020 36990
rect 33852 35810 34020 35812
rect 33852 35758 33854 35810
rect 33906 35758 34020 35810
rect 33852 35756 34020 35758
rect 33852 35746 33908 35756
rect 34076 35588 34132 37102
rect 34076 35522 34132 35532
rect 34188 35476 34244 37324
rect 34524 37154 34580 37166
rect 34524 37102 34526 37154
rect 34578 37102 34580 37154
rect 34524 37044 34580 37102
rect 34524 36978 34580 36988
rect 34412 36372 34468 36382
rect 34412 36370 34580 36372
rect 34412 36318 34414 36370
rect 34466 36318 34580 36370
rect 34412 36316 34580 36318
rect 34412 36306 34468 36316
rect 34188 35410 34244 35420
rect 34300 36258 34356 36270
rect 34300 36206 34302 36258
rect 34354 36206 34356 36258
rect 34076 34244 34132 34254
rect 34076 34150 34132 34188
rect 34188 34020 34244 34030
rect 34188 33460 34244 33964
rect 34300 33572 34356 36206
rect 34412 34130 34468 34142
rect 34412 34078 34414 34130
rect 34466 34078 34468 34130
rect 34412 33684 34468 34078
rect 34412 33618 34468 33628
rect 34300 33506 34356 33516
rect 34188 33394 34244 33404
rect 34300 33236 34356 33246
rect 33404 33180 34244 33236
rect 33404 32900 33460 33180
rect 33404 32562 33460 32844
rect 33740 32676 33796 32686
rect 33404 32510 33406 32562
rect 33458 32510 33460 32562
rect 33404 32498 33460 32510
rect 33628 32674 33796 32676
rect 33628 32622 33742 32674
rect 33794 32622 33796 32674
rect 33628 32620 33796 32622
rect 33404 32338 33460 32350
rect 33404 32286 33406 32338
rect 33458 32286 33460 32338
rect 33404 32004 33460 32286
rect 33404 31938 33460 31948
rect 33180 31838 33182 31890
rect 33234 31838 33236 31890
rect 33180 31826 33236 31838
rect 33068 31276 33460 31332
rect 33292 31106 33348 31118
rect 33292 31054 33294 31106
rect 33346 31054 33348 31106
rect 32396 30996 32452 31006
rect 32396 30994 32564 30996
rect 32396 30942 32398 30994
rect 32450 30942 32564 30994
rect 32396 30940 32564 30942
rect 32396 30930 32452 30940
rect 32172 30882 32228 30894
rect 32172 30830 32174 30882
rect 32226 30830 32228 30882
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 31836 30146 31892 30158
rect 32060 30770 32116 30782
rect 32060 30718 32062 30770
rect 32114 30718 32116 30770
rect 31500 29708 31780 29764
rect 31388 29598 31390 29650
rect 31442 29598 31444 29650
rect 31388 29586 31444 29598
rect 31612 29540 31668 29550
rect 31052 29374 31054 29426
rect 31106 29374 31108 29426
rect 31052 29362 31108 29374
rect 31500 29484 31612 29540
rect 30828 29314 30884 29326
rect 30828 29262 30830 29314
rect 30882 29262 30884 29314
rect 30828 28868 30884 29262
rect 30828 28802 30884 28812
rect 30940 28644 30996 28654
rect 30940 27858 30996 28588
rect 30940 27806 30942 27858
rect 30994 27806 30996 27858
rect 30940 27794 30996 27806
rect 30716 27300 30772 27310
rect 30716 27298 31444 27300
rect 30716 27246 30718 27298
rect 30770 27246 31444 27298
rect 30716 27244 31444 27246
rect 30716 27234 30772 27244
rect 31164 26962 31220 26974
rect 31164 26910 31166 26962
rect 31218 26910 31220 26962
rect 30604 26852 30772 26908
rect 30268 26628 30324 26796
rect 30156 26572 30324 26628
rect 30156 26180 30212 26572
rect 30268 26404 30324 26414
rect 30268 26310 30324 26348
rect 30156 26124 30324 26180
rect 29708 25618 29876 25620
rect 29708 25566 29710 25618
rect 29762 25566 29876 25618
rect 29708 25564 29876 25566
rect 29708 25554 29764 25564
rect 29708 24724 29764 24734
rect 29148 24722 29764 24724
rect 29148 24670 29150 24722
rect 29202 24670 29710 24722
rect 29762 24670 29764 24722
rect 29148 24668 29764 24670
rect 29148 24658 29204 24668
rect 29484 24164 29540 24174
rect 29484 24070 29540 24108
rect 29708 24164 29764 24668
rect 29708 24098 29764 24108
rect 29820 24052 29876 25564
rect 30268 24162 30324 26124
rect 30716 25844 30772 26852
rect 31052 26850 31108 26862
rect 31052 26798 31054 26850
rect 31106 26798 31108 26850
rect 30828 26404 30884 26414
rect 31052 26404 31108 26798
rect 30884 26348 31108 26404
rect 30828 26338 30884 26348
rect 31164 26068 31220 26910
rect 31164 26002 31220 26012
rect 31276 25844 31332 25854
rect 30716 25788 31108 25844
rect 30716 25620 30772 25630
rect 30716 25526 30772 25564
rect 30604 25396 30660 25406
rect 30380 25394 30660 25396
rect 30380 25342 30606 25394
rect 30658 25342 30660 25394
rect 30380 25340 30660 25342
rect 30380 24834 30436 25340
rect 30604 25330 30660 25340
rect 30380 24782 30382 24834
rect 30434 24782 30436 24834
rect 30380 24770 30436 24782
rect 30268 24110 30270 24162
rect 30322 24110 30324 24162
rect 30268 24098 30324 24110
rect 30044 24052 30100 24062
rect 29820 24050 30100 24052
rect 29820 23998 30046 24050
rect 30098 23998 30100 24050
rect 29820 23996 30100 23998
rect 29708 23940 29764 23950
rect 29820 23940 29876 23996
rect 30044 23986 30100 23996
rect 29484 23938 29876 23940
rect 29484 23886 29710 23938
rect 29762 23886 29876 23938
rect 29484 23884 29876 23886
rect 29148 23716 29204 23726
rect 29148 23714 29316 23716
rect 29148 23662 29150 23714
rect 29202 23662 29316 23714
rect 29148 23660 29316 23662
rect 29148 23650 29204 23660
rect 28812 23314 28868 23324
rect 28588 23202 28644 23212
rect 28476 23090 28532 23100
rect 29148 23042 29204 23054
rect 29148 22990 29150 23042
rect 29202 22990 29204 23042
rect 28364 22932 28420 22942
rect 27804 22540 28308 22596
rect 28028 22372 28084 22382
rect 27356 22370 28084 22372
rect 27356 22318 28030 22370
rect 28082 22318 28084 22370
rect 27356 22316 28084 22318
rect 27356 22258 27412 22316
rect 28028 22306 28084 22316
rect 27356 22206 27358 22258
rect 27410 22206 27412 22258
rect 27356 22194 27412 22206
rect 27244 21812 27300 21822
rect 27244 20692 27300 21756
rect 27244 20598 27300 20636
rect 27356 20690 27412 20702
rect 27356 20638 27358 20690
rect 27410 20638 27412 20690
rect 27356 20356 27412 20638
rect 26908 20188 27188 20244
rect 27244 20300 27412 20356
rect 27804 20578 27860 20590
rect 27804 20526 27806 20578
rect 27858 20526 27860 20578
rect 26460 20018 26628 20020
rect 26460 19966 26462 20018
rect 26514 19966 26628 20018
rect 26460 19964 26628 19966
rect 26684 20018 26740 20030
rect 26684 19966 26686 20018
rect 26738 19966 26740 20018
rect 26348 19348 26404 19358
rect 26348 18450 26404 19292
rect 26348 18398 26350 18450
rect 26402 18398 26404 18450
rect 26348 18386 26404 18398
rect 26012 18162 26068 18172
rect 26460 17780 26516 19964
rect 26684 18564 26740 19966
rect 26796 20020 26852 20030
rect 26796 19926 26852 19964
rect 26740 18508 26852 18564
rect 26684 18498 26740 18508
rect 26684 17780 26740 17790
rect 26460 17778 26740 17780
rect 26460 17726 26686 17778
rect 26738 17726 26740 17778
rect 26460 17724 26740 17726
rect 26684 17714 26740 17724
rect 25452 17042 25508 17052
rect 26348 17108 26404 17118
rect 24780 16940 25284 16996
rect 24332 16884 24388 16894
rect 24332 16770 24388 16828
rect 24332 16718 24334 16770
rect 24386 16718 24388 16770
rect 24332 16706 24388 16718
rect 24668 16212 24724 16222
rect 24780 16212 24836 16940
rect 25452 16884 25508 16894
rect 25452 16790 25508 16828
rect 26124 16882 26180 16894
rect 26124 16830 26126 16882
rect 26178 16830 26180 16882
rect 24668 16210 24836 16212
rect 24668 16158 24670 16210
rect 24722 16158 24836 16210
rect 24668 16156 24836 16158
rect 26124 16212 26180 16830
rect 26348 16882 26404 17052
rect 26348 16830 26350 16882
rect 26402 16830 26404 16882
rect 26348 16818 26404 16830
rect 26796 16548 26852 18508
rect 26908 17108 26964 20188
rect 27020 20020 27076 20030
rect 27244 20020 27300 20300
rect 27804 20242 27860 20526
rect 27804 20190 27806 20242
rect 27858 20190 27860 20242
rect 27804 20178 27860 20190
rect 28140 20578 28196 20590
rect 28140 20526 28142 20578
rect 28194 20526 28196 20578
rect 28140 20244 28196 20526
rect 28252 20580 28308 22540
rect 28252 20514 28308 20524
rect 28252 20244 28308 20254
rect 28140 20188 28252 20244
rect 28252 20178 28308 20188
rect 27356 20132 27412 20142
rect 27356 20038 27412 20076
rect 27020 20018 27300 20020
rect 27020 19966 27022 20018
rect 27074 19966 27300 20018
rect 27020 19964 27300 19966
rect 27580 20020 27636 20030
rect 27020 19796 27076 19964
rect 27580 19926 27636 19964
rect 27692 19908 27748 19918
rect 27692 19814 27748 19852
rect 28252 19906 28308 19918
rect 28252 19854 28254 19906
rect 28306 19854 28308 19906
rect 27020 19730 27076 19740
rect 28252 18564 28308 19854
rect 28252 18498 28308 18508
rect 27132 18340 27188 18350
rect 27916 18340 27972 18350
rect 27132 18338 27860 18340
rect 27132 18286 27134 18338
rect 27186 18286 27860 18338
rect 27132 18284 27860 18286
rect 27132 18274 27188 18284
rect 27804 17890 27860 18284
rect 27804 17838 27806 17890
rect 27858 17838 27860 17890
rect 27804 17826 27860 17838
rect 27916 17778 27972 18284
rect 27916 17726 27918 17778
rect 27970 17726 27972 17778
rect 27916 17714 27972 17726
rect 26908 17042 26964 17052
rect 27692 17108 27748 17118
rect 27692 17014 27748 17052
rect 27132 16996 27188 17006
rect 27020 16994 27188 16996
rect 27020 16942 27134 16994
rect 27186 16942 27188 16994
rect 27020 16940 27188 16942
rect 26796 16492 26964 16548
rect 26796 16212 26852 16222
rect 24668 16146 24724 16156
rect 26124 16146 26180 16156
rect 26572 16156 26796 16212
rect 26460 15540 26516 15550
rect 25788 15538 26516 15540
rect 25788 15486 26462 15538
rect 26514 15486 26516 15538
rect 25788 15484 26516 15486
rect 25340 15316 25396 15326
rect 25228 15204 25284 15242
rect 24220 15092 24388 15148
rect 25228 15138 25284 15148
rect 23100 14478 23102 14530
rect 23154 14478 23156 14530
rect 23100 14466 23156 14478
rect 23548 13972 23604 13982
rect 23548 13858 23604 13916
rect 23884 13972 23940 15092
rect 24332 14308 24388 15092
rect 23884 13970 24276 13972
rect 23884 13918 23886 13970
rect 23938 13918 24276 13970
rect 23884 13916 24276 13918
rect 23884 13906 23940 13916
rect 23548 13806 23550 13858
rect 23602 13806 23604 13858
rect 22988 13748 23044 13758
rect 22988 13524 23044 13692
rect 23548 13636 23604 13806
rect 23660 13860 23716 13870
rect 23660 13766 23716 13804
rect 24220 13746 24276 13916
rect 24220 13694 24222 13746
rect 24274 13694 24276 13746
rect 24220 13682 24276 13694
rect 23548 13580 24052 13636
rect 22988 13468 23604 13524
rect 23548 13074 23604 13468
rect 23548 13022 23550 13074
rect 23602 13022 23604 13074
rect 22876 12292 22932 12302
rect 22876 12178 22932 12236
rect 22876 12126 22878 12178
rect 22930 12126 22932 12178
rect 22876 12114 22932 12126
rect 23212 11956 23268 11966
rect 22988 11954 23268 11956
rect 22988 11902 23214 11954
rect 23266 11902 23268 11954
rect 22988 11900 23268 11902
rect 22876 11844 22932 11854
rect 22652 10556 22820 10612
rect 22316 10500 22372 10510
rect 22316 10498 22708 10500
rect 22316 10446 22318 10498
rect 22370 10446 22708 10498
rect 22316 10444 22708 10446
rect 22316 10434 22372 10444
rect 22652 9714 22708 10444
rect 22652 9662 22654 9714
rect 22706 9662 22708 9714
rect 22652 9650 22708 9662
rect 22204 9550 22206 9602
rect 22258 9550 22260 9602
rect 22204 9380 22260 9550
rect 22764 9604 22820 10556
rect 22764 9538 22820 9548
rect 22204 9314 22260 9324
rect 22764 8930 22820 8942
rect 22764 8878 22766 8930
rect 22818 8878 22820 8930
rect 22316 8484 22372 8494
rect 22652 8484 22708 8494
rect 22316 8482 22708 8484
rect 22316 8430 22318 8482
rect 22370 8430 22654 8482
rect 22706 8430 22708 8482
rect 22316 8428 22708 8430
rect 22316 8418 22372 8428
rect 22652 8418 22708 8428
rect 21980 8372 22036 8382
rect 21980 8258 22036 8316
rect 21980 8206 21982 8258
rect 22034 8206 22036 8258
rect 21980 8194 22036 8206
rect 22428 8258 22484 8270
rect 22428 8206 22430 8258
rect 22482 8206 22484 8258
rect 21756 8148 21812 8158
rect 21756 8054 21812 8092
rect 22316 7924 22372 7934
rect 21532 7532 21700 7588
rect 22204 7588 22260 7598
rect 21532 7140 21588 7532
rect 22204 7494 22260 7532
rect 21868 7474 21924 7486
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 21644 7364 21700 7374
rect 21868 7364 21924 7422
rect 21700 7308 21924 7364
rect 22092 7362 22148 7374
rect 22092 7310 22094 7362
rect 22146 7310 22148 7362
rect 21644 7270 21700 7308
rect 21532 7084 21812 7140
rect 21420 7074 21476 7084
rect 20972 6804 21028 6814
rect 20524 6066 20580 6076
rect 20748 6468 20804 6478
rect 20748 5684 20804 6412
rect 20748 5618 20804 5628
rect 20636 5572 20692 5582
rect 20636 5122 20692 5516
rect 20636 5070 20638 5122
rect 20690 5070 20692 5122
rect 20636 5058 20692 5070
rect 20860 5348 20916 5358
rect 20412 4958 20414 5010
rect 20466 4958 20468 5010
rect 20412 4946 20468 4958
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18732 4386 18788 4396
rect 18060 4286 18062 4338
rect 18114 4286 18116 4338
rect 18060 4274 18116 4286
rect 18732 4228 18788 4238
rect 18732 4134 18788 4172
rect 20860 4226 20916 5292
rect 20860 4174 20862 4226
rect 20914 4174 20916 4226
rect 20860 4162 20916 4174
rect 18620 3666 18676 3678
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17276 3490 17332 3502
rect 17612 3556 17668 3566
rect 17612 3462 17668 3500
rect 18620 3388 18676 3614
rect 16828 924 17220 980
rect 18396 3332 18676 3388
rect 20076 3668 20132 3678
rect 20076 3332 20132 3612
rect 20972 3554 21028 6748
rect 21644 6692 21700 6702
rect 21756 6692 21812 7084
rect 21868 6916 21924 6926
rect 21868 6914 22036 6916
rect 21868 6862 21870 6914
rect 21922 6862 22036 6914
rect 21868 6860 22036 6862
rect 21868 6850 21924 6860
rect 21868 6692 21924 6702
rect 21756 6690 21924 6692
rect 21756 6638 21870 6690
rect 21922 6638 21924 6690
rect 21756 6636 21924 6638
rect 21308 6578 21364 6590
rect 21308 6526 21310 6578
rect 21362 6526 21364 6578
rect 21308 6132 21364 6526
rect 21532 6580 21588 6590
rect 21532 6486 21588 6524
rect 21308 6066 21364 6076
rect 21644 6020 21700 6636
rect 21420 6018 21700 6020
rect 21420 5966 21646 6018
rect 21698 5966 21700 6018
rect 21420 5964 21700 5966
rect 21308 5124 21364 5134
rect 21420 5124 21476 5964
rect 21644 5954 21700 5964
rect 21756 6466 21812 6478
rect 21756 6414 21758 6466
rect 21810 6414 21812 6466
rect 21364 5122 21476 5124
rect 21364 5070 21422 5122
rect 21474 5070 21476 5122
rect 21364 5068 21476 5070
rect 21308 4338 21364 5068
rect 21420 5058 21476 5068
rect 21308 4286 21310 4338
rect 21362 4286 21364 4338
rect 21308 4274 21364 4286
rect 21532 4452 21588 4462
rect 21756 4452 21812 6414
rect 21868 6468 21924 6636
rect 21868 6402 21924 6412
rect 21980 5124 22036 6860
rect 22092 5234 22148 7310
rect 22316 7028 22372 7868
rect 22428 7476 22484 8206
rect 22540 8036 22596 8046
rect 22764 8036 22820 8878
rect 22540 8034 22820 8036
rect 22540 7982 22542 8034
rect 22594 7982 22820 8034
rect 22540 7980 22820 7982
rect 22876 8148 22932 11788
rect 22988 9826 23044 11900
rect 23212 11890 23268 11900
rect 23548 11396 23604 13022
rect 23996 12292 24052 13580
rect 23996 12198 24052 12236
rect 24108 12404 24164 12414
rect 23660 12178 23716 12190
rect 23660 12126 23662 12178
rect 23714 12126 23716 12178
rect 23660 12068 23716 12126
rect 23884 12180 23940 12190
rect 23884 12086 23940 12124
rect 24108 12178 24164 12348
rect 24108 12126 24110 12178
rect 24162 12126 24164 12178
rect 24108 12114 24164 12126
rect 23660 12002 23716 12012
rect 23772 11396 23828 11406
rect 23604 11394 23828 11396
rect 23604 11342 23774 11394
rect 23826 11342 23828 11394
rect 23604 11340 23828 11342
rect 23548 11302 23604 11340
rect 23772 11330 23828 11340
rect 24332 10276 24388 14252
rect 24556 13972 24612 13982
rect 24556 13970 24724 13972
rect 24556 13918 24558 13970
rect 24610 13918 24724 13970
rect 24556 13916 24724 13918
rect 24556 13906 24612 13916
rect 24556 13748 24612 13758
rect 24556 13654 24612 13692
rect 24444 13524 24500 13534
rect 24444 13430 24500 13468
rect 24444 11956 24500 11966
rect 24444 10498 24500 11900
rect 24556 11508 24612 11518
rect 24668 11508 24724 13916
rect 25228 13524 25284 13534
rect 25228 13430 25284 13468
rect 25340 12178 25396 15260
rect 25788 15314 25844 15484
rect 26460 15474 26516 15484
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15250 25844 15262
rect 26236 15314 26292 15326
rect 26236 15262 26238 15314
rect 26290 15262 26292 15314
rect 25564 15204 25620 15242
rect 26236 15148 26292 15262
rect 26460 15316 26516 15326
rect 26572 15316 26628 16156
rect 26796 16118 26852 16156
rect 26908 15988 26964 16492
rect 26460 15314 26628 15316
rect 26460 15262 26462 15314
rect 26514 15262 26628 15314
rect 26460 15260 26628 15262
rect 26684 15932 26964 15988
rect 26684 15316 26740 15932
rect 26460 15250 26516 15260
rect 26684 15222 26740 15260
rect 26796 15204 26852 15214
rect 26908 15204 26964 15214
rect 26852 15202 26964 15204
rect 26852 15150 26910 15202
rect 26962 15150 26964 15202
rect 26852 15148 26964 15150
rect 25564 13746 25620 15148
rect 25900 15092 26292 15148
rect 25900 14642 25956 15092
rect 26236 15026 26292 15036
rect 26572 15092 26852 15148
rect 26908 15138 26964 15148
rect 26572 14754 26628 15092
rect 26572 14702 26574 14754
rect 26626 14702 26628 14754
rect 26572 14690 26628 14702
rect 26908 14756 26964 14766
rect 27020 14756 27076 16940
rect 27132 16930 27188 16940
rect 27580 16996 27636 17006
rect 27244 16884 27300 16894
rect 27244 16882 27524 16884
rect 27244 16830 27246 16882
rect 27298 16830 27524 16882
rect 27244 16828 27524 16830
rect 27244 16818 27300 16828
rect 27132 16660 27188 16670
rect 27132 16658 27300 16660
rect 27132 16606 27134 16658
rect 27186 16606 27300 16658
rect 27132 16604 27300 16606
rect 27132 16594 27188 16604
rect 27132 15874 27188 15886
rect 27132 15822 27134 15874
rect 27186 15822 27188 15874
rect 27132 15202 27188 15822
rect 27132 15150 27134 15202
rect 27186 15150 27188 15202
rect 27132 15138 27188 15150
rect 27132 14756 27188 14766
rect 27020 14754 27188 14756
rect 27020 14702 27134 14754
rect 27186 14702 27188 14754
rect 27020 14700 27188 14702
rect 25900 14590 25902 14642
rect 25954 14590 25956 14642
rect 25900 14578 25956 14590
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 14084 26404 14254
rect 26348 14018 26404 14028
rect 26460 14306 26516 14318
rect 26460 14254 26462 14306
rect 26514 14254 26516 14306
rect 25564 13694 25566 13746
rect 25618 13694 25620 13746
rect 25564 13682 25620 13694
rect 26460 13748 26516 14254
rect 26460 13682 26516 13692
rect 26572 14084 26628 14094
rect 26572 13746 26628 14028
rect 26796 13860 26852 13870
rect 26796 13766 26852 13804
rect 26908 13858 26964 14700
rect 27132 14690 27188 14700
rect 27244 14756 27300 16604
rect 27244 14690 27300 14700
rect 27356 15988 27412 15998
rect 27356 15314 27412 15932
rect 27468 15540 27524 16828
rect 27580 16098 27636 16940
rect 28140 16996 28196 17006
rect 28140 16902 28196 16940
rect 28364 16548 28420 22876
rect 29148 22258 29204 22990
rect 29148 22206 29150 22258
rect 29202 22206 29204 22258
rect 28588 22146 28644 22158
rect 29036 22148 29092 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 21476 28644 22094
rect 28700 22146 29092 22148
rect 28700 22094 29038 22146
rect 29090 22094 29092 22146
rect 28700 22092 29092 22094
rect 28700 21698 28756 22092
rect 29036 22082 29092 22092
rect 28700 21646 28702 21698
rect 28754 21646 28756 21698
rect 28700 21634 28756 21646
rect 28476 20580 28532 20590
rect 28476 20486 28532 20524
rect 28588 20244 28644 21420
rect 29036 21364 29092 21374
rect 29036 20802 29092 21308
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20738 29092 20750
rect 28588 20178 28644 20188
rect 29148 20132 29204 22206
rect 29148 20066 29204 20076
rect 28700 19908 28756 19918
rect 29148 19908 29204 19918
rect 28700 19906 29204 19908
rect 28700 19854 28702 19906
rect 28754 19854 29150 19906
rect 29202 19854 29204 19906
rect 28700 19852 29204 19854
rect 28700 19796 28756 19852
rect 29148 19842 29204 19852
rect 28588 17556 28644 17566
rect 28588 17462 28644 17500
rect 28364 16482 28420 16492
rect 28476 16770 28532 16782
rect 28476 16718 28478 16770
rect 28530 16718 28532 16770
rect 27580 16046 27582 16098
rect 27634 16046 27636 16098
rect 27580 16034 27636 16046
rect 27692 16212 27748 16222
rect 28476 16212 28532 16718
rect 28588 16212 28644 16222
rect 28476 16156 28588 16212
rect 27692 16098 27748 16156
rect 28588 16118 28644 16156
rect 27692 16046 27694 16098
rect 27746 16046 27748 16098
rect 27468 15474 27524 15484
rect 27580 15652 27636 15662
rect 27580 15316 27636 15596
rect 27692 15540 27748 16046
rect 27804 15988 27860 15998
rect 27804 15894 27860 15932
rect 28476 15876 28532 15886
rect 28364 15874 28532 15876
rect 28364 15822 28478 15874
rect 28530 15822 28532 15874
rect 28364 15820 28532 15822
rect 27804 15540 27860 15550
rect 27692 15538 27860 15540
rect 27692 15486 27806 15538
rect 27858 15486 27860 15538
rect 27692 15484 27860 15486
rect 27804 15474 27860 15484
rect 27916 15428 27972 15438
rect 27916 15334 27972 15372
rect 27356 15262 27358 15314
rect 27410 15262 27412 15314
rect 27356 15092 27412 15262
rect 27356 14644 27412 15036
rect 27356 14578 27412 14588
rect 27468 15314 27636 15316
rect 27468 15262 27582 15314
rect 27634 15262 27636 15314
rect 27468 15260 27636 15262
rect 27132 14532 27188 14542
rect 27132 14418 27188 14476
rect 27132 14366 27134 14418
rect 27186 14366 27188 14418
rect 27132 14354 27188 14366
rect 27244 14420 27300 14430
rect 27468 14420 27524 15260
rect 27580 15250 27636 15260
rect 28028 15316 28084 15326
rect 28028 15222 28084 15260
rect 28364 15316 28420 15820
rect 28476 15810 28532 15820
rect 28476 15652 28532 15662
rect 28476 15538 28532 15596
rect 28476 15486 28478 15538
rect 28530 15486 28532 15538
rect 28476 15474 28532 15486
rect 28364 15250 28420 15260
rect 28588 15314 28644 15326
rect 28588 15262 28590 15314
rect 28642 15262 28644 15314
rect 27244 14418 27524 14420
rect 27244 14366 27246 14418
rect 27298 14366 27524 14418
rect 27244 14364 27524 14366
rect 27692 15092 27748 15102
rect 27692 14420 27748 15036
rect 28364 15092 28420 15102
rect 27244 14354 27300 14364
rect 27692 14326 27748 14364
rect 28028 14530 28084 14542
rect 28028 14478 28030 14530
rect 28082 14478 28084 14530
rect 28028 14084 28084 14478
rect 28028 14018 28084 14028
rect 26908 13806 26910 13858
rect 26962 13806 26964 13858
rect 26908 13794 26964 13806
rect 27692 13860 27748 13870
rect 28028 13860 28084 13870
rect 27692 13858 27860 13860
rect 27692 13806 27694 13858
rect 27746 13806 27860 13858
rect 27692 13804 27860 13806
rect 27692 13794 27748 13804
rect 26572 13694 26574 13746
rect 26626 13694 26628 13746
rect 25788 13636 25844 13646
rect 25788 13542 25844 13580
rect 26572 13636 26628 13694
rect 26460 13524 26516 13534
rect 25340 12126 25342 12178
rect 25394 12126 25396 12178
rect 25340 12114 25396 12126
rect 25564 12404 25620 12414
rect 25564 12178 25620 12348
rect 26460 12292 26516 13468
rect 25564 12126 25566 12178
rect 25618 12126 25620 12178
rect 25564 12114 25620 12126
rect 25788 12180 25844 12190
rect 25788 12086 25844 12124
rect 26460 12178 26516 12236
rect 26460 12126 26462 12178
rect 26514 12126 26516 12178
rect 26460 12114 26516 12126
rect 24556 11506 24724 11508
rect 24556 11454 24558 11506
rect 24610 11454 24724 11506
rect 24556 11452 24724 11454
rect 25676 12066 25732 12078
rect 25676 12014 25678 12066
rect 25730 12014 25732 12066
rect 24556 11442 24612 11452
rect 25676 10724 25732 12014
rect 26124 12068 26180 12078
rect 26124 11974 26180 12012
rect 26572 11508 26628 13580
rect 27468 13746 27524 13758
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13300 27524 13694
rect 27804 13524 27860 13804
rect 28028 13766 28084 13804
rect 27804 13468 28084 13524
rect 27916 13300 27972 13310
rect 27020 13244 27860 13300
rect 27020 13186 27076 13244
rect 27020 13134 27022 13186
rect 27074 13134 27076 13186
rect 27020 13122 27076 13134
rect 27692 13076 27748 13086
rect 27356 12964 27412 12974
rect 27356 12962 27636 12964
rect 27356 12910 27358 12962
rect 27410 12910 27636 12962
rect 27356 12908 27636 12910
rect 27356 12898 27412 12908
rect 26908 12852 26964 12862
rect 26908 12850 27076 12852
rect 26908 12798 26910 12850
rect 26962 12798 27076 12850
rect 26908 12796 27076 12798
rect 26908 12786 26964 12796
rect 27020 12292 27076 12796
rect 27468 12740 27524 12750
rect 27132 12292 27188 12302
rect 27020 12290 27188 12292
rect 27020 12238 27134 12290
rect 27186 12238 27188 12290
rect 27020 12236 27188 12238
rect 26908 12180 26964 12190
rect 26908 12086 26964 12124
rect 26684 12066 26740 12078
rect 26684 12014 26686 12066
rect 26738 12014 26740 12066
rect 26684 11956 26740 12014
rect 26684 11890 26740 11900
rect 27132 11956 27188 12236
rect 27244 12292 27300 12302
rect 27244 12198 27300 12236
rect 27132 11890 27188 11900
rect 26684 11508 26740 11518
rect 26572 11506 26740 11508
rect 26572 11454 26686 11506
rect 26738 11454 26740 11506
rect 26572 11452 26740 11454
rect 26684 11442 26740 11452
rect 27244 11172 27300 11182
rect 27244 11078 27300 11116
rect 27244 10948 27300 10958
rect 26012 10724 26068 10734
rect 25676 10722 26068 10724
rect 25676 10670 26014 10722
rect 26066 10670 26068 10722
rect 25676 10668 26068 10670
rect 26012 10658 26068 10668
rect 24444 10446 24446 10498
rect 24498 10446 24500 10498
rect 24444 10434 24500 10446
rect 25340 10610 25396 10622
rect 25340 10558 25342 10610
rect 25394 10558 25396 10610
rect 24332 10220 24500 10276
rect 22988 9774 22990 9826
rect 23042 9774 23044 9826
rect 22988 9762 23044 9774
rect 23324 9938 23380 9950
rect 23324 9886 23326 9938
rect 23378 9886 23380 9938
rect 23324 8482 23380 9886
rect 24220 9940 24276 9950
rect 24220 9846 24276 9884
rect 23660 9716 23716 9726
rect 23660 9714 24388 9716
rect 23660 9662 23662 9714
rect 23714 9662 24388 9714
rect 23660 9660 24388 9662
rect 23660 9650 23716 9660
rect 23436 9604 23492 9614
rect 23436 9492 23492 9548
rect 23436 9436 23716 9492
rect 23324 8430 23326 8482
rect 23378 8430 23380 8482
rect 23324 8418 23380 8430
rect 23548 9042 23604 9054
rect 23548 8990 23550 9042
rect 23602 8990 23604 9042
rect 22540 7970 22596 7980
rect 22876 7812 22932 8092
rect 23212 8036 23268 8046
rect 23212 7942 23268 7980
rect 22876 7756 23044 7812
rect 22988 7698 23044 7756
rect 22988 7646 22990 7698
rect 23042 7646 23044 7698
rect 22988 7634 23044 7646
rect 22876 7588 22932 7598
rect 22876 7494 22932 7532
rect 22428 7410 22484 7420
rect 22652 7474 22708 7486
rect 22652 7422 22654 7474
rect 22706 7422 22708 7474
rect 22652 7364 22708 7422
rect 22652 7298 22708 7308
rect 22764 7474 22820 7486
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22316 6972 22708 7028
rect 22652 6914 22708 6972
rect 22652 6862 22654 6914
rect 22706 6862 22708 6914
rect 22652 6850 22708 6862
rect 22764 5572 22820 7422
rect 23212 7476 23268 7486
rect 23212 7474 23492 7476
rect 23212 7422 23214 7474
rect 23266 7422 23492 7474
rect 23212 7420 23492 7422
rect 23212 7410 23268 7420
rect 23100 7252 23156 7262
rect 22764 5506 22820 5516
rect 22876 6580 22932 6590
rect 23100 6580 23156 7196
rect 23324 7252 23380 7262
rect 22876 6578 23156 6580
rect 22876 6526 22878 6578
rect 22930 6526 23156 6578
rect 22876 6524 23156 6526
rect 23212 6802 23268 6814
rect 23212 6750 23214 6802
rect 23266 6750 23268 6802
rect 22092 5182 22094 5234
rect 22146 5182 22148 5234
rect 22092 5170 22148 5182
rect 22876 5236 22932 6524
rect 23212 5908 23268 6750
rect 23324 6468 23380 7196
rect 23436 6914 23492 7420
rect 23436 6862 23438 6914
rect 23490 6862 23492 6914
rect 23436 6804 23492 6862
rect 23436 6738 23492 6748
rect 23548 6692 23604 8990
rect 23660 8932 23716 9436
rect 24332 9044 24388 9660
rect 23996 8932 24052 8942
rect 23660 8930 24052 8932
rect 23660 8878 23998 8930
rect 24050 8878 24052 8930
rect 23660 8876 24052 8878
rect 23660 8372 23716 8382
rect 23660 8278 23716 8316
rect 23660 8148 23716 8158
rect 23660 7698 23716 8092
rect 23996 8036 24052 8876
rect 24108 8260 24164 8270
rect 24108 8166 24164 8204
rect 24332 8258 24388 8988
rect 24444 8820 24500 10220
rect 25340 10052 25396 10558
rect 25340 9986 25396 9996
rect 27132 10052 27188 10062
rect 25004 9940 25060 9950
rect 24780 9268 24836 9278
rect 24780 9174 24836 9212
rect 24444 8754 24500 8764
rect 25004 9156 25060 9884
rect 26572 9940 26628 9950
rect 25228 9716 25284 9726
rect 24332 8206 24334 8258
rect 24386 8206 24388 8258
rect 24332 8194 24388 8206
rect 25004 8258 25060 9100
rect 25116 9660 25228 9716
rect 25116 8370 25172 9660
rect 25228 9650 25284 9660
rect 26348 9716 26404 9726
rect 26348 9622 26404 9660
rect 25228 9268 25284 9278
rect 25228 9042 25284 9212
rect 26572 9266 26628 9884
rect 27132 9826 27188 9996
rect 27132 9774 27134 9826
rect 27186 9774 27188 9826
rect 27132 9762 27188 9774
rect 26572 9214 26574 9266
rect 26626 9214 26628 9266
rect 26572 9202 26628 9214
rect 27132 9268 27188 9278
rect 27244 9268 27300 10892
rect 27132 9266 27300 9268
rect 27132 9214 27134 9266
rect 27186 9214 27300 9266
rect 27132 9212 27300 9214
rect 27356 9268 27412 9278
rect 27132 9202 27188 9212
rect 25788 9154 25844 9166
rect 26012 9156 26068 9166
rect 25788 9102 25790 9154
rect 25842 9102 25844 9154
rect 25228 8990 25230 9042
rect 25282 8990 25284 9042
rect 25228 8978 25284 8990
rect 25564 9044 25620 9054
rect 25564 8950 25620 8988
rect 25116 8318 25118 8370
rect 25170 8318 25172 8370
rect 25116 8306 25172 8318
rect 25676 8930 25732 8942
rect 25676 8878 25678 8930
rect 25730 8878 25732 8930
rect 25004 8206 25006 8258
rect 25058 8206 25060 8258
rect 25004 8194 25060 8206
rect 25564 8260 25620 8270
rect 25676 8260 25732 8878
rect 25564 8258 25732 8260
rect 25564 8206 25566 8258
rect 25618 8206 25732 8258
rect 25564 8204 25732 8206
rect 25564 8194 25620 8204
rect 25340 8148 25396 8158
rect 23996 7980 24164 8036
rect 23660 7646 23662 7698
rect 23714 7646 23716 7698
rect 23660 7634 23716 7646
rect 23548 6626 23604 6636
rect 23660 7140 23716 7150
rect 23548 6468 23604 6478
rect 23324 6466 23604 6468
rect 23324 6414 23550 6466
rect 23602 6414 23604 6466
rect 23324 6412 23604 6414
rect 23548 6402 23604 6412
rect 23212 5842 23268 5852
rect 23660 5906 23716 7084
rect 23660 5854 23662 5906
rect 23714 5854 23716 5906
rect 23660 5842 23716 5854
rect 23996 6690 24052 6702
rect 23996 6638 23998 6690
rect 24050 6638 24052 6690
rect 22876 5170 22932 5180
rect 23660 5460 23716 5470
rect 21980 5058 22036 5068
rect 21980 4452 22036 4462
rect 21756 4450 22036 4452
rect 21756 4398 21982 4450
rect 22034 4398 22036 4450
rect 21756 4396 22036 4398
rect 20972 3502 20974 3554
rect 21026 3502 21028 3554
rect 20972 3490 21028 3502
rect 16828 800 16884 924
rect 18396 800 18452 3332
rect 20076 3276 20244 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 2996 20244 3276
rect 19964 2940 20244 2996
rect 19964 800 20020 2940
rect 21532 800 21588 4396
rect 21980 4386 22036 4396
rect 23660 3778 23716 5404
rect 23660 3726 23662 3778
rect 23714 3726 23716 3778
rect 23660 3714 23716 3726
rect 23772 5124 23828 5134
rect 21868 3668 21924 3678
rect 21868 3574 21924 3612
rect 23772 3666 23828 5068
rect 23996 4676 24052 6638
rect 24108 5684 24164 7980
rect 24444 8034 24500 8046
rect 24444 7982 24446 8034
rect 24498 7982 24500 8034
rect 24444 7924 24500 7982
rect 24444 7858 24500 7868
rect 24668 8034 24724 8046
rect 24668 7982 24670 8034
rect 24722 7982 24724 8034
rect 24668 7588 24724 7982
rect 25228 7588 25284 7598
rect 24668 7586 25284 7588
rect 24668 7534 25230 7586
rect 25282 7534 25284 7586
rect 24668 7532 25284 7534
rect 24332 7476 24388 7486
rect 24332 7382 24388 7420
rect 24556 7476 24612 7486
rect 24668 7476 24724 7532
rect 25228 7522 25284 7532
rect 24556 7474 24724 7476
rect 24556 7422 24558 7474
rect 24610 7422 24724 7474
rect 24556 7420 24724 7422
rect 24556 7410 24612 7420
rect 24220 7364 24276 7374
rect 24220 7270 24276 7308
rect 24668 7250 24724 7262
rect 24668 7198 24670 7250
rect 24722 7198 24724 7250
rect 24668 6802 24724 7198
rect 24668 6750 24670 6802
rect 24722 6750 24724 6802
rect 24668 6738 24724 6750
rect 24780 6692 24836 6702
rect 24780 6132 24836 6636
rect 24220 5684 24276 5694
rect 24108 5628 24220 5684
rect 24220 5618 24276 5628
rect 24556 5460 24612 5470
rect 24220 5236 24276 5246
rect 24220 5142 24276 5180
rect 24556 5234 24612 5404
rect 24556 5182 24558 5234
rect 24610 5182 24612 5234
rect 24556 5170 24612 5182
rect 24780 5234 24836 6076
rect 25340 6020 25396 8092
rect 25788 8148 25844 9102
rect 25788 8082 25844 8092
rect 25900 9100 26012 9156
rect 25900 8484 25956 9100
rect 26012 9062 26068 9100
rect 25900 8428 26292 8484
rect 25900 8146 25956 8428
rect 25900 8094 25902 8146
rect 25954 8094 25956 8146
rect 25900 8082 25956 8094
rect 26124 8258 26180 8270
rect 26124 8206 26126 8258
rect 26178 8206 26180 8258
rect 26124 8148 26180 8206
rect 26124 8082 26180 8092
rect 26012 8034 26068 8046
rect 26012 7982 26014 8034
rect 26066 7982 26068 8034
rect 25564 7586 25620 7598
rect 25564 7534 25566 7586
rect 25618 7534 25620 7586
rect 25564 6804 25620 7534
rect 26012 7476 26068 7982
rect 26236 7586 26292 8428
rect 27356 8370 27412 9212
rect 27468 9266 27524 12684
rect 27580 12404 27636 12908
rect 27580 11620 27636 12348
rect 27692 12962 27748 13020
rect 27692 12910 27694 12962
rect 27746 12910 27748 12962
rect 27692 12290 27748 12910
rect 27804 12962 27860 13244
rect 27916 13074 27972 13244
rect 27916 13022 27918 13074
rect 27970 13022 27972 13074
rect 27916 13010 27972 13022
rect 27804 12910 27806 12962
rect 27858 12910 27860 12962
rect 27804 12898 27860 12910
rect 28028 12964 28084 13468
rect 28028 12404 28084 12908
rect 28028 12348 28308 12404
rect 27692 12238 27694 12290
rect 27746 12238 27748 12290
rect 27692 12226 27748 12238
rect 27804 12290 27860 12302
rect 27804 12238 27806 12290
rect 27858 12238 27860 12290
rect 27804 11620 27860 12238
rect 28028 12180 28084 12190
rect 28028 12086 28084 12124
rect 27580 11618 27860 11620
rect 27580 11566 27582 11618
rect 27634 11566 27860 11618
rect 27580 11564 27860 11566
rect 27580 11554 27636 11564
rect 27692 11284 27748 11294
rect 27692 11282 27972 11284
rect 27692 11230 27694 11282
rect 27746 11230 27972 11282
rect 27692 11228 27972 11230
rect 27692 11218 27748 11228
rect 27468 9214 27470 9266
rect 27522 9214 27524 9266
rect 27468 8484 27524 9214
rect 27692 10724 27748 10734
rect 27692 10276 27748 10668
rect 27916 10500 27972 11228
rect 28028 11170 28084 11182
rect 28028 11118 28030 11170
rect 28082 11118 28084 11170
rect 28028 10724 28084 11118
rect 28028 10658 28084 10668
rect 28140 10500 28196 10510
rect 27916 10498 28196 10500
rect 27916 10446 28142 10498
rect 28194 10446 28196 10498
rect 27916 10444 28196 10446
rect 28252 10500 28308 12348
rect 28364 11394 28420 15036
rect 28588 14980 28644 15262
rect 28700 15316 28756 19740
rect 29036 19348 29092 19358
rect 28700 15250 28756 15260
rect 28812 19346 29092 19348
rect 28812 19294 29038 19346
rect 29090 19294 29092 19346
rect 28812 19292 29092 19294
rect 28812 15148 28868 19292
rect 29036 19282 29092 19292
rect 29260 19236 29316 23660
rect 29484 23154 29540 23884
rect 29708 23874 29764 23884
rect 30604 23716 30660 23726
rect 30604 23714 30996 23716
rect 30604 23662 30606 23714
rect 30658 23662 30996 23714
rect 30604 23660 30996 23662
rect 30604 23650 30660 23660
rect 29484 23102 29486 23154
rect 29538 23102 29540 23154
rect 29484 23090 29540 23102
rect 29708 23156 29764 23166
rect 29708 23062 29764 23100
rect 30492 23154 30548 23166
rect 30492 23102 30494 23154
rect 30546 23102 30548 23154
rect 30044 22932 30100 22942
rect 30044 22838 30100 22876
rect 30380 22484 30436 22494
rect 29372 22428 29764 22484
rect 29372 22370 29428 22428
rect 29372 22318 29374 22370
rect 29426 22318 29428 22370
rect 29372 22306 29428 22318
rect 29596 22258 29652 22270
rect 29596 22206 29598 22258
rect 29650 22206 29652 22258
rect 29484 21588 29540 21598
rect 29484 21494 29540 21532
rect 29596 20914 29652 22206
rect 29708 21810 29764 22428
rect 30268 22428 30380 22484
rect 30044 22372 30100 22382
rect 30044 22278 30100 22316
rect 29708 21758 29710 21810
rect 29762 21758 29764 21810
rect 29708 21746 29764 21758
rect 30044 21588 30100 21598
rect 29596 20862 29598 20914
rect 29650 20862 29652 20914
rect 29596 20850 29652 20862
rect 29932 21532 30044 21588
rect 29708 20804 29764 20814
rect 29708 20710 29764 20748
rect 29596 20692 29652 20702
rect 29484 20578 29540 20590
rect 29484 20526 29486 20578
rect 29538 20526 29540 20578
rect 29484 20468 29540 20526
rect 29484 20402 29540 20412
rect 29148 19180 29316 19236
rect 29372 20244 29428 20254
rect 29036 18900 29092 18910
rect 29036 15148 29092 18844
rect 29148 18452 29204 19180
rect 29260 19012 29316 19022
rect 29372 19012 29428 20188
rect 29596 19906 29652 20636
rect 29596 19854 29598 19906
rect 29650 19854 29652 19906
rect 29596 19458 29652 19854
rect 29596 19406 29598 19458
rect 29650 19406 29652 19458
rect 29596 19394 29652 19406
rect 29932 19234 29988 21532
rect 30044 21522 30100 21532
rect 30156 21588 30212 21598
rect 30268 21588 30324 22428
rect 30380 22418 30436 22428
rect 30492 22372 30548 23102
rect 30828 23044 30884 23054
rect 30828 22950 30884 22988
rect 30548 22316 30772 22372
rect 30492 22306 30548 22316
rect 30156 21586 30324 21588
rect 30156 21534 30158 21586
rect 30210 21534 30324 21586
rect 30156 21532 30324 21534
rect 30380 21812 30436 21822
rect 30156 20804 30212 21532
rect 30380 21364 30436 21756
rect 30716 21700 30772 22316
rect 30940 22036 30996 23660
rect 31052 23156 31108 25788
rect 31164 25620 31220 25658
rect 31164 25554 31220 25564
rect 31276 25506 31332 25788
rect 31276 25454 31278 25506
rect 31330 25454 31332 25506
rect 31276 25442 31332 25454
rect 31164 25396 31220 25406
rect 31164 25302 31220 25340
rect 31164 24164 31220 24174
rect 31164 23940 31220 24108
rect 31164 23938 31332 23940
rect 31164 23886 31166 23938
rect 31218 23886 31332 23938
rect 31164 23884 31332 23886
rect 31164 23874 31220 23884
rect 31164 23156 31220 23166
rect 31052 23100 31164 23156
rect 31164 23062 31220 23100
rect 31276 22260 31332 23884
rect 31388 23380 31444 27244
rect 31500 27188 31556 29484
rect 31612 29474 31668 29484
rect 31612 28980 31668 28990
rect 31612 28196 31668 28924
rect 31612 28082 31668 28140
rect 31612 28030 31614 28082
rect 31666 28030 31668 28082
rect 31612 28018 31668 28030
rect 31612 27188 31668 27198
rect 31500 27186 31668 27188
rect 31500 27134 31614 27186
rect 31666 27134 31668 27186
rect 31500 27132 31668 27134
rect 31612 27122 31668 27132
rect 31724 26964 31780 29708
rect 31612 26908 31780 26964
rect 31836 29314 31892 29326
rect 31836 29262 31838 29314
rect 31890 29262 31892 29314
rect 31500 25508 31556 25518
rect 31500 25414 31556 25452
rect 31612 23548 31668 26908
rect 31836 25844 31892 29262
rect 32060 28756 32116 30718
rect 32172 29876 32228 30830
rect 32508 30884 32564 30940
rect 32172 29810 32228 29820
rect 32396 30210 32452 30222
rect 32396 30158 32398 30210
rect 32450 30158 32452 30210
rect 32284 29652 32340 29662
rect 32060 28662 32116 28700
rect 32172 29596 32284 29652
rect 32172 28532 32228 29596
rect 32284 29586 32340 29596
rect 32284 29428 32340 29438
rect 32284 29334 32340 29372
rect 32396 28756 32452 30158
rect 31836 25778 31892 25788
rect 31948 28476 32228 28532
rect 32284 28700 32452 28756
rect 31948 28082 32004 28476
rect 32284 28308 32340 28700
rect 32508 28644 32564 30828
rect 32956 29986 33012 29998
rect 32956 29934 32958 29986
rect 33010 29934 33012 29986
rect 32956 29876 33012 29934
rect 32620 29428 32676 29438
rect 32676 29372 32900 29428
rect 32620 29362 32676 29372
rect 32732 28644 32788 28654
rect 32508 28642 32788 28644
rect 32508 28590 32734 28642
rect 32786 28590 32788 28642
rect 32508 28588 32788 28590
rect 32732 28578 32788 28588
rect 32396 28532 32452 28542
rect 32396 28438 32452 28476
rect 32508 28420 32564 28430
rect 32508 28326 32564 28364
rect 32284 28252 32452 28308
rect 31948 28030 31950 28082
rect 32002 28030 32004 28082
rect 31948 25508 32004 28030
rect 32060 28196 32116 28206
rect 32060 28082 32116 28140
rect 32060 28030 32062 28082
rect 32114 28030 32116 28082
rect 32060 28018 32116 28030
rect 32284 28084 32340 28094
rect 32284 27990 32340 28028
rect 32172 27748 32228 27786
rect 32172 27682 32228 27692
rect 32396 26404 32452 28252
rect 32508 27860 32564 27870
rect 32508 27766 32564 27804
rect 32844 27636 32900 29372
rect 32508 27580 32900 27636
rect 32508 27188 32564 27580
rect 32956 27524 33012 29820
rect 33180 29652 33236 29662
rect 33292 29652 33348 31054
rect 33404 30996 33460 31276
rect 33516 30996 33572 31006
rect 33404 30994 33572 30996
rect 33404 30942 33518 30994
rect 33570 30942 33572 30994
rect 33404 30940 33572 30942
rect 33404 30212 33460 30940
rect 33516 30930 33572 30940
rect 33628 30324 33684 32620
rect 33740 32610 33796 32620
rect 34076 32562 34132 32574
rect 34076 32510 34078 32562
rect 34130 32510 34132 32562
rect 34076 32004 34132 32510
rect 34076 31938 34132 31948
rect 33964 31778 34020 31790
rect 33964 31726 33966 31778
rect 34018 31726 34020 31778
rect 33404 30146 33460 30156
rect 33516 30268 33684 30324
rect 33852 31332 33908 31342
rect 33404 29988 33460 29998
rect 33404 29894 33460 29932
rect 33236 29596 33348 29652
rect 33404 29652 33460 29662
rect 33180 29558 33236 29596
rect 33404 29558 33460 29596
rect 33516 29650 33572 30268
rect 33740 30212 33796 30222
rect 33516 29598 33518 29650
rect 33570 29598 33572 29650
rect 33292 29428 33348 29438
rect 33180 28756 33236 28766
rect 33180 28662 33236 28700
rect 33292 28308 33348 29372
rect 33292 28242 33348 28252
rect 33404 28644 33460 28654
rect 33180 27860 33236 27870
rect 33404 27860 33460 28588
rect 33516 28084 33572 29598
rect 33628 30210 33796 30212
rect 33628 30158 33742 30210
rect 33794 30158 33796 30210
rect 33628 30156 33796 30158
rect 33628 29428 33684 30156
rect 33740 30146 33796 30156
rect 33628 29362 33684 29372
rect 33740 29426 33796 29438
rect 33740 29374 33742 29426
rect 33794 29374 33796 29426
rect 33740 28756 33796 29374
rect 33852 28868 33908 31276
rect 33964 30884 34020 31726
rect 34076 31220 34132 31230
rect 34188 31220 34244 33180
rect 34076 31218 34244 31220
rect 34076 31166 34078 31218
rect 34130 31166 34244 31218
rect 34076 31164 34244 31166
rect 34300 32452 34356 33180
rect 34524 32564 34580 36316
rect 34636 36260 34692 36270
rect 34636 36166 34692 36204
rect 34748 34916 34804 40910
rect 34860 40290 34916 40302
rect 34860 40238 34862 40290
rect 34914 40238 34916 40290
rect 34860 36596 34916 40238
rect 34972 40292 35028 41132
rect 35196 40852 35252 40862
rect 35084 40628 35140 40638
rect 35084 40514 35140 40572
rect 35196 40626 35252 40796
rect 35196 40574 35198 40626
rect 35250 40574 35252 40626
rect 35196 40562 35252 40574
rect 35084 40462 35086 40514
rect 35138 40462 35140 40514
rect 35084 40450 35140 40462
rect 35532 40516 35588 40526
rect 35532 40422 35588 40460
rect 34972 40236 35140 40292
rect 34972 39618 35028 39630
rect 34972 39566 34974 39618
rect 35026 39566 35028 39618
rect 34972 39172 35028 39566
rect 35084 39396 35140 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35756 39844 35812 42700
rect 35980 42196 36036 42812
rect 36092 42756 36148 42766
rect 36148 42700 36260 42756
rect 36092 42662 36148 42700
rect 35980 42140 36148 42196
rect 35980 41970 36036 41982
rect 35980 41918 35982 41970
rect 36034 41918 36036 41970
rect 35980 41300 36036 41918
rect 35868 40514 35924 40526
rect 35868 40462 35870 40514
rect 35922 40462 35924 40514
rect 35868 40180 35924 40462
rect 35868 40114 35924 40124
rect 35756 39788 35924 39844
rect 35756 39620 35812 39630
rect 35756 39526 35812 39564
rect 35196 39506 35252 39518
rect 35532 39508 35588 39518
rect 35196 39454 35198 39506
rect 35250 39454 35252 39506
rect 35196 39396 35252 39454
rect 35140 39340 35252 39396
rect 35308 39506 35588 39508
rect 35308 39454 35534 39506
rect 35586 39454 35588 39506
rect 35308 39452 35588 39454
rect 35084 39330 35140 39340
rect 35308 39172 35364 39452
rect 35532 39442 35588 39452
rect 35868 39508 35924 39788
rect 35868 39442 35924 39452
rect 34972 39106 35028 39116
rect 35084 39116 35364 39172
rect 35084 39058 35140 39116
rect 35084 39006 35086 39058
rect 35138 39006 35140 39058
rect 35084 38994 35140 39006
rect 34972 38836 35028 38846
rect 34972 38742 35028 38780
rect 35756 38836 35812 38846
rect 35980 38836 36036 41244
rect 36092 41410 36148 42140
rect 36204 42084 36260 42700
rect 36316 42530 36372 43036
rect 36316 42478 36318 42530
rect 36370 42478 36372 42530
rect 36316 42420 36372 42478
rect 36316 42354 36372 42364
rect 36204 42018 36260 42028
rect 36092 41358 36094 41410
rect 36146 41358 36148 41410
rect 36092 39620 36148 41358
rect 36316 41970 36372 41982
rect 36316 41918 36318 41970
rect 36370 41918 36372 41970
rect 36204 40962 36260 40974
rect 36204 40910 36206 40962
rect 36258 40910 36260 40962
rect 36204 40404 36260 40910
rect 36316 40516 36372 41918
rect 36428 41860 36484 41870
rect 36428 41186 36484 41804
rect 36540 41300 36596 43484
rect 37100 43428 37156 43438
rect 37100 43334 37156 43372
rect 37212 42530 37268 42542
rect 37212 42478 37214 42530
rect 37266 42478 37268 42530
rect 36652 42420 36708 42430
rect 36652 42194 36708 42364
rect 36652 42142 36654 42194
rect 36706 42142 36708 42194
rect 36652 42130 36708 42142
rect 37100 41972 37156 41982
rect 37100 41878 37156 41916
rect 36988 41860 37044 41870
rect 36988 41766 37044 41804
rect 37212 41524 37268 42478
rect 37324 41972 37380 43820
rect 39116 43540 39172 43550
rect 37996 43428 38052 43438
rect 37548 42754 37604 42766
rect 37772 42756 37828 42766
rect 37548 42702 37550 42754
rect 37602 42702 37604 42754
rect 37548 42420 37604 42702
rect 37548 42354 37604 42364
rect 37660 42754 37828 42756
rect 37660 42702 37774 42754
rect 37826 42702 37828 42754
rect 37660 42700 37828 42702
rect 37436 41972 37492 41982
rect 37324 41970 37492 41972
rect 37324 41918 37438 41970
rect 37490 41918 37492 41970
rect 37324 41916 37492 41918
rect 37436 41906 37492 41916
rect 36540 41234 36596 41244
rect 37100 41468 37268 41524
rect 36428 41134 36430 41186
rect 36482 41134 36484 41186
rect 36428 41122 36484 41134
rect 36316 40450 36372 40460
rect 36764 40626 36820 40638
rect 36764 40574 36766 40626
rect 36818 40574 36820 40626
rect 36764 40516 36820 40574
rect 36764 40450 36820 40460
rect 36204 40338 36260 40348
rect 36876 40292 36932 40302
rect 36876 40198 36932 40236
rect 36988 39844 37044 39854
rect 36092 39554 36148 39564
rect 36540 39842 37044 39844
rect 36540 39790 36990 39842
rect 37042 39790 37044 39842
rect 36540 39788 37044 39790
rect 35756 38834 36036 38836
rect 35756 38782 35758 38834
rect 35810 38782 36036 38834
rect 35756 38780 36036 38782
rect 36092 39394 36148 39406
rect 36092 39342 36094 39394
rect 36146 39342 36148 39394
rect 35084 38724 35140 38734
rect 34972 38388 35028 38398
rect 34972 38050 35028 38332
rect 35084 38276 35140 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 38276 35252 38286
rect 35084 38274 35252 38276
rect 35084 38222 35198 38274
rect 35250 38222 35252 38274
rect 35084 38220 35252 38222
rect 35196 38210 35252 38220
rect 35756 38164 35812 38780
rect 34972 37998 34974 38050
rect 35026 37998 35028 38050
rect 34972 37044 35028 37998
rect 35420 38108 35812 38164
rect 35308 37268 35364 37278
rect 35420 37268 35476 38108
rect 35980 38052 36036 38062
rect 35980 37958 36036 37996
rect 36092 38050 36148 39342
rect 36540 38946 36596 39788
rect 36988 39778 37044 39788
rect 37100 39620 37156 41468
rect 37212 41300 37268 41310
rect 37212 41206 37268 41244
rect 37660 40404 37716 42700
rect 37772 42690 37828 42700
rect 37996 42754 38052 43372
rect 38444 42980 38500 42990
rect 38444 42886 38500 42924
rect 39116 42978 39172 43484
rect 39228 43426 39284 43932
rect 39900 43988 39956 43998
rect 39900 43650 39956 43932
rect 40124 43876 40180 44270
rect 40908 44210 40964 44222
rect 40908 44158 40910 44210
rect 40962 44158 40964 44210
rect 40124 43708 40180 43820
rect 40460 44100 40516 44110
rect 40124 43652 40292 43708
rect 39900 43598 39902 43650
rect 39954 43598 39956 43650
rect 39900 43586 39956 43598
rect 39228 43374 39230 43426
rect 39282 43374 39284 43426
rect 39228 43362 39284 43374
rect 39452 43538 39508 43550
rect 39452 43486 39454 43538
rect 39506 43486 39508 43538
rect 39452 43092 39508 43486
rect 40012 43538 40068 43550
rect 40012 43486 40014 43538
rect 40066 43486 40068 43538
rect 39676 43428 39732 43438
rect 39676 43334 39732 43372
rect 39452 43026 39508 43036
rect 39564 43316 39620 43326
rect 39116 42926 39118 42978
rect 39170 42926 39172 42978
rect 39116 42914 39172 42926
rect 39452 42868 39508 42878
rect 39564 42868 39620 43260
rect 39452 42866 39620 42868
rect 39452 42814 39454 42866
rect 39506 42814 39620 42866
rect 39452 42812 39620 42814
rect 39452 42802 39508 42812
rect 37996 42702 37998 42754
rect 38050 42702 38052 42754
rect 37996 42690 38052 42702
rect 38556 42754 38612 42766
rect 38556 42702 38558 42754
rect 38610 42702 38612 42754
rect 37884 42532 37940 42542
rect 37884 42438 37940 42476
rect 38220 41858 38276 41870
rect 38220 41806 38222 41858
rect 38274 41806 38276 41858
rect 38220 41188 38276 41806
rect 38220 41122 38276 41132
rect 38556 41860 38612 42702
rect 37660 40338 37716 40348
rect 37884 40516 37940 40526
rect 37884 40402 37940 40460
rect 37884 40350 37886 40402
rect 37938 40350 37940 40402
rect 37884 40338 37940 40350
rect 38332 40404 38388 40414
rect 37212 40290 37268 40302
rect 37212 40238 37214 40290
rect 37266 40238 37268 40290
rect 37212 39844 37268 40238
rect 37772 40292 37828 40302
rect 37324 39844 37380 39854
rect 37212 39842 37380 39844
rect 37212 39790 37326 39842
rect 37378 39790 37380 39842
rect 37212 39788 37380 39790
rect 37324 39778 37380 39788
rect 37772 39732 37828 40236
rect 38108 40292 38164 40302
rect 38108 40198 38164 40236
rect 38332 40180 38388 40348
rect 38556 40180 38612 41804
rect 38780 42754 38836 42766
rect 38780 42702 38782 42754
rect 38834 42702 38836 42754
rect 38780 40516 38836 42702
rect 39004 42756 39060 42766
rect 39004 42754 39172 42756
rect 39004 42702 39006 42754
rect 39058 42702 39172 42754
rect 39004 42700 39172 42702
rect 39004 42690 39060 42700
rect 38780 40450 38836 40460
rect 38892 40964 38948 40974
rect 38892 40404 38948 40908
rect 38892 40310 38948 40348
rect 39116 40402 39172 42700
rect 40012 41972 40068 43486
rect 40012 40740 40068 41916
rect 40012 40674 40068 40684
rect 40124 42980 40180 42990
rect 40124 42644 40180 42924
rect 39116 40350 39118 40402
rect 39170 40350 39172 40402
rect 39004 40180 39060 40190
rect 38556 40124 38724 40180
rect 38332 40114 38388 40124
rect 37772 39730 38276 39732
rect 37772 39678 37774 39730
rect 37826 39678 38276 39730
rect 37772 39676 38276 39678
rect 37772 39666 37828 39676
rect 36540 38894 36542 38946
rect 36594 38894 36596 38946
rect 36540 38882 36596 38894
rect 36876 39564 37156 39620
rect 36092 37998 36094 38050
rect 36146 37998 36148 38050
rect 36092 37986 36148 37998
rect 35532 37940 35588 37950
rect 35868 37940 35924 37950
rect 35532 37938 35924 37940
rect 35532 37886 35534 37938
rect 35586 37886 35870 37938
rect 35922 37886 35924 37938
rect 35532 37884 35924 37886
rect 35532 37874 35588 37884
rect 35868 37874 35924 37884
rect 36428 37940 36484 37950
rect 36428 37846 36484 37884
rect 35308 37266 35476 37268
rect 35308 37214 35310 37266
rect 35362 37214 35476 37266
rect 35308 37212 35476 37214
rect 36092 37828 36148 37838
rect 35308 37202 35364 37212
rect 35980 37156 36036 37166
rect 34972 36978 35028 36988
rect 35868 37154 36036 37156
rect 35868 37102 35982 37154
rect 36034 37102 36036 37154
rect 35868 37100 36036 37102
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 34860 36530 34916 36540
rect 34972 36484 35028 36494
rect 35644 36484 35700 36494
rect 34972 36482 35252 36484
rect 34972 36430 34974 36482
rect 35026 36430 35252 36482
rect 34972 36428 35252 36430
rect 34972 36418 35028 36428
rect 35196 36372 35252 36428
rect 35700 36428 35812 36484
rect 35644 36418 35700 36428
rect 35308 36372 35364 36382
rect 35196 36370 35364 36372
rect 35196 36318 35310 36370
rect 35362 36318 35364 36370
rect 35196 36316 35364 36318
rect 34860 36258 34916 36270
rect 34860 36206 34862 36258
rect 34914 36206 34916 36258
rect 34860 35140 34916 36206
rect 35196 35476 35252 36316
rect 35308 36036 35364 36316
rect 35308 35970 35364 35980
rect 35420 36258 35476 36270
rect 35420 36206 35422 36258
rect 35474 36206 35476 36258
rect 35420 35924 35476 36206
rect 35420 35858 35476 35868
rect 35644 36258 35700 36270
rect 35644 36206 35646 36258
rect 35698 36206 35700 36258
rect 35084 35420 35252 35476
rect 35084 35140 35140 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35532 35140 35588 35150
rect 35644 35140 35700 36206
rect 35084 35084 35252 35140
rect 34860 35074 34916 35084
rect 34748 34914 35140 34916
rect 34748 34862 34750 34914
rect 34802 34862 35140 34914
rect 34748 34860 35140 34862
rect 34748 34850 34804 34860
rect 34860 34244 34916 34254
rect 34860 34150 34916 34188
rect 34636 34132 34692 34142
rect 34636 33236 34692 34076
rect 35084 34020 35140 34860
rect 35196 34242 35252 35084
rect 35532 35138 35700 35140
rect 35532 35086 35534 35138
rect 35586 35086 35700 35138
rect 35532 35084 35700 35086
rect 35532 35074 35588 35084
rect 35644 34916 35700 34926
rect 35532 34804 35588 34814
rect 35532 34354 35588 34748
rect 35532 34302 35534 34354
rect 35586 34302 35588 34354
rect 35532 34290 35588 34302
rect 35644 34356 35700 34860
rect 35644 34290 35700 34300
rect 35756 34356 35812 36428
rect 35868 35026 35924 37100
rect 35980 37090 36036 37100
rect 35980 35586 36036 35598
rect 35980 35534 35982 35586
rect 36034 35534 36036 35586
rect 35980 35476 36036 35534
rect 35980 35410 36036 35420
rect 36092 35138 36148 37772
rect 36876 37492 36932 39564
rect 37212 39508 37268 39518
rect 37100 39396 37156 39406
rect 37212 39396 37268 39452
rect 37100 39394 37268 39396
rect 37100 39342 37102 39394
rect 37154 39342 37268 39394
rect 37100 39340 37268 39342
rect 37100 39330 37156 39340
rect 38220 38836 38276 39676
rect 38668 39618 38724 40124
rect 39004 40086 39060 40124
rect 38668 39566 38670 39618
rect 38722 39566 38724 39618
rect 38668 39554 38724 39566
rect 38780 39508 38836 39518
rect 38780 39414 38836 39452
rect 39116 39508 39172 40350
rect 39116 39442 39172 39452
rect 39340 40402 39396 40414
rect 39340 40350 39342 40402
rect 39394 40350 39396 40402
rect 38332 39396 38388 39406
rect 38332 39394 38612 39396
rect 38332 39342 38334 39394
rect 38386 39342 38612 39394
rect 38332 39340 38612 39342
rect 38332 39330 38388 39340
rect 37884 38050 37940 38062
rect 37884 37998 37886 38050
rect 37938 37998 37940 38050
rect 37324 37940 37380 37950
rect 37324 37938 37828 37940
rect 37324 37886 37326 37938
rect 37378 37886 37828 37938
rect 37324 37884 37828 37886
rect 37324 37874 37380 37884
rect 37212 37828 37268 37838
rect 37212 37734 37268 37772
rect 37772 37492 37828 37884
rect 37884 37828 37940 37998
rect 37884 37762 37940 37772
rect 37772 37436 38164 37492
rect 36876 37426 36932 37436
rect 36876 37156 36932 37166
rect 36204 36932 36260 36942
rect 36204 36594 36260 36876
rect 36204 36542 36206 36594
rect 36258 36542 36260 36594
rect 36204 36530 36260 36542
rect 36428 36370 36484 36382
rect 36428 36318 36430 36370
rect 36482 36318 36484 36370
rect 36428 35252 36484 36318
rect 36652 35812 36708 35822
rect 36652 35698 36708 35756
rect 36652 35646 36654 35698
rect 36706 35646 36708 35698
rect 36652 35634 36708 35646
rect 36876 35698 36932 37100
rect 38108 37154 38164 37436
rect 38108 37102 38110 37154
rect 38162 37102 38164 37154
rect 38108 37090 38164 37102
rect 38220 36932 38276 38780
rect 38556 38724 38612 39340
rect 39340 39284 39396 40350
rect 39452 40404 39508 40414
rect 39452 40402 39956 40404
rect 39452 40350 39454 40402
rect 39506 40350 39956 40402
rect 39452 40348 39956 40350
rect 39452 40338 39508 40348
rect 39340 39218 39396 39228
rect 39900 39060 39956 40348
rect 40124 40402 40180 42588
rect 40124 40350 40126 40402
rect 40178 40350 40180 40402
rect 40124 40338 40180 40350
rect 40236 40404 40292 43652
rect 40348 41860 40404 41870
rect 40348 41766 40404 41804
rect 40348 40628 40404 40638
rect 40460 40628 40516 44044
rect 40908 43708 40964 44158
rect 41468 44212 41524 44222
rect 40796 43652 40964 43708
rect 41356 43988 41412 43998
rect 40348 40626 40516 40628
rect 40348 40574 40350 40626
rect 40402 40574 40516 40626
rect 40348 40572 40516 40574
rect 40572 40740 40628 40750
rect 40348 40562 40404 40572
rect 40236 40338 40292 40348
rect 40348 40292 40404 40302
rect 40012 39060 40068 39070
rect 39900 39058 40068 39060
rect 39900 39006 40014 39058
rect 40066 39006 40068 39058
rect 39900 39004 40068 39006
rect 40012 38994 40068 39004
rect 40236 38946 40292 38958
rect 40236 38894 40238 38946
rect 40290 38894 40292 38946
rect 39116 38834 39172 38846
rect 39116 38782 39118 38834
rect 39170 38782 39172 38834
rect 38668 38724 38724 38734
rect 38556 38722 38724 38724
rect 38556 38670 38670 38722
rect 38722 38670 38724 38722
rect 38556 38668 38724 38670
rect 38668 38612 39060 38668
rect 38332 38052 38388 38062
rect 38332 37958 38388 37996
rect 38892 38050 38948 38062
rect 38892 37998 38894 38050
rect 38946 37998 38948 38050
rect 38556 37938 38612 37950
rect 38556 37886 38558 37938
rect 38610 37886 38612 37938
rect 37996 36876 38276 36932
rect 38444 37492 38500 37502
rect 37996 36594 38052 36876
rect 37996 36542 37998 36594
rect 38050 36542 38052 36594
rect 37996 36530 38052 36542
rect 37212 36484 37268 36494
rect 37100 36036 37156 36046
rect 36988 35924 37044 35934
rect 36988 35830 37044 35868
rect 36876 35646 36878 35698
rect 36930 35646 36932 35698
rect 36876 35634 36932 35646
rect 36428 35186 36484 35196
rect 36092 35086 36094 35138
rect 36146 35086 36148 35138
rect 36092 35074 36148 35086
rect 35868 34974 35870 35026
rect 35922 34974 35924 35026
rect 35868 34962 35924 34974
rect 36316 35028 36372 35038
rect 36316 34934 36372 34972
rect 36988 34804 37044 34814
rect 36988 34710 37044 34748
rect 35756 34300 36036 34356
rect 35196 34190 35198 34242
rect 35250 34190 35252 34242
rect 35196 34178 35252 34190
rect 35308 34242 35364 34254
rect 35308 34190 35310 34242
rect 35362 34190 35364 34242
rect 35308 34132 35364 34190
rect 35756 34132 35812 34300
rect 35308 34076 35812 34132
rect 35868 34132 35924 34142
rect 35868 34038 35924 34076
rect 34972 33964 35140 34020
rect 34748 33906 34804 33918
rect 34748 33854 34750 33906
rect 34802 33854 34804 33906
rect 34748 33796 34804 33854
rect 34748 33730 34804 33740
rect 34860 33458 34916 33470
rect 34860 33406 34862 33458
rect 34914 33406 34916 33458
rect 34860 33236 34916 33406
rect 34636 33180 34916 33236
rect 34524 32498 34580 32508
rect 34748 32562 34804 32574
rect 34748 32510 34750 32562
rect 34802 32510 34804 32562
rect 34300 31778 34356 32396
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34076 31154 34132 31164
rect 33964 30818 34020 30828
rect 34300 30436 34356 31726
rect 34188 30380 34356 30436
rect 34412 31892 34468 31902
rect 34076 29428 34132 29438
rect 33852 28802 33908 28812
rect 33964 29426 34132 29428
rect 33964 29374 34078 29426
rect 34130 29374 34132 29426
rect 33964 29372 34132 29374
rect 33740 28690 33796 28700
rect 33516 28018 33572 28028
rect 33180 27858 33460 27860
rect 33180 27806 33182 27858
rect 33234 27806 33460 27858
rect 33180 27804 33460 27806
rect 33180 27794 33236 27804
rect 32508 27094 32564 27132
rect 32844 27468 33012 27524
rect 33068 27748 33124 27758
rect 32396 26338 32452 26348
rect 32396 26178 32452 26190
rect 32396 26126 32398 26178
rect 32450 26126 32452 26178
rect 32172 26068 32228 26078
rect 32172 25618 32228 26012
rect 32396 25844 32452 26126
rect 32396 25788 32676 25844
rect 32172 25566 32174 25618
rect 32226 25566 32228 25618
rect 32172 25554 32228 25566
rect 32060 25508 32116 25518
rect 31948 25506 32116 25508
rect 31948 25454 32062 25506
rect 32114 25454 32116 25506
rect 31948 25452 32116 25454
rect 31724 25394 31780 25406
rect 31724 25342 31726 25394
rect 31778 25342 31780 25394
rect 31724 24612 31780 25342
rect 31948 25396 32004 25452
rect 32060 25442 32116 25452
rect 32508 25508 32564 25518
rect 32620 25508 32676 25788
rect 32732 25508 32788 25518
rect 32620 25452 32732 25508
rect 32508 25414 32564 25452
rect 32732 25414 32788 25452
rect 31948 25330 32004 25340
rect 32284 25284 32340 25294
rect 32284 25190 32340 25228
rect 31724 24546 31780 24556
rect 32508 24612 32564 24622
rect 32508 24518 32564 24556
rect 31836 24500 31892 24510
rect 31836 24050 31892 24444
rect 31836 23998 31838 24050
rect 31890 23998 31892 24050
rect 31836 23986 31892 23998
rect 31612 23492 31780 23548
rect 31388 23324 31556 23380
rect 31388 22260 31444 22270
rect 31276 22204 31388 22260
rect 30940 21970 30996 21980
rect 30716 21644 31220 21700
rect 30156 20738 30212 20748
rect 30268 21362 30436 21364
rect 30268 21310 30382 21362
rect 30434 21310 30436 21362
rect 30268 21308 30436 21310
rect 30044 20580 30100 20590
rect 30044 20242 30100 20524
rect 30268 20580 30324 21308
rect 30380 21298 30436 21308
rect 30604 21474 30660 21486
rect 30604 21422 30606 21474
rect 30658 21422 30660 21474
rect 30604 21364 30660 21422
rect 30604 21298 30660 21308
rect 30716 20692 30772 20702
rect 30716 20598 30772 20636
rect 30268 20514 30324 20524
rect 30380 20578 30436 20590
rect 30380 20526 30382 20578
rect 30434 20526 30436 20578
rect 30044 20190 30046 20242
rect 30098 20190 30100 20242
rect 30044 20178 30100 20190
rect 30380 19908 30436 20526
rect 30828 20580 30884 20590
rect 30828 20486 30884 20524
rect 30940 20356 30996 21644
rect 31164 21586 31220 21644
rect 31164 21534 31166 21586
rect 31218 21534 31220 21586
rect 31164 21522 31220 21534
rect 31388 21588 31444 22204
rect 31388 20802 31444 21532
rect 31500 21812 31556 23324
rect 31724 23268 31780 23492
rect 31724 23202 31780 23212
rect 31612 23154 31668 23166
rect 31612 23102 31614 23154
rect 31666 23102 31668 23154
rect 31612 21924 31668 23102
rect 31836 23154 31892 23166
rect 31836 23102 31838 23154
rect 31890 23102 31892 23154
rect 31724 23044 31780 23054
rect 31724 22950 31780 22988
rect 31836 22484 31892 23102
rect 32396 23156 32452 23166
rect 32396 23062 32452 23100
rect 31836 22418 31892 22428
rect 31612 21858 31668 21868
rect 31948 22036 32004 22046
rect 31500 21586 31556 21756
rect 31500 21534 31502 21586
rect 31554 21534 31556 21586
rect 31500 21522 31556 21534
rect 31724 21476 31780 21486
rect 31724 21474 31892 21476
rect 31724 21422 31726 21474
rect 31778 21422 31892 21474
rect 31724 21420 31892 21422
rect 31724 21410 31780 21420
rect 31388 20750 31390 20802
rect 31442 20750 31444 20802
rect 31388 20738 31444 20750
rect 30716 20300 30996 20356
rect 30716 20242 30772 20300
rect 30716 20190 30718 20242
rect 30770 20190 30772 20242
rect 30716 20178 30772 20190
rect 31724 20244 31780 20254
rect 31724 20150 31780 20188
rect 31836 20020 31892 21420
rect 29932 19182 29934 19234
rect 29986 19182 29988 19234
rect 29932 19170 29988 19182
rect 30268 19852 30380 19908
rect 29316 18956 29428 19012
rect 29260 18918 29316 18956
rect 30044 18564 30100 18574
rect 30044 18470 30100 18508
rect 29148 17890 29204 18396
rect 29596 18450 29652 18462
rect 29596 18398 29598 18450
rect 29650 18398 29652 18450
rect 29148 17838 29150 17890
rect 29202 17838 29204 17890
rect 29148 17826 29204 17838
rect 29260 18340 29316 18350
rect 29596 18340 29652 18398
rect 29260 18338 29652 18340
rect 29260 18286 29262 18338
rect 29314 18286 29652 18338
rect 29260 18284 29652 18286
rect 29820 18450 29876 18462
rect 29820 18398 29822 18450
rect 29874 18398 29876 18450
rect 29260 15540 29316 18284
rect 29484 17780 29540 17790
rect 29820 17780 29876 18398
rect 30156 18452 30212 18462
rect 30156 18358 30212 18396
rect 29932 18340 29988 18350
rect 29932 18246 29988 18284
rect 29484 17778 29876 17780
rect 29484 17726 29486 17778
rect 29538 17726 29876 17778
rect 29484 17724 29876 17726
rect 29484 17714 29540 17724
rect 29820 17666 29876 17724
rect 29820 17614 29822 17666
rect 29874 17614 29876 17666
rect 29820 17602 29876 17614
rect 29484 17556 29540 17566
rect 29372 17444 29428 17454
rect 29484 17444 29540 17500
rect 30156 17444 30212 17454
rect 29372 17442 29540 17444
rect 29372 17390 29374 17442
rect 29426 17390 29540 17442
rect 29372 17388 29540 17390
rect 29708 17442 30212 17444
rect 29708 17390 30158 17442
rect 30210 17390 30212 17442
rect 29708 17388 30212 17390
rect 29372 17378 29428 17388
rect 29484 16212 29540 16222
rect 29484 16098 29540 16156
rect 29484 16046 29486 16098
rect 29538 16046 29540 16098
rect 29484 16034 29540 16046
rect 29708 16100 29764 17388
rect 30156 17378 30212 17388
rect 30268 16772 30324 19852
rect 30380 19842 30436 19852
rect 31276 19908 31332 19918
rect 31276 19906 31780 19908
rect 31276 19854 31278 19906
rect 31330 19854 31780 19906
rect 31276 19852 31780 19854
rect 31276 19842 31332 19852
rect 31164 19796 31220 19806
rect 30828 19794 31220 19796
rect 30828 19742 31166 19794
rect 31218 19742 31220 19794
rect 30828 19740 31220 19742
rect 30716 19348 30772 19358
rect 30828 19348 30884 19740
rect 31164 19730 31220 19740
rect 30716 19346 30884 19348
rect 30716 19294 30718 19346
rect 30770 19294 30884 19346
rect 30716 19292 30884 19294
rect 30716 19282 30772 19292
rect 31724 18674 31780 19852
rect 31724 18622 31726 18674
rect 31778 18622 31780 18674
rect 31724 18610 31780 18622
rect 31836 18674 31892 19964
rect 31836 18622 31838 18674
rect 31890 18622 31892 18674
rect 31836 18610 31892 18622
rect 30716 18564 30772 18574
rect 30716 18340 30772 18508
rect 30716 18246 30772 18284
rect 30828 18452 30884 18462
rect 30828 17666 30884 18396
rect 31500 18452 31556 18462
rect 31500 18358 31556 18396
rect 31612 18450 31668 18462
rect 31948 18452 32004 21980
rect 32060 21812 32116 21822
rect 32060 21718 32116 21756
rect 32396 21698 32452 21710
rect 32396 21646 32398 21698
rect 32450 21646 32452 21698
rect 32172 20916 32228 20926
rect 32060 20860 32172 20916
rect 32060 20802 32116 20860
rect 32172 20850 32228 20860
rect 32060 20750 32062 20802
rect 32114 20750 32116 20802
rect 32060 20738 32116 20750
rect 32396 20132 32452 21646
rect 32060 19348 32116 19358
rect 32060 18562 32116 19292
rect 32060 18510 32062 18562
rect 32114 18510 32116 18562
rect 32060 18498 32116 18510
rect 31612 18398 31614 18450
rect 31666 18398 31668 18450
rect 31388 18004 31444 18014
rect 31388 17778 31444 17948
rect 31388 17726 31390 17778
rect 31442 17726 31444 17778
rect 31388 17714 31444 17726
rect 30828 17614 30830 17666
rect 30882 17614 30884 17666
rect 30828 17602 30884 17614
rect 31500 17668 31556 17678
rect 29932 16716 30268 16772
rect 29708 16098 29876 16100
rect 29708 16046 29710 16098
rect 29762 16046 29876 16098
rect 29708 16044 29876 16046
rect 29708 16034 29764 16044
rect 29820 15652 29876 16044
rect 29932 16098 29988 16716
rect 30268 16678 30324 16716
rect 30492 17442 30548 17454
rect 30492 17390 30494 17442
rect 30546 17390 30548 17442
rect 30492 16436 30548 17390
rect 31388 17108 31444 17118
rect 31276 16882 31332 16894
rect 31276 16830 31278 16882
rect 31330 16830 31332 16882
rect 30492 16370 30548 16380
rect 30604 16770 30660 16782
rect 30604 16718 30606 16770
rect 30658 16718 30660 16770
rect 30604 16322 30660 16718
rect 30604 16270 30606 16322
rect 30658 16270 30660 16322
rect 30604 16258 30660 16270
rect 30044 16212 30100 16222
rect 30492 16212 30548 16222
rect 30044 16210 30548 16212
rect 30044 16158 30046 16210
rect 30098 16158 30494 16210
rect 30546 16158 30548 16210
rect 30044 16156 30548 16158
rect 30044 16146 30100 16156
rect 30492 16146 30548 16156
rect 29932 16046 29934 16098
rect 29986 16046 29988 16098
rect 29932 16034 29988 16046
rect 30044 15988 30100 15998
rect 30044 15894 30100 15932
rect 29820 15596 30100 15652
rect 28588 14914 28644 14924
rect 28700 15092 28868 15148
rect 28924 15092 29092 15148
rect 29148 15484 29316 15540
rect 28476 14532 28532 14542
rect 28476 14438 28532 14476
rect 28700 14084 28756 15092
rect 28476 13746 28532 13758
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28476 13188 28532 13694
rect 28476 13122 28532 13132
rect 28588 12852 28644 12862
rect 28588 12758 28644 12796
rect 28476 12068 28532 12078
rect 28476 11974 28532 12012
rect 28588 11954 28644 11966
rect 28588 11902 28590 11954
rect 28642 11902 28644 11954
rect 28588 11620 28644 11902
rect 28588 11554 28644 11564
rect 28700 11956 28756 14028
rect 28924 13524 28980 15092
rect 29036 14306 29092 14318
rect 29036 14254 29038 14306
rect 29090 14254 29092 14306
rect 29036 13746 29092 14254
rect 29036 13694 29038 13746
rect 29090 13694 29092 13746
rect 29036 13682 29092 13694
rect 28924 13468 29092 13524
rect 28924 12964 28980 12974
rect 28364 11342 28366 11394
rect 28418 11342 28420 11394
rect 28364 11172 28420 11342
rect 28588 11396 28644 11406
rect 28700 11396 28756 11900
rect 28588 11394 28756 11396
rect 28588 11342 28590 11394
rect 28642 11342 28756 11394
rect 28588 11340 28756 11342
rect 28812 12852 28868 12862
rect 28812 11844 28868 12796
rect 28924 12290 28980 12908
rect 28924 12238 28926 12290
rect 28978 12238 28980 12290
rect 28924 12226 28980 12238
rect 28588 11330 28644 11340
rect 28812 11284 28868 11788
rect 28364 10724 28420 11116
rect 28364 10658 28420 10668
rect 28700 11228 28868 11284
rect 28476 10500 28532 10510
rect 28252 10498 28532 10500
rect 28252 10446 28478 10498
rect 28530 10446 28532 10498
rect 28252 10444 28532 10446
rect 28140 10434 28196 10444
rect 28476 10434 28532 10444
rect 27692 9938 27748 10220
rect 27692 9886 27694 9938
rect 27746 9886 27748 9938
rect 27468 8418 27524 8428
rect 27580 9044 27636 9054
rect 27356 8318 27358 8370
rect 27410 8318 27412 8370
rect 27356 8306 27412 8318
rect 26236 7534 26238 7586
rect 26290 7534 26292 7586
rect 26236 7522 26292 7534
rect 26348 8258 26404 8270
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 26348 7588 26404 8206
rect 27468 8260 27524 8270
rect 27580 8260 27636 8988
rect 27468 8258 27636 8260
rect 27468 8206 27470 8258
rect 27522 8206 27636 8258
rect 27468 8204 27636 8206
rect 27692 8260 27748 9886
rect 28476 10276 28532 10286
rect 28476 9940 28532 10220
rect 28588 9940 28644 9950
rect 28476 9938 28644 9940
rect 28476 9886 28590 9938
rect 28642 9886 28644 9938
rect 28476 9884 28644 9886
rect 28588 9874 28644 9884
rect 28140 9604 28196 9614
rect 28140 9510 28196 9548
rect 27916 9268 27972 9278
rect 27916 9174 27972 9212
rect 28700 9044 28756 11228
rect 29036 11060 29092 13468
rect 29148 13076 29204 15484
rect 29260 15202 29316 15214
rect 29260 15150 29262 15202
rect 29314 15150 29316 15202
rect 29260 14980 29316 15150
rect 29260 14914 29316 14924
rect 29820 14980 29876 14990
rect 29372 14756 29428 14766
rect 29708 14756 29764 14766
rect 29372 14530 29428 14700
rect 29372 14478 29374 14530
rect 29426 14478 29428 14530
rect 29372 14466 29428 14478
rect 29484 14700 29708 14756
rect 29484 14420 29540 14700
rect 29708 14690 29764 14700
rect 29820 14530 29876 14924
rect 29820 14478 29822 14530
rect 29874 14478 29876 14530
rect 29820 14466 29876 14478
rect 30044 14532 30100 15596
rect 31276 15316 31332 16830
rect 31388 16210 31444 17052
rect 31388 16158 31390 16210
rect 31442 16158 31444 16210
rect 31388 16146 31444 16158
rect 31276 15250 31332 15260
rect 31388 15202 31444 15214
rect 31388 15150 31390 15202
rect 31442 15150 31444 15202
rect 31388 15148 31444 15150
rect 31052 15092 31444 15148
rect 30380 14644 30436 14682
rect 30380 14578 30436 14588
rect 30828 14644 30884 14654
rect 30828 14550 30884 14588
rect 30940 14644 30996 14654
rect 31052 14644 31108 15092
rect 31500 14868 31556 17612
rect 30940 14642 31108 14644
rect 30940 14590 30942 14642
rect 30994 14590 31108 14642
rect 30940 14588 31108 14590
rect 31164 14812 31556 14868
rect 30940 14578 30996 14588
rect 30044 14530 30212 14532
rect 30044 14478 30046 14530
rect 30098 14478 30212 14530
rect 30044 14476 30212 14478
rect 30044 14466 30100 14476
rect 29260 14308 29316 14318
rect 29260 14214 29316 14252
rect 29148 13010 29204 13020
rect 29260 12850 29316 12862
rect 29260 12798 29262 12850
rect 29314 12798 29316 12850
rect 29260 12404 29316 12798
rect 29372 12852 29428 12862
rect 29372 12758 29428 12796
rect 29260 12338 29316 12348
rect 29148 12292 29204 12302
rect 29148 12198 29204 12236
rect 29372 12178 29428 12190
rect 29372 12126 29374 12178
rect 29426 12126 29428 12178
rect 29260 12068 29316 12078
rect 29260 11974 29316 12012
rect 29372 11844 29428 12126
rect 29372 11778 29428 11788
rect 29036 10994 29092 11004
rect 29484 10836 29540 14364
rect 29596 13972 29652 13982
rect 29596 13970 30100 13972
rect 29596 13918 29598 13970
rect 29650 13918 30100 13970
rect 29596 13916 30100 13918
rect 29596 13906 29652 13916
rect 29820 13746 29876 13758
rect 29820 13694 29822 13746
rect 29874 13694 29876 13746
rect 29820 13524 29876 13694
rect 30044 13746 30100 13916
rect 30044 13694 30046 13746
rect 30098 13694 30100 13746
rect 30044 13682 30100 13694
rect 29820 13458 29876 13468
rect 29708 13188 29764 13198
rect 29708 13076 29764 13132
rect 29708 13074 29988 13076
rect 29708 13022 29710 13074
rect 29762 13022 29988 13074
rect 29708 13020 29988 13022
rect 29708 13010 29764 13020
rect 29596 12516 29652 12526
rect 29596 12178 29652 12460
rect 29932 12290 29988 13020
rect 29932 12238 29934 12290
rect 29986 12238 29988 12290
rect 29932 12226 29988 12238
rect 30156 12402 30212 14476
rect 30380 14420 30436 14430
rect 30940 14420 30996 14430
rect 30436 14364 30548 14420
rect 30380 14326 30436 14364
rect 30268 14306 30324 14318
rect 30268 14254 30270 14306
rect 30322 14254 30324 14306
rect 30268 14084 30324 14254
rect 30268 14018 30324 14028
rect 30268 13860 30324 13870
rect 30268 13766 30324 13804
rect 30492 12516 30548 14364
rect 30156 12350 30158 12402
rect 30210 12350 30212 12402
rect 30156 12292 30212 12350
rect 30268 12404 30324 12414
rect 30268 12310 30324 12348
rect 30492 12402 30548 12460
rect 30492 12350 30494 12402
rect 30546 12350 30548 12402
rect 30492 12338 30548 12350
rect 30828 13746 30884 13758
rect 30828 13694 30830 13746
rect 30882 13694 30884 13746
rect 30156 12226 30212 12236
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29596 12114 29652 12126
rect 30380 12178 30436 12190
rect 30380 12126 30382 12178
rect 30434 12126 30436 12178
rect 30380 11956 30436 12126
rect 30828 12180 30884 13694
rect 30828 12114 30884 12124
rect 30828 11956 30884 11966
rect 30380 11954 30884 11956
rect 30380 11902 30830 11954
rect 30882 11902 30884 11954
rect 30380 11900 30884 11902
rect 30828 11890 30884 11900
rect 28812 10780 29540 10836
rect 30604 11620 30660 11630
rect 28812 9266 28868 10780
rect 30604 10722 30660 11564
rect 30604 10670 30606 10722
rect 30658 10670 30660 10722
rect 30604 10658 30660 10670
rect 29372 10612 29428 10622
rect 29260 10052 29316 10062
rect 29260 9826 29316 9996
rect 29260 9774 29262 9826
rect 29314 9774 29316 9826
rect 29260 9762 29316 9774
rect 28812 9214 28814 9266
rect 28866 9214 28868 9266
rect 28812 9202 28868 9214
rect 28700 8988 28868 9044
rect 28476 8932 28532 8942
rect 28476 8838 28532 8876
rect 27468 8194 27524 8204
rect 27692 8194 27748 8204
rect 27804 8372 27860 8382
rect 28140 8372 28196 8382
rect 27804 8258 27860 8316
rect 27804 8206 27806 8258
rect 27858 8206 27860 8258
rect 27804 8194 27860 8206
rect 28028 8370 28196 8372
rect 28028 8318 28142 8370
rect 28194 8318 28196 8370
rect 28028 8316 28196 8318
rect 27692 8034 27748 8046
rect 27692 7982 27694 8034
rect 27746 7982 27748 8034
rect 26348 7586 26740 7588
rect 26348 7534 26350 7586
rect 26402 7534 26740 7586
rect 26348 7532 26740 7534
rect 26348 7522 26404 7532
rect 26012 7410 26068 7420
rect 26124 7474 26180 7486
rect 26124 7422 26126 7474
rect 26178 7422 26180 7474
rect 25564 6738 25620 6748
rect 25564 6020 25620 6030
rect 25340 6018 25620 6020
rect 25340 5966 25566 6018
rect 25618 5966 25620 6018
rect 25340 5964 25620 5966
rect 25228 5908 25284 5918
rect 24780 5182 24782 5234
rect 24834 5182 24836 5234
rect 24780 5170 24836 5182
rect 25116 5852 25228 5908
rect 25116 5124 25172 5852
rect 25228 5814 25284 5852
rect 25564 5124 25620 5964
rect 26012 5908 26068 5918
rect 26124 5908 26180 7422
rect 26684 6804 26740 7532
rect 27356 7474 27412 7486
rect 27356 7422 27358 7474
rect 27410 7422 27412 7474
rect 26796 7364 26852 7374
rect 26796 7270 26852 7308
rect 26796 6804 26852 6814
rect 26684 6802 26852 6804
rect 26684 6750 26798 6802
rect 26850 6750 26852 6802
rect 26684 6748 26852 6750
rect 26796 6738 26852 6748
rect 26908 6804 26964 6814
rect 26348 6580 26404 6590
rect 26908 6580 26964 6748
rect 26236 6132 26292 6142
rect 26236 6038 26292 6076
rect 26068 5852 26180 5908
rect 26012 5842 26068 5852
rect 25676 5572 25732 5582
rect 25676 5346 25732 5516
rect 25676 5294 25678 5346
rect 25730 5294 25732 5346
rect 25676 5282 25732 5294
rect 26348 5346 26404 6524
rect 26796 6524 26964 6580
rect 26572 5908 26628 5918
rect 26572 5814 26628 5852
rect 26684 5572 26740 5582
rect 26796 5572 26852 6524
rect 26740 5516 26852 5572
rect 26684 5506 26740 5516
rect 26348 5294 26350 5346
rect 26402 5294 26404 5346
rect 26348 5282 26404 5294
rect 26796 5346 26852 5516
rect 26796 5294 26798 5346
rect 26850 5294 26852 5346
rect 26796 5282 26852 5294
rect 27356 6018 27412 7422
rect 27692 6692 27748 7982
rect 28028 7586 28084 8316
rect 28140 8306 28196 8316
rect 28364 8260 28420 8270
rect 28028 7534 28030 7586
rect 28082 7534 28084 7586
rect 28028 7522 28084 7534
rect 28252 8034 28308 8046
rect 28252 7982 28254 8034
rect 28306 7982 28308 8034
rect 28252 6804 28308 7982
rect 28252 6738 28308 6748
rect 28364 7364 28420 8204
rect 28476 8148 28532 8158
rect 28476 8054 28532 8092
rect 28140 6692 28196 6702
rect 27692 6636 28140 6692
rect 28140 6598 28196 6636
rect 28364 6690 28420 7308
rect 28364 6638 28366 6690
rect 28418 6638 28420 6690
rect 28364 6626 28420 6638
rect 28588 6580 28644 6590
rect 28588 6486 28644 6524
rect 27356 5966 27358 6018
rect 27410 5966 27412 6018
rect 26012 5234 26068 5246
rect 26012 5182 26014 5234
rect 26066 5182 26068 5234
rect 25564 5068 25956 5124
rect 25116 5030 25172 5068
rect 25900 5010 25956 5068
rect 25900 4958 25902 5010
rect 25954 4958 25956 5010
rect 25900 4946 25956 4958
rect 23996 4610 24052 4620
rect 25228 4676 25284 4686
rect 24444 4452 24500 4462
rect 24444 4358 24500 4396
rect 25228 4338 25284 4620
rect 26012 4450 26068 5182
rect 26460 5236 26516 5246
rect 26460 5142 26516 5180
rect 26236 5124 26292 5134
rect 27244 5124 27300 5134
rect 26236 5012 26292 5068
rect 27020 5068 27244 5124
rect 26236 4956 26404 5012
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 23772 3614 23774 3666
rect 23826 3614 23828 3666
rect 23772 3602 23828 3614
rect 24108 4226 24164 4238
rect 24108 4174 24110 4226
rect 24162 4174 24164 4226
rect 23996 3556 24052 3566
rect 24108 3556 24164 4174
rect 24052 3500 24164 3556
rect 23996 3462 24052 3500
rect 26012 3444 26068 3454
rect 23100 3332 23156 3342
rect 24892 3332 24948 3342
rect 23100 800 23156 3276
rect 24668 3330 24948 3332
rect 24668 3278 24894 3330
rect 24946 3278 24948 3330
rect 24668 3276 24948 3278
rect 24668 800 24724 3276
rect 24892 3266 24948 3276
rect 25340 3332 25396 3342
rect 25340 3238 25396 3276
rect 26012 3330 26068 3388
rect 26348 3442 26404 4956
rect 27020 5010 27076 5068
rect 27020 4958 27022 5010
rect 27074 4958 27076 5010
rect 27020 4946 27076 4958
rect 26908 4900 26964 4910
rect 26908 4806 26964 4844
rect 27244 3780 27300 5068
rect 27356 4676 27412 5966
rect 27580 5908 27636 5918
rect 27468 5460 27524 5470
rect 27468 5234 27524 5404
rect 27468 5182 27470 5234
rect 27522 5182 27524 5234
rect 27468 5170 27524 5182
rect 27580 5348 27636 5852
rect 27580 5122 27636 5292
rect 27580 5070 27582 5122
rect 27634 5070 27636 5122
rect 27580 5058 27636 5070
rect 27804 5124 27860 5134
rect 27804 5030 27860 5068
rect 27356 4610 27412 4620
rect 28588 4676 28644 4686
rect 28588 4340 28644 4620
rect 28812 4340 28868 8988
rect 29260 8932 29316 8942
rect 29372 8932 29428 10556
rect 30604 10500 30660 10510
rect 29932 9716 29988 9726
rect 29932 9714 30548 9716
rect 29932 9662 29934 9714
rect 29986 9662 30548 9714
rect 29932 9660 30548 9662
rect 29932 9650 29988 9660
rect 30492 9266 30548 9660
rect 30492 9214 30494 9266
rect 30546 9214 30548 9266
rect 30492 9202 30548 9214
rect 30156 9156 30212 9166
rect 30156 9062 30212 9100
rect 30604 9154 30660 10444
rect 30940 9604 30996 14364
rect 31052 12066 31108 12078
rect 31052 12014 31054 12066
rect 31106 12014 31108 12066
rect 31052 11956 31108 12014
rect 31164 11956 31220 14812
rect 31612 14644 31668 18398
rect 31724 18396 32004 18452
rect 32396 18452 32452 20076
rect 32844 19572 32900 27468
rect 33068 27188 33124 27692
rect 33292 27300 33348 27310
rect 33292 27206 33348 27244
rect 33180 27188 33236 27198
rect 33068 27186 33236 27188
rect 33068 27134 33182 27186
rect 33234 27134 33236 27186
rect 33068 27132 33236 27134
rect 33180 27122 33236 27132
rect 32956 26404 33012 26414
rect 32956 25284 33012 26348
rect 33404 26290 33460 27804
rect 33852 27746 33908 27758
rect 33852 27694 33854 27746
rect 33906 27694 33908 27746
rect 33852 27300 33908 27694
rect 33852 27234 33908 27244
rect 33404 26238 33406 26290
rect 33458 26238 33460 26290
rect 33404 26226 33460 26238
rect 33740 27076 33796 27086
rect 33964 27076 34020 29372
rect 34076 29362 34132 29372
rect 34076 28756 34132 28766
rect 34076 27300 34132 28700
rect 34188 28532 34244 30380
rect 34300 30212 34356 30222
rect 34412 30212 34468 31836
rect 34748 30884 34804 32510
rect 34860 31778 34916 31790
rect 34860 31726 34862 31778
rect 34914 31726 34916 31778
rect 34860 31332 34916 31726
rect 34860 31266 34916 31276
rect 34748 30818 34804 30828
rect 34300 30210 34468 30212
rect 34300 30158 34302 30210
rect 34354 30158 34468 30210
rect 34300 30156 34468 30158
rect 34300 30146 34356 30156
rect 34188 28476 34356 28532
rect 34076 27234 34132 27244
rect 34188 28308 34244 28318
rect 34188 27186 34244 28252
rect 34188 27134 34190 27186
rect 34242 27134 34244 27186
rect 34188 27122 34244 27134
rect 33740 27074 34020 27076
rect 33740 27022 33742 27074
rect 33794 27022 34020 27074
rect 33740 27020 34020 27022
rect 33180 25844 33236 25854
rect 33180 25618 33236 25788
rect 33180 25566 33182 25618
rect 33234 25566 33236 25618
rect 33180 25554 33236 25566
rect 32956 25218 33012 25228
rect 33628 25284 33684 25294
rect 33628 25190 33684 25228
rect 31724 17892 31780 18396
rect 32396 18386 32452 18396
rect 32508 19516 32900 19572
rect 32956 23828 33012 23838
rect 32508 18452 32564 19516
rect 32844 19348 32900 19358
rect 32844 19254 32900 19292
rect 32956 19124 33012 23772
rect 33740 23828 33796 27020
rect 34300 26908 34356 28476
rect 34076 26852 34356 26908
rect 34412 26908 34468 30156
rect 34860 30210 34916 30222
rect 34860 30158 34862 30210
rect 34914 30158 34916 30210
rect 34860 29876 34916 30158
rect 34860 29810 34916 29820
rect 34972 29540 35028 33964
rect 35868 33908 35924 33918
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 33572 35252 33582
rect 35252 33516 35476 33572
rect 35196 33506 35252 33516
rect 35084 33460 35140 33470
rect 35084 33236 35140 33404
rect 35420 33348 35476 33516
rect 35420 33346 35812 33348
rect 35420 33294 35422 33346
rect 35474 33294 35812 33346
rect 35420 33292 35812 33294
rect 35420 33282 35476 33292
rect 35196 33236 35252 33246
rect 35084 33234 35252 33236
rect 35084 33182 35198 33234
rect 35250 33182 35252 33234
rect 35084 33180 35252 33182
rect 35084 33124 35140 33180
rect 35196 33170 35252 33180
rect 35084 33058 35140 33068
rect 35420 32452 35476 32462
rect 35420 32450 35700 32452
rect 35420 32398 35422 32450
rect 35474 32398 35700 32450
rect 35420 32396 35700 32398
rect 35420 32386 35476 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35644 31890 35700 32396
rect 35644 31838 35646 31890
rect 35698 31838 35700 31890
rect 35644 31826 35700 31838
rect 35756 31892 35812 33292
rect 35868 32228 35924 33852
rect 35980 32564 36036 34300
rect 36540 34244 36596 34254
rect 36540 34150 36596 34188
rect 36204 33236 36260 33246
rect 36204 33142 36260 33180
rect 36988 33236 37044 33246
rect 37100 33236 37156 35980
rect 37212 35698 37268 36428
rect 38444 36482 38500 37436
rect 38444 36430 38446 36482
rect 38498 36430 38500 36482
rect 37212 35646 37214 35698
rect 37266 35646 37268 35698
rect 37212 35634 37268 35646
rect 37548 35700 37604 35710
rect 37548 35698 37716 35700
rect 37548 35646 37550 35698
rect 37602 35646 37716 35698
rect 37548 35644 37716 35646
rect 37548 35634 37604 35644
rect 37548 35140 37604 35150
rect 37548 35046 37604 35084
rect 37212 34916 37268 34926
rect 37212 34356 37268 34860
rect 37212 34290 37268 34300
rect 37324 34802 37380 34814
rect 37324 34750 37326 34802
rect 37378 34750 37380 34802
rect 37324 34244 37380 34750
rect 37324 34178 37380 34188
rect 37660 34132 37716 35644
rect 38220 35586 38276 35598
rect 38220 35534 38222 35586
rect 38274 35534 38276 35586
rect 37772 35252 37828 35262
rect 37828 35196 37940 35252
rect 37772 35186 37828 35196
rect 37660 34066 37716 34076
rect 37772 35028 37828 35038
rect 37772 34914 37828 34972
rect 37772 34862 37774 34914
rect 37826 34862 37828 34914
rect 36988 33234 37156 33236
rect 36988 33182 36990 33234
rect 37042 33182 37156 33234
rect 36988 33180 37156 33182
rect 37212 33346 37268 33358
rect 37212 33294 37214 33346
rect 37266 33294 37268 33346
rect 36988 33170 37044 33180
rect 36092 33122 36148 33134
rect 36092 33070 36094 33122
rect 36146 33070 36148 33122
rect 36092 32676 36148 33070
rect 36092 32620 36260 32676
rect 35980 32498 36036 32508
rect 35868 32162 35924 32172
rect 36092 32452 36148 32462
rect 35756 31826 35812 31836
rect 35532 31780 35588 31790
rect 35532 31686 35588 31724
rect 36092 31778 36148 32396
rect 36092 31726 36094 31778
rect 36146 31726 36148 31778
rect 36092 31714 36148 31726
rect 35868 31666 35924 31678
rect 35868 31614 35870 31666
rect 35922 31614 35924 31666
rect 35868 31220 35924 31614
rect 35084 30772 35140 30782
rect 35084 30324 35140 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 30324 35252 30334
rect 35084 30322 35252 30324
rect 35084 30270 35198 30322
rect 35250 30270 35252 30322
rect 35084 30268 35252 30270
rect 35196 30258 35252 30268
rect 35756 30098 35812 30110
rect 35756 30046 35758 30098
rect 35810 30046 35812 30098
rect 35644 29988 35700 29998
rect 34972 29474 35028 29484
rect 35532 29986 35700 29988
rect 35532 29934 35646 29986
rect 35698 29934 35700 29986
rect 35532 29932 35700 29934
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35308 28756 35364 28766
rect 35532 28756 35588 29932
rect 35644 29922 35700 29932
rect 35756 29652 35812 30046
rect 35756 29586 35812 29596
rect 35308 28754 35588 28756
rect 35308 28702 35310 28754
rect 35362 28702 35588 28754
rect 35308 28700 35588 28702
rect 35308 28690 35364 28700
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34860 27188 34916 27198
rect 34860 27074 34916 27132
rect 34860 27022 34862 27074
rect 34914 27022 34916 27074
rect 34860 27010 34916 27022
rect 35308 27186 35364 27198
rect 35308 27134 35310 27186
rect 35362 27134 35364 27186
rect 35308 27076 35364 27134
rect 35308 27010 35364 27020
rect 34412 26852 34804 26908
rect 33740 23762 33796 23772
rect 33964 24050 34020 24062
rect 33964 23998 33966 24050
rect 34018 23998 34020 24050
rect 33964 23940 34020 23998
rect 33964 23604 34020 23884
rect 33516 23548 34020 23604
rect 33516 23154 33572 23548
rect 34076 23492 34132 26852
rect 34188 26178 34244 26190
rect 34188 26126 34190 26178
rect 34242 26126 34244 26178
rect 34188 25732 34244 26126
rect 34188 25666 34244 25676
rect 34188 24612 34244 24622
rect 34188 24276 34244 24556
rect 34300 24500 34356 24510
rect 34636 24500 34692 24510
rect 34300 24498 34692 24500
rect 34300 24446 34302 24498
rect 34354 24446 34638 24498
rect 34690 24446 34692 24498
rect 34300 24444 34692 24446
rect 34300 24434 34356 24444
rect 34636 24434 34692 24444
rect 34188 24220 34468 24276
rect 34412 24050 34468 24220
rect 34412 23998 34414 24050
rect 34466 23998 34468 24050
rect 34412 23986 34468 23998
rect 34636 23940 34692 23950
rect 34636 23846 34692 23884
rect 34076 23426 34132 23436
rect 33516 23102 33518 23154
rect 33570 23102 33572 23154
rect 33516 23090 33572 23102
rect 33628 23380 33684 23390
rect 33628 21812 33684 23324
rect 34188 23380 34244 23390
rect 33740 23268 33796 23278
rect 33740 23174 33796 23212
rect 34188 23154 34244 23324
rect 34188 23102 34190 23154
rect 34242 23102 34244 23154
rect 34188 23090 34244 23102
rect 34636 23156 34692 23166
rect 34636 23062 34692 23100
rect 33852 22260 33908 22270
rect 33852 22166 33908 22204
rect 34524 22260 34580 22270
rect 33740 21812 33796 21822
rect 33628 21810 33796 21812
rect 33628 21758 33742 21810
rect 33794 21758 33796 21810
rect 33628 21756 33796 21758
rect 33180 21476 33236 21486
rect 33180 21474 33460 21476
rect 33180 21422 33182 21474
rect 33234 21422 33460 21474
rect 33180 21420 33460 21422
rect 33180 21410 33236 21420
rect 33068 21362 33124 21374
rect 33068 21310 33070 21362
rect 33122 21310 33124 21362
rect 33068 20916 33124 21310
rect 33068 20850 33124 20860
rect 33404 20242 33460 21420
rect 33404 20190 33406 20242
rect 33458 20190 33460 20242
rect 33404 20178 33460 20190
rect 33628 20916 33684 20926
rect 33068 20132 33124 20142
rect 33068 20018 33124 20076
rect 33068 19966 33070 20018
rect 33122 19966 33124 20018
rect 33068 19954 33124 19966
rect 33292 20018 33348 20030
rect 33292 19966 33294 20018
rect 33346 19966 33348 20018
rect 33292 19908 33348 19966
rect 33516 20020 33572 20030
rect 33516 19926 33572 19964
rect 33628 20018 33684 20860
rect 33628 19966 33630 20018
rect 33682 19966 33684 20018
rect 33628 19954 33684 19966
rect 33740 20244 33796 21756
rect 34524 21586 34580 22204
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34524 21522 34580 21534
rect 34188 20916 34244 20926
rect 34188 20822 34244 20860
rect 34748 20804 34804 26852
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35308 25620 35364 25630
rect 35308 25618 35812 25620
rect 35308 25566 35310 25618
rect 35362 25566 35812 25618
rect 35308 25564 35812 25566
rect 35308 25554 35364 25564
rect 35756 25506 35812 25564
rect 35756 25454 35758 25506
rect 35810 25454 35812 25506
rect 35756 25442 35812 25454
rect 35420 25396 35476 25406
rect 35308 25394 35476 25396
rect 35308 25342 35422 25394
rect 35474 25342 35476 25394
rect 35308 25340 35476 25342
rect 35196 25284 35252 25294
rect 35196 25190 35252 25228
rect 34860 24834 34916 24846
rect 34860 24782 34862 24834
rect 34914 24782 34916 24834
rect 34860 23268 34916 24782
rect 34972 24724 35028 24734
rect 34972 24610 35028 24668
rect 34972 24558 34974 24610
rect 35026 24558 35028 24610
rect 34972 24546 35028 24558
rect 35308 24500 35364 25340
rect 35420 25330 35476 25340
rect 35868 24836 35924 31164
rect 36204 31332 36260 32620
rect 35980 30884 36036 30894
rect 35980 30212 36036 30828
rect 35980 28644 36036 30156
rect 36092 30100 36148 30110
rect 36092 30006 36148 30044
rect 36092 29540 36148 29550
rect 36092 29446 36148 29484
rect 35980 28550 36036 28588
rect 36092 27972 36148 27982
rect 36204 27972 36260 31276
rect 36988 32004 37044 32014
rect 36988 31108 37044 31948
rect 37100 31892 37156 31902
rect 37100 31798 37156 31836
rect 37212 31444 37268 33294
rect 37660 33124 37716 33134
rect 37772 33124 37828 34862
rect 37436 33122 37828 33124
rect 37436 33070 37662 33122
rect 37714 33070 37828 33122
rect 37436 33068 37828 33070
rect 37324 31780 37380 31790
rect 37436 31780 37492 33068
rect 37660 33058 37716 33068
rect 37884 32676 37940 35196
rect 38220 34244 38276 35534
rect 38444 35140 38500 36430
rect 38556 36260 38612 37886
rect 38892 37940 38948 37998
rect 38892 37874 38948 37884
rect 38892 37492 38948 37502
rect 38892 37398 38948 37436
rect 39004 37266 39060 38612
rect 39116 37492 39172 38782
rect 39340 38836 39396 38846
rect 39340 38742 39396 38780
rect 40236 38836 40292 38894
rect 40348 38946 40404 40236
rect 40348 38894 40350 38946
rect 40402 38894 40404 38946
rect 40348 38882 40404 38894
rect 40236 38770 40292 38780
rect 39116 37426 39172 37436
rect 39228 38722 39284 38734
rect 39228 38670 39230 38722
rect 39282 38670 39284 38722
rect 39004 37214 39006 37266
rect 39058 37214 39060 37266
rect 39004 37202 39060 37214
rect 39228 37156 39284 38670
rect 39564 38724 39620 38734
rect 39788 38724 39844 38734
rect 39564 38722 39732 38724
rect 39564 38670 39566 38722
rect 39618 38670 39732 38722
rect 39564 38668 39732 38670
rect 39564 38658 39620 38668
rect 39340 38050 39396 38062
rect 39340 37998 39342 38050
rect 39394 37998 39396 38050
rect 39340 37604 39396 37998
rect 39340 37538 39396 37548
rect 39564 37828 39620 37838
rect 39564 37266 39620 37772
rect 39564 37214 39566 37266
rect 39618 37214 39620 37266
rect 39564 37202 39620 37214
rect 39676 37492 39732 38668
rect 39788 38722 40180 38724
rect 39788 38670 39790 38722
rect 39842 38670 40180 38722
rect 39788 38668 40180 38670
rect 40572 38668 40628 40684
rect 40684 40516 40740 40526
rect 40684 39618 40740 40460
rect 40684 39566 40686 39618
rect 40738 39566 40740 39618
rect 40684 39554 40740 39566
rect 39788 38658 39844 38668
rect 40124 38612 40628 38668
rect 39228 37090 39284 37100
rect 39452 37154 39508 37166
rect 39452 37102 39454 37154
rect 39506 37102 39508 37154
rect 39452 36484 39508 37102
rect 39452 36390 39508 36428
rect 39564 37044 39620 37054
rect 38780 36260 38836 36270
rect 38556 36204 38724 36260
rect 38668 35812 38724 36204
rect 38836 36204 38948 36260
rect 38780 36194 38836 36204
rect 38668 35746 38724 35756
rect 38444 35026 38500 35084
rect 38444 34974 38446 35026
rect 38498 34974 38500 35026
rect 38444 34962 38500 34974
rect 38220 34178 38276 34188
rect 38668 34802 38724 34814
rect 38668 34750 38670 34802
rect 38722 34750 38724 34802
rect 38668 34018 38724 34750
rect 38892 34244 38948 36204
rect 39004 35812 39060 35822
rect 39004 34914 39060 35756
rect 39564 35026 39620 36988
rect 39676 36932 39732 37436
rect 39788 38276 39844 38286
rect 39788 38162 39844 38220
rect 39788 38110 39790 38162
rect 39842 38110 39844 38162
rect 39788 37378 39844 38110
rect 40236 37604 40292 37614
rect 39788 37326 39790 37378
rect 39842 37326 39844 37378
rect 39788 37314 39844 37326
rect 40124 37548 40236 37604
rect 39676 36866 39732 36876
rect 39564 34974 39566 35026
rect 39618 34974 39620 35026
rect 39564 34962 39620 34974
rect 39676 35476 39732 35486
rect 39004 34862 39006 34914
rect 39058 34862 39060 34914
rect 39004 34850 39060 34862
rect 39676 34802 39732 35420
rect 39676 34750 39678 34802
rect 39730 34750 39732 34802
rect 39676 34738 39732 34750
rect 39116 34356 39172 34366
rect 40124 34356 40180 37548
rect 40236 37538 40292 37548
rect 40236 36594 40292 36606
rect 40236 36542 40238 36594
rect 40290 36542 40292 36594
rect 40236 34916 40292 36542
rect 40572 36482 40628 38612
rect 40796 38388 40852 43652
rect 41020 43538 41076 43550
rect 41020 43486 41022 43538
rect 41074 43486 41076 43538
rect 41020 43428 41076 43486
rect 41020 43362 41076 43372
rect 41132 43538 41188 43550
rect 41132 43486 41134 43538
rect 41186 43486 41188 43538
rect 41132 42756 41188 43486
rect 41244 43540 41300 43550
rect 41244 43446 41300 43484
rect 41132 42690 41188 42700
rect 41356 40852 41412 43932
rect 41468 41300 41524 44156
rect 41692 43652 41748 47200
rect 42924 45108 42980 45118
rect 42364 44100 42420 44110
rect 41692 43586 41748 43596
rect 42252 43876 42308 43886
rect 42140 43540 42196 43550
rect 42140 43446 42196 43484
rect 41692 43316 41748 43326
rect 42028 43316 42084 43326
rect 41692 43222 41748 43260
rect 41804 43314 42084 43316
rect 41804 43262 42030 43314
rect 42082 43262 42084 43314
rect 41804 43260 42084 43262
rect 41580 42868 41636 42878
rect 41804 42868 41860 43260
rect 42028 43250 42084 43260
rect 42252 43092 42308 43820
rect 42364 43538 42420 44044
rect 42364 43486 42366 43538
rect 42418 43486 42420 43538
rect 42364 43474 42420 43486
rect 42476 43316 42532 43326
rect 42532 43260 42868 43316
rect 42476 43222 42532 43260
rect 41580 42866 41860 42868
rect 41580 42814 41582 42866
rect 41634 42814 41860 42866
rect 41580 42812 41860 42814
rect 42140 43036 42308 43092
rect 41580 42802 41636 42812
rect 41468 41234 41524 41244
rect 41692 42532 41748 42542
rect 41356 40796 41524 40852
rect 41356 40628 41412 40638
rect 41020 40404 41076 40414
rect 41020 40310 41076 40348
rect 41244 39508 41300 39518
rect 41020 39452 41244 39508
rect 41020 39058 41076 39452
rect 41244 39414 41300 39452
rect 41020 39006 41022 39058
rect 41074 39006 41076 39058
rect 41020 38994 41076 39006
rect 40796 38322 40852 38332
rect 40908 38834 40964 38846
rect 40908 38782 40910 38834
rect 40962 38782 40964 38834
rect 40908 38276 40964 38782
rect 40908 38210 40964 38220
rect 41356 38722 41412 40572
rect 41356 38670 41358 38722
rect 41410 38670 41412 38722
rect 41356 38052 41412 38670
rect 41356 37986 41412 37996
rect 41468 37716 41524 40796
rect 41692 40514 41748 42476
rect 41916 41972 41972 41982
rect 41916 41188 41972 41916
rect 41692 40462 41694 40514
rect 41746 40462 41748 40514
rect 41692 40450 41748 40462
rect 41804 41186 41972 41188
rect 41804 41134 41918 41186
rect 41970 41134 41972 41186
rect 41804 41132 41972 41134
rect 41356 37660 41524 37716
rect 40572 36430 40574 36482
rect 40626 36430 40628 36482
rect 40572 36418 40628 36430
rect 41020 37380 41076 37390
rect 40908 36036 40964 36046
rect 40908 35810 40964 35980
rect 40908 35758 40910 35810
rect 40962 35758 40964 35810
rect 40908 35746 40964 35758
rect 41020 35922 41076 37324
rect 41020 35870 41022 35922
rect 41074 35870 41076 35922
rect 40236 34850 40292 34860
rect 40348 35586 40404 35598
rect 40348 35534 40350 35586
rect 40402 35534 40404 35586
rect 40236 34356 40292 34366
rect 39004 34244 39060 34254
rect 38892 34242 39060 34244
rect 38892 34190 39006 34242
rect 39058 34190 39060 34242
rect 38892 34188 39060 34190
rect 39004 34178 39060 34188
rect 39116 34130 39172 34300
rect 39564 34354 40292 34356
rect 39564 34302 40238 34354
rect 40290 34302 40292 34354
rect 39564 34300 40292 34302
rect 39340 34244 39396 34254
rect 39340 34150 39396 34188
rect 39116 34078 39118 34130
rect 39170 34078 39172 34130
rect 39116 34066 39172 34078
rect 39564 34130 39620 34300
rect 40236 34290 40292 34300
rect 40348 34242 40404 35534
rect 41020 35364 41076 35870
rect 41020 35298 41076 35308
rect 41244 35698 41300 35710
rect 41244 35646 41246 35698
rect 41298 35646 41300 35698
rect 41244 35140 41300 35646
rect 41244 35074 41300 35084
rect 41132 34916 41188 34926
rect 41132 34822 41188 34860
rect 41356 34692 41412 37660
rect 41468 37492 41524 37502
rect 41468 36482 41524 37436
rect 41804 37268 41860 41132
rect 41916 41122 41972 41132
rect 41916 40180 41972 40190
rect 41916 39730 41972 40124
rect 41916 39678 41918 39730
rect 41970 39678 41972 39730
rect 41916 39666 41972 39678
rect 41916 39284 41972 39294
rect 41916 38162 41972 39228
rect 42140 38948 42196 43036
rect 42140 38882 42196 38892
rect 42252 42924 42532 42980
rect 42252 38668 42308 42924
rect 42364 42754 42420 42766
rect 42364 42702 42366 42754
rect 42418 42702 42420 42754
rect 42364 41860 42420 42702
rect 42476 42644 42532 42924
rect 42812 42868 42868 43260
rect 42924 42980 42980 45052
rect 43036 44436 43092 44446
rect 43036 44342 43092 44380
rect 45164 44436 45220 44446
rect 44156 44324 44212 44334
rect 43596 44212 43652 44222
rect 43596 44118 43652 44156
rect 43708 44098 43764 44110
rect 43708 44046 43710 44098
rect 43762 44046 43764 44098
rect 43708 43876 43764 44046
rect 43708 43810 43764 43820
rect 43148 43764 43204 43774
rect 44156 43708 44212 44268
rect 45164 44322 45220 44380
rect 45164 44270 45166 44322
rect 45218 44270 45220 44322
rect 42924 42914 42980 42924
rect 43036 43652 43204 43708
rect 43820 43652 44212 43708
rect 44268 44210 44324 44222
rect 44268 44158 44270 44210
rect 44322 44158 44324 44210
rect 42812 42774 42868 42812
rect 43036 42754 43092 43652
rect 43036 42702 43038 42754
rect 43090 42702 43092 42754
rect 43036 42644 43092 42702
rect 42476 42588 43092 42644
rect 43148 43540 43204 43550
rect 43148 42420 43204 43484
rect 43148 42354 43204 42364
rect 43260 43538 43316 43550
rect 43260 43486 43262 43538
rect 43314 43486 43316 43538
rect 42700 41860 42756 41870
rect 43260 41860 43316 43486
rect 43484 42868 43540 42878
rect 43484 42308 43540 42812
rect 43708 42644 43764 42654
rect 43484 42242 43540 42252
rect 43596 42642 43764 42644
rect 43596 42590 43710 42642
rect 43762 42590 43764 42642
rect 43596 42588 43764 42590
rect 43596 42084 43652 42588
rect 43708 42578 43764 42588
rect 43820 42532 43876 43652
rect 43932 43540 43988 43550
rect 43932 42756 43988 43484
rect 44268 43540 44324 44158
rect 44940 44210 44996 44222
rect 44940 44158 44942 44210
rect 44994 44158 44996 44210
rect 44380 44100 44436 44110
rect 44380 44006 44436 44044
rect 44492 44098 44548 44110
rect 44492 44046 44494 44098
rect 44546 44046 44548 44098
rect 44268 43474 44324 43484
rect 44044 43426 44100 43438
rect 44044 43374 44046 43426
rect 44098 43374 44100 43426
rect 44044 42868 44100 43374
rect 44492 43428 44548 44046
rect 44940 43764 44996 44158
rect 44940 43698 44996 43708
rect 44492 43362 44548 43372
rect 44044 42812 44660 42868
rect 43932 42700 44100 42756
rect 43820 42466 43876 42476
rect 43932 42530 43988 42542
rect 43932 42478 43934 42530
rect 43986 42478 43988 42530
rect 43820 42308 43876 42318
rect 43596 42018 43652 42028
rect 43708 42196 43764 42206
rect 42364 41858 43316 41860
rect 42364 41806 42702 41858
rect 42754 41806 43316 41858
rect 42364 41804 43316 41806
rect 43484 41860 43540 41870
rect 42588 41186 42644 41198
rect 42588 41134 42590 41186
rect 42642 41134 42644 41186
rect 42588 40740 42644 41134
rect 42588 40674 42644 40684
rect 42700 40404 42756 41804
rect 43484 41186 43540 41804
rect 43484 41134 43486 41186
rect 43538 41134 43540 41186
rect 42252 38612 42420 38668
rect 41916 38110 41918 38162
rect 41970 38110 41972 38162
rect 41916 38098 41972 38110
rect 41468 36430 41470 36482
rect 41522 36430 41524 36482
rect 41468 36418 41524 36430
rect 41692 37266 41860 37268
rect 41692 37214 41806 37266
rect 41858 37214 41860 37266
rect 41692 37212 41860 37214
rect 41356 34626 41412 34636
rect 41580 36148 41636 36158
rect 40348 34190 40350 34242
rect 40402 34190 40404 34242
rect 40348 34178 40404 34190
rect 39564 34078 39566 34130
rect 39618 34078 39620 34130
rect 39564 34066 39620 34078
rect 40460 34132 40516 34142
rect 38668 33966 38670 34018
rect 38722 33966 38724 34018
rect 38668 33954 38724 33966
rect 39788 33906 39844 33918
rect 39788 33854 39790 33906
rect 39842 33854 39844 33906
rect 38668 33796 38724 33806
rect 38668 33234 38724 33740
rect 39788 33796 39844 33854
rect 39788 33730 39844 33740
rect 40460 33458 40516 34076
rect 40908 34132 40964 34142
rect 40908 34038 40964 34076
rect 40460 33406 40462 33458
rect 40514 33406 40516 33458
rect 38668 33182 38670 33234
rect 38722 33182 38724 33234
rect 38668 33170 38724 33182
rect 39788 33236 39844 33246
rect 37996 33124 38052 33134
rect 38332 33124 38388 33134
rect 37996 33122 38388 33124
rect 37996 33070 37998 33122
rect 38050 33070 38334 33122
rect 38386 33070 38388 33122
rect 37996 33068 38388 33070
rect 37996 33058 38052 33068
rect 37548 32674 37940 32676
rect 37548 32622 37886 32674
rect 37938 32622 37940 32674
rect 37548 32620 37940 32622
rect 37548 32450 37604 32620
rect 37884 32610 37940 32620
rect 38108 32676 38164 32686
rect 38108 32562 38164 32620
rect 38108 32510 38110 32562
rect 38162 32510 38164 32562
rect 38108 32498 38164 32510
rect 37548 32398 37550 32450
rect 37602 32398 37604 32450
rect 37548 32386 37604 32398
rect 37996 32452 38052 32462
rect 37996 32358 38052 32396
rect 37884 32340 37940 32350
rect 37380 31724 37492 31780
rect 37660 32116 37716 32126
rect 37660 31778 37716 32060
rect 37660 31726 37662 31778
rect 37714 31726 37716 31778
rect 37324 31686 37380 31724
rect 37548 31668 37604 31678
rect 37548 31574 37604 31612
rect 37212 31378 37268 31388
rect 37660 31332 37716 31726
rect 37884 31778 37940 32284
rect 37884 31726 37886 31778
rect 37938 31726 37940 31778
rect 37884 31714 37940 31726
rect 38332 31554 38388 33068
rect 38892 32788 38948 32798
rect 38444 32564 38500 32574
rect 38892 32564 38948 32732
rect 39788 32786 39844 33180
rect 39788 32734 39790 32786
rect 39842 32734 39844 32786
rect 39788 32722 39844 32734
rect 39452 32676 39508 32686
rect 38444 32562 38948 32564
rect 38444 32510 38446 32562
rect 38498 32510 38894 32562
rect 38946 32510 38948 32562
rect 38444 32508 38948 32510
rect 38444 32498 38500 32508
rect 38668 31666 38724 32508
rect 38892 32498 38948 32508
rect 39004 32564 39060 32574
rect 39004 32470 39060 32508
rect 39452 32562 39508 32620
rect 39452 32510 39454 32562
rect 39506 32510 39508 32562
rect 39452 32498 39508 32510
rect 39228 32452 39284 32462
rect 39228 32358 39284 32396
rect 40236 32450 40292 32462
rect 40236 32398 40238 32450
rect 40290 32398 40292 32450
rect 39340 31892 39396 31902
rect 39340 31778 39396 31836
rect 39340 31726 39342 31778
rect 39394 31726 39396 31778
rect 39340 31714 39396 31726
rect 38668 31614 38670 31666
rect 38722 31614 38724 31666
rect 38668 31602 38724 31614
rect 40012 31668 40068 31678
rect 40012 31574 40068 31612
rect 38332 31502 38334 31554
rect 38386 31502 38388 31554
rect 38332 31444 38388 31502
rect 38332 31378 38388 31388
rect 37660 31266 37716 31276
rect 40236 31220 40292 32398
rect 40460 31892 40516 33406
rect 41020 32450 41076 32462
rect 41020 32398 41022 32450
rect 41074 32398 41076 32450
rect 41020 32116 41076 32398
rect 41468 32452 41524 32462
rect 41468 32358 41524 32396
rect 41020 32050 41076 32060
rect 41580 31892 41636 36092
rect 41692 34468 41748 37212
rect 41804 37202 41860 37212
rect 42364 36594 42420 38612
rect 42700 38050 42756 40348
rect 43148 40962 43204 40974
rect 43148 40910 43150 40962
rect 43202 40910 43204 40962
rect 43148 39844 43204 40910
rect 43484 40740 43540 41134
rect 43708 41186 43764 42140
rect 43708 41134 43710 41186
rect 43762 41134 43764 41186
rect 43708 41122 43764 41134
rect 43820 41076 43876 42252
rect 43932 41636 43988 42478
rect 43932 41570 43988 41580
rect 43932 41412 43988 41422
rect 43932 41298 43988 41356
rect 43932 41246 43934 41298
rect 43986 41246 43988 41298
rect 43932 41234 43988 41246
rect 44044 41300 44100 42700
rect 44268 42644 44324 42654
rect 44268 42550 44324 42588
rect 44156 42532 44212 42542
rect 44604 42532 44660 42812
rect 44828 42644 44884 42654
rect 44884 42588 45108 42644
rect 44828 42550 44884 42588
rect 44156 42438 44212 42476
rect 44492 42476 44660 42532
rect 44044 41244 44212 41300
rect 44044 41076 44100 41086
rect 43820 41074 44100 41076
rect 43820 41022 44046 41074
rect 44098 41022 44100 41074
rect 43820 41020 44100 41022
rect 44044 41010 44100 41020
rect 43484 40674 43540 40684
rect 42924 39788 43148 39844
rect 42700 37998 42702 38050
rect 42754 37998 42756 38050
rect 42700 37986 42756 37998
rect 42812 39506 42868 39518
rect 42812 39454 42814 39506
rect 42866 39454 42868 39506
rect 42812 37268 42868 39454
rect 42924 38052 42980 39788
rect 43148 39778 43204 39788
rect 43484 40516 43540 40526
rect 43036 39620 43092 39630
rect 43036 39618 43316 39620
rect 43036 39566 43038 39618
rect 43090 39566 43316 39618
rect 43036 39564 43316 39566
rect 43036 39554 43092 39564
rect 43260 38164 43316 39564
rect 43372 39618 43428 39630
rect 43372 39566 43374 39618
rect 43426 39566 43428 39618
rect 43372 38500 43428 39566
rect 43484 38946 43540 40460
rect 43820 40290 43876 40302
rect 43820 40238 43822 40290
rect 43874 40238 43876 40290
rect 43820 39732 43876 40238
rect 44156 40180 44212 41244
rect 44156 40114 44212 40124
rect 43820 39666 43876 39676
rect 44268 39620 44324 39630
rect 44268 39526 44324 39564
rect 44044 39508 44100 39518
rect 43484 38894 43486 38946
rect 43538 38894 43540 38946
rect 43484 38882 43540 38894
rect 43820 39506 44100 39508
rect 43820 39454 44046 39506
rect 44098 39454 44100 39506
rect 43820 39452 44100 39454
rect 43820 38668 43876 39452
rect 44044 39442 44100 39452
rect 44156 38836 44212 38846
rect 43372 38434 43428 38444
rect 43596 38612 43876 38668
rect 43932 38834 44212 38836
rect 43932 38782 44158 38834
rect 44210 38782 44212 38834
rect 43932 38780 44212 38782
rect 43372 38164 43428 38174
rect 43260 38162 43428 38164
rect 43260 38110 43374 38162
rect 43426 38110 43428 38162
rect 43260 38108 43428 38110
rect 43372 38098 43428 38108
rect 43036 38052 43092 38062
rect 42924 38050 43092 38052
rect 42924 37998 43038 38050
rect 43090 37998 43092 38050
rect 42924 37996 43092 37998
rect 43036 37986 43092 37996
rect 43484 38052 43540 38062
rect 43484 37958 43540 37996
rect 43036 37828 43092 37838
rect 42700 37212 42868 37268
rect 42924 37772 43036 37828
rect 42364 36542 42366 36594
rect 42418 36542 42420 36594
rect 41916 36372 41972 36382
rect 41916 36278 41972 36316
rect 41804 36258 41860 36270
rect 41804 36206 41806 36258
rect 41858 36206 41860 36258
rect 41804 35924 41860 36206
rect 41804 35858 41860 35868
rect 42028 36258 42084 36270
rect 42028 36206 42030 36258
rect 42082 36206 42084 36258
rect 42028 35476 42084 36206
rect 42252 35924 42308 35934
rect 42028 35382 42084 35420
rect 42140 35868 42252 35924
rect 42140 35586 42196 35868
rect 42252 35858 42308 35868
rect 42252 35700 42308 35710
rect 42364 35700 42420 36542
rect 42476 37044 42532 37054
rect 42476 36482 42532 36988
rect 42476 36430 42478 36482
rect 42530 36430 42532 36482
rect 42476 36418 42532 36430
rect 42252 35698 42420 35700
rect 42252 35646 42254 35698
rect 42306 35646 42420 35698
rect 42252 35644 42420 35646
rect 42252 35634 42308 35644
rect 42140 35534 42142 35586
rect 42194 35534 42196 35586
rect 42140 35028 42196 35534
rect 42028 34972 42196 35028
rect 42364 35364 42420 35374
rect 41692 34412 41860 34468
rect 41692 34244 41748 34254
rect 41692 34150 41748 34188
rect 41804 33348 41860 34412
rect 41804 33282 41860 33292
rect 41916 32900 41972 32910
rect 41804 32788 41860 32798
rect 41804 32674 41860 32732
rect 41916 32786 41972 32844
rect 41916 32734 41918 32786
rect 41970 32734 41972 32786
rect 41916 32722 41972 32734
rect 41804 32622 41806 32674
rect 41858 32622 41860 32674
rect 41804 32610 41860 32622
rect 42028 32676 42084 34972
rect 42140 34804 42196 34814
rect 42140 32786 42196 34748
rect 42140 32734 42142 32786
rect 42194 32734 42196 32786
rect 42140 32722 42196 32734
rect 42252 33348 42308 33358
rect 40516 31836 40852 31892
rect 40460 31826 40516 31836
rect 40236 31154 40292 31164
rect 36988 31052 37156 31108
rect 36428 29988 36484 29998
rect 36428 29894 36484 29932
rect 36148 27916 36260 27972
rect 36988 28754 37044 28766
rect 36988 28702 36990 28754
rect 37042 28702 37044 28754
rect 36988 27972 37044 28702
rect 36092 27906 36148 27916
rect 36988 27906 37044 27916
rect 35980 27860 36036 27870
rect 35980 27746 36036 27804
rect 35980 27694 35982 27746
rect 36034 27694 36036 27746
rect 35980 27186 36036 27694
rect 35980 27134 35982 27186
rect 36034 27134 36036 27186
rect 35980 27122 36036 27134
rect 36428 27746 36484 27758
rect 36428 27694 36430 27746
rect 36482 27694 36484 27746
rect 36428 27188 36484 27694
rect 36092 26850 36148 26862
rect 36092 26798 36094 26850
rect 36146 26798 36148 26850
rect 35980 26516 36036 26526
rect 35980 25730 36036 26460
rect 35980 25678 35982 25730
rect 36034 25678 36036 25730
rect 35980 25666 36036 25678
rect 36092 25396 36148 26798
rect 36316 26180 36372 26190
rect 36316 26086 36372 26124
rect 36316 25732 36372 25742
rect 36316 25638 36372 25676
rect 36092 25330 36148 25340
rect 36204 25506 36260 25518
rect 36204 25454 36206 25506
rect 36258 25454 36260 25506
rect 35868 24770 35924 24780
rect 35420 24724 35476 24734
rect 35420 24722 35700 24724
rect 35420 24670 35422 24722
rect 35474 24670 35700 24722
rect 35420 24668 35700 24670
rect 35420 24658 35476 24668
rect 35532 24500 35588 24510
rect 35308 24498 35588 24500
rect 35308 24446 35534 24498
rect 35586 24446 35588 24498
rect 35308 24444 35588 24446
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35308 23940 35364 23950
rect 35196 23938 35364 23940
rect 35196 23886 35310 23938
rect 35362 23886 35364 23938
rect 35196 23884 35364 23886
rect 35532 23940 35588 24444
rect 35644 24164 35700 24668
rect 35756 24498 35812 24510
rect 35756 24446 35758 24498
rect 35810 24446 35812 24498
rect 35756 24276 35812 24446
rect 35868 24500 35924 24510
rect 35868 24406 35924 24444
rect 35868 24276 35924 24286
rect 35756 24220 35868 24276
rect 35868 24210 35924 24220
rect 36204 24276 36260 25454
rect 36204 24210 36260 24220
rect 36316 24836 36372 24846
rect 35644 24108 35812 24164
rect 35756 24052 35812 24108
rect 35756 23996 35924 24052
rect 35644 23940 35700 23950
rect 35532 23938 35700 23940
rect 35532 23886 35646 23938
rect 35698 23886 35700 23938
rect 35532 23884 35700 23886
rect 35196 23828 35252 23884
rect 35308 23874 35364 23884
rect 35644 23874 35700 23884
rect 35196 23762 35252 23772
rect 35868 23492 35924 23996
rect 35644 23436 35924 23492
rect 35980 23996 36260 24052
rect 35644 23378 35700 23436
rect 35644 23326 35646 23378
rect 35698 23326 35700 23378
rect 35644 23314 35700 23326
rect 34972 23268 35028 23278
rect 34860 23212 34972 23268
rect 34972 23202 35028 23212
rect 35868 23268 35924 23278
rect 35420 23156 35476 23166
rect 35756 23156 35812 23166
rect 35420 23154 35588 23156
rect 35420 23102 35422 23154
rect 35474 23102 35588 23154
rect 35420 23100 35588 23102
rect 35420 23090 35476 23100
rect 35084 23042 35140 23054
rect 35084 22990 35086 23042
rect 35138 22990 35140 23042
rect 35084 20914 35140 22990
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22484 35588 23100
rect 35756 22932 35812 23100
rect 35868 23154 35924 23212
rect 35868 23102 35870 23154
rect 35922 23102 35924 23154
rect 35868 23090 35924 23102
rect 35980 22932 36036 23996
rect 36204 23940 36260 23996
rect 36204 23846 36260 23884
rect 35756 22876 36036 22932
rect 36092 23826 36148 23838
rect 36092 23774 36094 23826
rect 36146 23774 36148 23826
rect 36092 23042 36148 23774
rect 36316 23826 36372 24780
rect 36316 23774 36318 23826
rect 36370 23774 36372 23826
rect 36316 23716 36372 23774
rect 36204 23660 36372 23716
rect 36204 23268 36260 23660
rect 36428 23268 36484 27132
rect 37100 27074 37156 31052
rect 39564 30996 39620 31006
rect 38332 30772 38388 30782
rect 37548 30212 37604 30222
rect 37548 30118 37604 30156
rect 38332 30210 38388 30716
rect 38332 30158 38334 30210
rect 38386 30158 38388 30210
rect 38332 30146 38388 30158
rect 37212 29986 37268 29998
rect 37212 29934 37214 29986
rect 37266 29934 37268 29986
rect 37212 29876 37268 29934
rect 37212 27188 37268 29820
rect 38444 28868 38500 28878
rect 38500 28812 38612 28868
rect 38444 28802 38500 28812
rect 38444 28644 38500 28654
rect 37436 28420 37492 28430
rect 37324 27860 37380 27870
rect 37324 27766 37380 27804
rect 37324 27188 37380 27198
rect 37212 27132 37324 27188
rect 37324 27122 37380 27132
rect 37100 27022 37102 27074
rect 37154 27022 37156 27074
rect 37100 27010 37156 27022
rect 37436 26962 37492 28364
rect 38332 27972 38388 27982
rect 38220 27970 38388 27972
rect 38220 27918 38334 27970
rect 38386 27918 38388 27970
rect 38220 27916 38388 27918
rect 37436 26910 37438 26962
rect 37490 26910 37492 26962
rect 37436 26898 37492 26910
rect 37548 27860 37604 27870
rect 37548 26908 37604 27804
rect 37660 27858 37716 27870
rect 37660 27806 37662 27858
rect 37714 27806 37716 27858
rect 37660 27076 37716 27806
rect 37772 27748 37828 27758
rect 38108 27748 38164 27758
rect 37772 27746 38164 27748
rect 37772 27694 37774 27746
rect 37826 27694 38110 27746
rect 38162 27694 38164 27746
rect 37772 27692 38164 27694
rect 37772 27682 37828 27692
rect 38108 27682 38164 27692
rect 37996 27300 38052 27310
rect 37884 27188 37940 27198
rect 37884 27094 37940 27132
rect 37660 27020 37828 27076
rect 37772 26964 37828 27020
rect 37772 26908 37940 26964
rect 37548 26852 37716 26908
rect 37660 26516 37716 26852
rect 37772 26516 37828 26526
rect 37660 26514 37828 26516
rect 37660 26462 37774 26514
rect 37826 26462 37828 26514
rect 37660 26460 37828 26462
rect 37772 26450 37828 26460
rect 37884 26516 37940 26908
rect 37884 26450 37940 26460
rect 36876 26292 36932 26302
rect 37324 26292 37380 26302
rect 37548 26292 37604 26302
rect 36876 26290 37380 26292
rect 36876 26238 36878 26290
rect 36930 26238 37326 26290
rect 37378 26238 37380 26290
rect 36876 26236 37380 26238
rect 36876 26226 36932 26236
rect 36764 26180 36820 26190
rect 36652 26124 36764 26180
rect 36652 25284 36708 26124
rect 36764 26086 36820 26124
rect 37100 25618 37156 26236
rect 37324 26226 37380 26236
rect 37436 26290 37604 26292
rect 37436 26238 37550 26290
rect 37602 26238 37604 26290
rect 37436 26236 37604 26238
rect 37100 25566 37102 25618
rect 37154 25566 37156 25618
rect 37100 25554 37156 25566
rect 37324 25732 37380 25742
rect 37436 25732 37492 26236
rect 37548 26226 37604 26236
rect 37996 26290 38052 27244
rect 38220 26908 38276 27916
rect 38332 27906 38388 27916
rect 38332 27748 38388 27758
rect 38444 27748 38500 28588
rect 38332 27746 38500 27748
rect 38332 27694 38334 27746
rect 38386 27694 38500 27746
rect 38332 27692 38500 27694
rect 38332 27682 38388 27692
rect 38556 27636 38612 28812
rect 39116 28644 39172 28654
rect 39116 28550 39172 28588
rect 39564 28420 39620 30940
rect 39788 30994 39844 31006
rect 39788 30942 39790 30994
rect 39842 30942 39844 30994
rect 39788 30212 39844 30942
rect 40236 30882 40292 30894
rect 40236 30830 40238 30882
rect 40290 30830 40292 30882
rect 40124 30772 40180 30782
rect 40124 30678 40180 30716
rect 39676 29988 39732 29998
rect 39676 29428 39732 29932
rect 39788 29764 39844 30156
rect 40236 29764 40292 30830
rect 40460 30322 40516 30334
rect 40460 30270 40462 30322
rect 40514 30270 40516 30322
rect 39788 29698 39844 29708
rect 40012 29708 40292 29764
rect 40348 30212 40404 30222
rect 39788 29428 39844 29438
rect 39676 29426 39844 29428
rect 39676 29374 39790 29426
rect 39842 29374 39844 29426
rect 39676 29372 39844 29374
rect 39788 28980 39844 29372
rect 39788 28914 39844 28924
rect 39900 29426 39956 29438
rect 39900 29374 39902 29426
rect 39954 29374 39956 29426
rect 39900 28868 39956 29374
rect 40012 29426 40068 29708
rect 40348 29652 40404 30156
rect 40236 29596 40404 29652
rect 40012 29374 40014 29426
rect 40066 29374 40068 29426
rect 40012 29362 40068 29374
rect 40124 29426 40180 29438
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 39900 28802 39956 28812
rect 39900 28644 39956 28654
rect 39900 28550 39956 28588
rect 39564 28354 39620 28364
rect 40124 28420 40180 29374
rect 40124 28354 40180 28364
rect 39564 28084 39620 28094
rect 39116 28082 39620 28084
rect 39116 28030 39566 28082
rect 39618 28030 39620 28082
rect 39116 28028 39620 28030
rect 38892 27972 38948 27982
rect 38892 27878 38948 27916
rect 38780 27860 38836 27870
rect 38780 27766 38836 27804
rect 38444 27580 38612 27636
rect 38444 27186 38500 27580
rect 38444 27134 38446 27186
rect 38498 27134 38500 27186
rect 38444 26908 38500 27134
rect 38780 27300 38836 27310
rect 38780 27186 38836 27244
rect 38892 27300 38948 27310
rect 39116 27300 39172 28028
rect 39564 28018 39620 28028
rect 38892 27298 39172 27300
rect 38892 27246 38894 27298
rect 38946 27246 39172 27298
rect 38892 27244 39172 27246
rect 39228 27860 39284 27870
rect 38892 27234 38948 27244
rect 38780 27134 38782 27186
rect 38834 27134 38836 27186
rect 38780 27122 38836 27134
rect 39228 27074 39284 27804
rect 39452 27860 39508 27870
rect 39452 27858 39620 27860
rect 39452 27806 39454 27858
rect 39506 27806 39620 27858
rect 39452 27804 39620 27806
rect 39452 27794 39508 27804
rect 39228 27022 39230 27074
rect 39282 27022 39284 27074
rect 39228 27010 39284 27022
rect 37996 26238 37998 26290
rect 38050 26238 38052 26290
rect 37996 26226 38052 26238
rect 38108 26852 38276 26908
rect 38332 26852 38500 26908
rect 37660 26180 37716 26190
rect 37660 26086 37716 26124
rect 37324 25730 37492 25732
rect 37324 25678 37326 25730
rect 37378 25678 37492 25730
rect 37324 25676 37492 25678
rect 37324 25508 37380 25676
rect 37324 25442 37380 25452
rect 37548 25508 37604 25518
rect 36652 24722 36708 25228
rect 37436 25396 37492 25406
rect 37100 25172 37156 25182
rect 37100 25060 37156 25116
rect 36876 25004 37156 25060
rect 36764 24836 36820 24846
rect 36764 24742 36820 24780
rect 36652 24670 36654 24722
rect 36706 24670 36708 24722
rect 36652 24658 36708 24670
rect 36204 23202 36260 23212
rect 36316 23212 36484 23268
rect 36540 24276 36596 24286
rect 36092 22990 36094 23042
rect 36146 22990 36148 23042
rect 35532 22428 35812 22484
rect 35644 22260 35700 22270
rect 35308 22148 35364 22158
rect 35308 21698 35364 22092
rect 35308 21646 35310 21698
rect 35362 21646 35364 21698
rect 35308 21634 35364 21646
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35308 21028 35364 21038
rect 35308 20934 35364 20972
rect 35644 21026 35700 22204
rect 35644 20974 35646 21026
rect 35698 20974 35700 21026
rect 35644 20962 35700 20974
rect 35756 21028 35812 22428
rect 35980 22370 36036 22382
rect 35980 22318 35982 22370
rect 36034 22318 36036 22370
rect 35980 22146 36036 22318
rect 35980 22094 35982 22146
rect 36034 22094 36036 22146
rect 35980 22082 36036 22094
rect 35868 21028 35924 21038
rect 35756 21026 35924 21028
rect 35756 20974 35870 21026
rect 35922 20974 35924 21026
rect 35756 20972 35924 20974
rect 35084 20862 35086 20914
rect 35138 20862 35140 20914
rect 35084 20850 35140 20862
rect 34748 20748 34916 20804
rect 34748 20578 34804 20590
rect 34748 20526 34750 20578
rect 34802 20526 34804 20578
rect 34748 20244 34804 20526
rect 33292 19842 33348 19852
rect 33740 19796 33796 20188
rect 34300 20188 34804 20244
rect 34188 20132 34244 20142
rect 34188 20038 34244 20076
rect 33740 19730 33796 19740
rect 34300 20018 34356 20188
rect 34300 19966 34302 20018
rect 34354 19966 34356 20018
rect 33516 19346 33572 19358
rect 33516 19294 33518 19346
rect 33570 19294 33572 19346
rect 33516 19236 33572 19294
rect 33516 19180 34020 19236
rect 32956 19068 33572 19124
rect 33404 18676 33460 18686
rect 33292 18452 33348 18462
rect 32508 18450 32900 18452
rect 32508 18398 32510 18450
rect 32562 18398 32900 18450
rect 32508 18396 32900 18398
rect 32508 18386 32564 18396
rect 31724 17798 31780 17836
rect 31948 18004 32004 18014
rect 31836 17556 31892 17566
rect 31724 16996 31780 17006
rect 31724 16902 31780 16940
rect 31500 14588 31668 14644
rect 31724 16548 31780 16558
rect 31276 14532 31332 14542
rect 31276 13746 31332 14476
rect 31276 13694 31278 13746
rect 31330 13694 31332 13746
rect 31276 13682 31332 13694
rect 31500 13748 31556 14588
rect 31724 14532 31780 16492
rect 31836 16210 31892 17500
rect 31948 17554 32004 17948
rect 31948 17502 31950 17554
rect 32002 17502 32004 17554
rect 31948 17490 32004 17502
rect 32060 17778 32116 17790
rect 32060 17726 32062 17778
rect 32114 17726 32116 17778
rect 31836 16158 31838 16210
rect 31890 16158 31892 16210
rect 31836 16146 31892 16158
rect 31948 16772 32004 16782
rect 31948 15148 32004 16716
rect 32060 16436 32116 17726
rect 32396 17668 32452 17678
rect 32396 17574 32452 17612
rect 32844 17666 32900 18396
rect 32844 17614 32846 17666
rect 32898 17614 32900 17666
rect 32060 16370 32116 16380
rect 32284 16884 32340 16894
rect 32060 16212 32116 16222
rect 32060 16118 32116 16156
rect 32172 15314 32228 15326
rect 32172 15262 32174 15314
rect 32226 15262 32228 15314
rect 32172 15204 32228 15262
rect 31948 15092 32116 15148
rect 32172 15138 32228 15148
rect 31500 13682 31556 13692
rect 31612 14476 31780 14532
rect 31948 14532 32004 14542
rect 31388 13636 31444 13646
rect 31276 11956 31332 11966
rect 31164 11954 31332 11956
rect 31164 11902 31278 11954
rect 31330 11902 31332 11954
rect 31164 11900 31332 11902
rect 31052 11890 31108 11900
rect 31276 11890 31332 11900
rect 31276 11282 31332 11294
rect 31276 11230 31278 11282
rect 31330 11230 31332 11282
rect 31276 10612 31332 11230
rect 31388 10948 31444 13580
rect 31500 12066 31556 12078
rect 31500 12014 31502 12066
rect 31554 12014 31556 12066
rect 31500 11954 31556 12014
rect 31500 11902 31502 11954
rect 31554 11902 31556 11954
rect 31500 11890 31556 11902
rect 31388 10882 31444 10892
rect 31276 10052 31332 10556
rect 31500 10052 31556 10062
rect 31276 9986 31332 9996
rect 31388 9996 31500 10052
rect 30940 9538 30996 9548
rect 31164 9940 31220 9950
rect 30604 9102 30606 9154
rect 30658 9102 30660 9154
rect 30604 9090 30660 9102
rect 31164 9268 31220 9884
rect 30492 9044 30548 9054
rect 29708 8932 29764 8942
rect 29260 8930 29540 8932
rect 29260 8878 29262 8930
rect 29314 8878 29540 8930
rect 29260 8876 29540 8878
rect 29260 8866 29316 8876
rect 29036 8260 29092 8270
rect 29036 8166 29092 8204
rect 29372 8258 29428 8270
rect 29372 8206 29374 8258
rect 29426 8206 29428 8258
rect 29260 8148 29316 8158
rect 29260 8054 29316 8092
rect 29148 6804 29204 6814
rect 29372 6804 29428 8206
rect 29484 7812 29540 8876
rect 29708 8930 29876 8932
rect 29708 8878 29710 8930
rect 29762 8878 29876 8930
rect 29708 8876 29876 8878
rect 29708 8866 29764 8876
rect 29820 8820 29876 8876
rect 29484 7746 29540 7756
rect 29596 8372 29652 8382
rect 29596 8258 29652 8316
rect 29596 8206 29598 8258
rect 29650 8206 29652 8258
rect 29148 6802 29428 6804
rect 29148 6750 29150 6802
rect 29202 6750 29428 6802
rect 29148 6748 29428 6750
rect 29148 6738 29204 6748
rect 29260 6692 29316 6748
rect 29148 5348 29204 5358
rect 29148 5254 29204 5292
rect 29260 5124 29316 6636
rect 29484 5348 29540 5358
rect 29596 5348 29652 8206
rect 29484 5346 29652 5348
rect 29484 5294 29486 5346
rect 29538 5294 29652 5346
rect 29484 5292 29652 5294
rect 29484 5282 29540 5292
rect 29708 5124 29764 5134
rect 29260 5122 29764 5124
rect 29260 5070 29710 5122
rect 29762 5070 29764 5122
rect 29260 5068 29764 5070
rect 29708 5058 29764 5068
rect 28588 4338 28756 4340
rect 28588 4286 28590 4338
rect 28642 4286 28756 4338
rect 28588 4284 28756 4286
rect 28588 4274 28644 4284
rect 28140 4226 28196 4238
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 27468 3780 27524 3790
rect 27244 3778 27524 3780
rect 27244 3726 27470 3778
rect 27522 3726 27524 3778
rect 27244 3724 27524 3726
rect 27468 3714 27524 3724
rect 26684 3668 26740 3678
rect 26684 3554 26740 3612
rect 27580 3668 27636 3678
rect 27580 3574 27636 3612
rect 28140 3668 28196 4174
rect 28140 3602 28196 3612
rect 26684 3502 26686 3554
rect 26738 3502 26740 3554
rect 26684 3490 26740 3502
rect 28700 3554 28756 4284
rect 28812 4274 28868 4284
rect 29484 4900 29540 4910
rect 29260 4228 29316 4238
rect 29260 4134 29316 4172
rect 29484 3666 29540 4844
rect 29820 4564 29876 8764
rect 29932 8372 29988 8382
rect 29988 8316 30100 8372
rect 29932 8306 29988 8316
rect 30044 7364 30100 8316
rect 30492 8260 30548 8988
rect 30492 8258 30884 8260
rect 30492 8206 30494 8258
rect 30546 8206 30884 8258
rect 30492 8204 30884 8206
rect 30492 8194 30548 8204
rect 30156 8034 30212 8046
rect 30156 7982 30158 8034
rect 30210 7982 30212 8034
rect 30156 7924 30212 7982
rect 30156 7858 30212 7868
rect 30828 7698 30884 8204
rect 30828 7646 30830 7698
rect 30882 7646 30884 7698
rect 30828 7634 30884 7646
rect 30940 8258 30996 8270
rect 30940 8206 30942 8258
rect 30994 8206 30996 8258
rect 30156 7364 30212 7374
rect 30044 7362 30212 7364
rect 30044 7310 30158 7362
rect 30210 7310 30212 7362
rect 30044 7308 30212 7310
rect 30156 7298 30212 7308
rect 30268 6804 30324 6814
rect 30044 6580 30100 6590
rect 30044 5346 30100 6524
rect 30044 5294 30046 5346
rect 30098 5294 30100 5346
rect 30044 5282 30100 5294
rect 30268 5124 30324 6748
rect 30940 6692 30996 8206
rect 30380 5348 30436 5358
rect 30380 5254 30436 5292
rect 30380 5124 30436 5134
rect 30268 5122 30436 5124
rect 30268 5070 30382 5122
rect 30434 5070 30436 5122
rect 30268 5068 30436 5070
rect 30380 5058 30436 5068
rect 30940 5124 30996 6636
rect 31164 5906 31220 9212
rect 31388 9156 31444 9996
rect 31500 9986 31556 9996
rect 31388 9042 31444 9100
rect 31612 9044 31668 14476
rect 31948 14418 32004 14476
rect 31948 14366 31950 14418
rect 32002 14366 32004 14418
rect 31948 14354 32004 14366
rect 31724 14306 31780 14318
rect 31724 14254 31726 14306
rect 31778 14254 31780 14306
rect 31724 12516 31780 14254
rect 31836 12852 31892 12862
rect 31836 12758 31892 12796
rect 31724 12450 31780 12460
rect 31388 8990 31390 9042
rect 31442 8990 31444 9042
rect 31388 8978 31444 8990
rect 31500 8988 31668 9044
rect 31724 11954 31780 11966
rect 31724 11902 31726 11954
rect 31778 11902 31780 11954
rect 31500 8930 31556 8988
rect 31500 8878 31502 8930
rect 31554 8878 31556 8930
rect 31500 8820 31556 8878
rect 31724 8932 31780 11902
rect 31948 10948 32004 10958
rect 31948 10834 32004 10892
rect 31948 10782 31950 10834
rect 32002 10782 32004 10834
rect 31948 10770 32004 10782
rect 32060 10834 32116 15092
rect 32284 14530 32340 16828
rect 32620 16884 32676 16894
rect 32284 14478 32286 14530
rect 32338 14478 32340 14530
rect 32284 14466 32340 14478
rect 32396 16548 32452 16558
rect 32172 13972 32228 13982
rect 32172 13878 32228 13916
rect 32396 12852 32452 16492
rect 32620 16098 32676 16828
rect 32620 16046 32622 16098
rect 32674 16046 32676 16098
rect 32620 16034 32676 16046
rect 32732 14532 32788 14542
rect 32732 14438 32788 14476
rect 32508 13636 32564 13646
rect 32508 13542 32564 13580
rect 32844 13188 32900 17614
rect 33292 17666 33348 18396
rect 33404 17778 33460 18620
rect 33516 18452 33572 19068
rect 33964 18564 34020 19180
rect 33852 18452 33908 18462
rect 33516 18450 33908 18452
rect 33516 18398 33518 18450
rect 33570 18398 33854 18450
rect 33906 18398 33908 18450
rect 33516 18396 33908 18398
rect 33516 18386 33572 18396
rect 33852 18386 33908 18396
rect 33740 18228 33796 18238
rect 33404 17726 33406 17778
rect 33458 17726 33460 17778
rect 33404 17714 33460 17726
rect 33628 17892 33684 17902
rect 33292 17614 33294 17666
rect 33346 17614 33348 17666
rect 33292 17602 33348 17614
rect 33516 17442 33572 17454
rect 33516 17390 33518 17442
rect 33570 17390 33572 17442
rect 33068 17108 33124 17118
rect 33516 17108 33572 17390
rect 33068 16994 33124 17052
rect 33068 16942 33070 16994
rect 33122 16942 33124 16994
rect 33068 16930 33124 16942
rect 33404 17052 33572 17108
rect 33404 16548 33460 17052
rect 33404 16482 33460 16492
rect 33516 16884 33572 16894
rect 33180 16436 33236 16446
rect 33180 16100 33236 16380
rect 33180 16006 33236 16044
rect 32956 15874 33012 15886
rect 32956 15822 32958 15874
rect 33010 15822 33012 15874
rect 32956 15148 33012 15822
rect 32956 15092 33460 15148
rect 33180 14756 33236 14766
rect 33180 14642 33236 14700
rect 33180 14590 33182 14642
rect 33234 14590 33236 14642
rect 33180 14578 33236 14590
rect 33292 14420 33348 14430
rect 33180 14196 33236 14206
rect 32844 13122 32900 13132
rect 33068 14140 33180 14196
rect 32620 12964 32676 12974
rect 32620 12870 32676 12908
rect 32396 12796 32564 12852
rect 32508 12740 32564 12796
rect 32508 12684 32676 12740
rect 32396 12628 32452 12638
rect 32284 12572 32396 12628
rect 32172 12068 32228 12078
rect 32172 11974 32228 12012
rect 32060 10782 32062 10834
rect 32114 10782 32116 10834
rect 32060 10164 32116 10782
rect 32284 10834 32340 12572
rect 32396 12562 32452 12572
rect 32508 12180 32564 12190
rect 32396 12124 32508 12180
rect 32396 12066 32452 12124
rect 32508 12114 32564 12124
rect 32396 12014 32398 12066
rect 32450 12014 32452 12066
rect 32396 12002 32452 12014
rect 32508 11954 32564 11966
rect 32508 11902 32510 11954
rect 32562 11902 32564 11954
rect 32508 11172 32564 11902
rect 32508 11106 32564 11116
rect 32620 11844 32676 12684
rect 32284 10782 32286 10834
rect 32338 10782 32340 10834
rect 32284 10770 32340 10782
rect 32508 10836 32564 10846
rect 32508 10724 32564 10780
rect 32396 10722 32564 10724
rect 32396 10670 32510 10722
rect 32562 10670 32564 10722
rect 32396 10668 32564 10670
rect 32172 10500 32228 10510
rect 32172 10406 32228 10444
rect 32396 10164 32452 10668
rect 32508 10658 32564 10668
rect 31724 8866 31780 8876
rect 31948 10108 32116 10164
rect 32172 10108 32452 10164
rect 31276 8764 31556 8820
rect 31612 8820 31668 8830
rect 31276 7474 31332 8764
rect 31612 8370 31668 8764
rect 31612 8318 31614 8370
rect 31666 8318 31668 8370
rect 31612 8306 31668 8318
rect 31836 8818 31892 8830
rect 31836 8766 31838 8818
rect 31890 8766 31892 8818
rect 31836 7700 31892 8766
rect 31948 7700 32004 10108
rect 32060 9940 32116 9950
rect 32172 9940 32228 10108
rect 32060 9938 32228 9940
rect 32060 9886 32062 9938
rect 32114 9886 32228 9938
rect 32060 9884 32228 9886
rect 32508 9940 32564 9950
rect 32060 9874 32116 9884
rect 32508 9846 32564 9884
rect 32396 8930 32452 8942
rect 32396 8878 32398 8930
rect 32450 8878 32452 8930
rect 32284 8820 32340 8830
rect 32284 8726 32340 8764
rect 32060 7700 32116 7710
rect 31948 7698 32116 7700
rect 31948 7646 32062 7698
rect 32114 7646 32116 7698
rect 31948 7644 32116 7646
rect 31836 7634 31892 7644
rect 32060 7634 32116 7644
rect 32172 7700 32228 7710
rect 32396 7700 32452 8878
rect 32620 8372 32676 11788
rect 33068 12178 33124 14140
rect 33180 14130 33236 14140
rect 33292 13970 33348 14364
rect 33292 13918 33294 13970
rect 33346 13918 33348 13970
rect 33292 13906 33348 13918
rect 33292 13748 33348 13758
rect 33180 12740 33236 12750
rect 33180 12404 33236 12684
rect 33180 12338 33236 12348
rect 33068 12126 33070 12178
rect 33122 12126 33124 12178
rect 33068 10948 33124 12126
rect 33180 12180 33236 12190
rect 33180 12066 33236 12124
rect 33292 12180 33348 13692
rect 33404 12628 33460 15092
rect 33516 14418 33572 16828
rect 33628 16100 33684 17836
rect 33740 17666 33796 18172
rect 33740 17614 33742 17666
rect 33794 17614 33796 17666
rect 33740 17602 33796 17614
rect 33964 17666 34020 18508
rect 34300 18340 34356 19966
rect 34524 20020 34580 20030
rect 34524 19926 34580 19964
rect 34748 20018 34804 20030
rect 34748 19966 34750 20018
rect 34802 19966 34804 20018
rect 34412 19908 34468 19918
rect 34412 19814 34468 19852
rect 34524 19796 34580 19806
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 33964 17602 34020 17614
rect 34188 18284 34356 18340
rect 34412 18452 34468 18462
rect 34188 17668 34244 18284
rect 34188 17602 34244 17612
rect 34300 17556 34356 17566
rect 34300 17462 34356 17500
rect 34412 17332 34468 18396
rect 34076 17276 34468 17332
rect 34524 17666 34580 19740
rect 34748 19236 34804 19966
rect 34748 19170 34804 19180
rect 34860 18452 34916 20748
rect 34860 18386 34916 18396
rect 34972 20580 35028 20590
rect 34524 17614 34526 17666
rect 34578 17614 34580 17666
rect 34076 17108 34132 17276
rect 34524 17220 34580 17614
rect 34076 16882 34132 17052
rect 34076 16830 34078 16882
rect 34130 16830 34132 16882
rect 34076 16818 34132 16830
rect 34188 17164 34580 17220
rect 34636 17612 34916 17668
rect 34188 16212 34244 17164
rect 34636 17108 34692 17612
rect 34860 17554 34916 17612
rect 34860 17502 34862 17554
rect 34914 17502 34916 17554
rect 34860 17490 34916 17502
rect 34412 17052 34692 17108
rect 34748 17444 34804 17454
rect 34300 16994 34356 17006
rect 34300 16942 34302 16994
rect 34354 16942 34356 16994
rect 34300 16548 34356 16942
rect 34300 16482 34356 16492
rect 34188 16146 34244 16156
rect 33852 16100 33908 16110
rect 33628 16098 33908 16100
rect 33628 16046 33854 16098
rect 33906 16046 33908 16098
rect 33628 16044 33908 16046
rect 33852 16034 33908 16044
rect 33628 15876 33684 15886
rect 33628 15874 33796 15876
rect 33628 15822 33630 15874
rect 33682 15822 33796 15874
rect 33628 15820 33796 15822
rect 33628 15810 33684 15820
rect 33516 14366 33518 14418
rect 33570 14366 33572 14418
rect 33516 14354 33572 14366
rect 33628 15204 33684 15242
rect 33628 12964 33684 15148
rect 33740 14196 33796 15820
rect 33740 14130 33796 14140
rect 33852 14420 33908 14430
rect 33740 13972 33796 13982
rect 33852 13972 33908 14364
rect 34188 14308 34244 14318
rect 33740 13970 33908 13972
rect 33740 13918 33742 13970
rect 33794 13918 33908 13970
rect 33740 13916 33908 13918
rect 33964 14306 34244 14308
rect 33964 14254 34190 14306
rect 34242 14254 34244 14306
rect 33964 14252 34244 14254
rect 33740 13906 33796 13916
rect 33628 12870 33684 12908
rect 33404 12404 33460 12572
rect 33516 12404 33572 12414
rect 33404 12402 33572 12404
rect 33404 12350 33518 12402
rect 33570 12350 33572 12402
rect 33404 12348 33572 12350
rect 33292 12178 33460 12180
rect 33292 12126 33294 12178
rect 33346 12126 33460 12178
rect 33292 12124 33460 12126
rect 33292 12114 33348 12124
rect 33180 12014 33182 12066
rect 33234 12014 33236 12066
rect 33180 12002 33236 12014
rect 33124 10892 33236 10948
rect 33068 10882 33124 10892
rect 33068 10612 33124 10622
rect 33068 10518 33124 10556
rect 32956 9940 33012 9950
rect 32956 9846 33012 9884
rect 33180 9042 33236 10892
rect 33292 10052 33348 10062
rect 33292 9938 33348 9996
rect 33292 9886 33294 9938
rect 33346 9886 33348 9938
rect 33292 9874 33348 9886
rect 33404 9716 33460 12124
rect 33180 8990 33182 9042
rect 33234 8990 33236 9042
rect 32620 8306 32676 8316
rect 33068 8932 33124 8942
rect 32172 7698 32452 7700
rect 32172 7646 32174 7698
rect 32226 7646 32452 7698
rect 32172 7644 32452 7646
rect 33068 7700 33124 8876
rect 33180 8260 33236 8990
rect 33180 8194 33236 8204
rect 33292 9660 33460 9716
rect 33292 7924 33348 9660
rect 33516 9268 33572 12348
rect 33964 12404 34020 14252
rect 34188 14242 34244 14252
rect 34300 13858 34356 13870
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 34076 13748 34132 13758
rect 34076 13746 34244 13748
rect 34076 13694 34078 13746
rect 34130 13694 34244 13746
rect 34076 13692 34244 13694
rect 34076 13682 34132 13692
rect 34188 12852 34244 13692
rect 34300 13074 34356 13806
rect 34300 13022 34302 13074
rect 34354 13022 34356 13074
rect 34300 13010 34356 13022
rect 34412 12964 34468 17052
rect 34636 16884 34692 16894
rect 34524 15092 34580 15102
rect 34524 14530 34580 15036
rect 34524 14478 34526 14530
rect 34578 14478 34580 14530
rect 34524 14466 34580 14478
rect 34636 13746 34692 16828
rect 34748 15204 34804 17388
rect 34972 17332 35028 20524
rect 35084 19906 35140 19918
rect 35084 19854 35086 19906
rect 35138 19854 35140 19906
rect 35084 18676 35140 19854
rect 35644 19908 35700 19918
rect 35196 19796 35252 19834
rect 35644 19814 35700 19852
rect 35196 19730 35252 19740
rect 35532 19794 35588 19806
rect 35532 19742 35534 19794
rect 35586 19742 35588 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 18610 35140 18620
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 19742
rect 35644 19684 35700 19694
rect 35644 19346 35700 19628
rect 35644 19294 35646 19346
rect 35698 19294 35700 19346
rect 35644 19282 35700 19294
rect 35420 17836 35588 17892
rect 35756 18676 35812 18686
rect 35196 17444 35252 17454
rect 35196 17350 35252 17388
rect 34748 15138 34804 15148
rect 34860 17276 35028 17332
rect 34860 14530 34916 17276
rect 34972 16996 35028 17006
rect 35028 16940 35140 16996
rect 34972 16930 35028 16940
rect 35084 16324 35140 16940
rect 35420 16994 35476 17836
rect 35756 17668 35812 18620
rect 35532 17612 35812 17668
rect 35532 17554 35588 17612
rect 35532 17502 35534 17554
rect 35586 17502 35588 17554
rect 35532 17490 35588 17502
rect 35420 16942 35422 16994
rect 35474 16942 35476 16994
rect 35420 16930 35476 16942
rect 35644 17444 35700 17454
rect 35532 16772 35588 16782
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 16268 35252 16324
rect 35196 16210 35252 16268
rect 35196 16158 35198 16210
rect 35250 16158 35252 16210
rect 35196 16146 35252 16158
rect 34860 14478 34862 14530
rect 34914 14478 34916 14530
rect 34860 14466 34916 14478
rect 35084 16098 35140 16110
rect 35084 16046 35086 16098
rect 35138 16046 35140 16098
rect 35084 15988 35140 16046
rect 34972 14308 35028 14318
rect 34636 13694 34638 13746
rect 34690 13694 34692 13746
rect 34636 13682 34692 13694
rect 34860 14306 35028 14308
rect 34860 14254 34974 14306
rect 35026 14254 35028 14306
rect 34860 14252 35028 14254
rect 34412 12908 34804 12964
rect 34188 12796 34468 12852
rect 33964 12338 34020 12348
rect 34412 12402 34468 12796
rect 34412 12350 34414 12402
rect 34466 12350 34468 12402
rect 34412 12338 34468 12350
rect 33740 12180 33796 12190
rect 33740 12086 33796 12124
rect 34300 12068 34356 12078
rect 33852 11172 33908 11182
rect 33852 10722 33908 11116
rect 33852 10670 33854 10722
rect 33906 10670 33908 10722
rect 33852 10658 33908 10670
rect 34300 9380 34356 12012
rect 34524 11506 34580 11518
rect 34524 11454 34526 11506
rect 34578 11454 34580 11506
rect 34412 11396 34468 11406
rect 34412 9940 34468 11340
rect 34412 9874 34468 9884
rect 34524 9604 34580 11454
rect 34748 10276 34804 12908
rect 34860 12290 34916 14252
rect 34972 14242 35028 14252
rect 35084 14306 35140 15932
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14254 35086 14306
rect 35138 14254 35140 14306
rect 34860 12238 34862 12290
rect 34914 12238 34916 12290
rect 34860 12226 34916 12238
rect 34972 13524 35028 13534
rect 34972 12290 35028 13468
rect 35084 13188 35140 14254
rect 35308 14306 35364 14318
rect 35308 14254 35310 14306
rect 35362 14254 35364 14306
rect 35308 13524 35364 14254
rect 35420 13860 35476 13870
rect 35532 13860 35588 16716
rect 35644 16210 35700 17388
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35644 16146 35700 16158
rect 35420 13858 35588 13860
rect 35420 13806 35422 13858
rect 35474 13806 35588 13858
rect 35420 13804 35588 13806
rect 35644 15428 35700 15438
rect 35756 15428 35812 17612
rect 35700 15372 35812 15428
rect 35420 13794 35476 13804
rect 35644 13636 35700 15372
rect 35868 14756 35924 20972
rect 36092 20356 36148 22990
rect 35980 20300 36148 20356
rect 36204 22146 36260 22158
rect 36204 22094 36206 22146
rect 36258 22094 36260 22146
rect 36204 20914 36260 22094
rect 36204 20862 36206 20914
rect 36258 20862 36260 20914
rect 35980 16996 36036 20300
rect 36092 20132 36148 20142
rect 36092 20038 36148 20076
rect 36204 19460 36260 20862
rect 36204 19394 36260 19404
rect 36316 17892 36372 23212
rect 36428 23042 36484 23054
rect 36428 22990 36430 23042
rect 36482 22990 36484 23042
rect 36428 22930 36484 22990
rect 36428 22878 36430 22930
rect 36482 22878 36484 22930
rect 36428 22866 36484 22878
rect 36428 22146 36484 22158
rect 36428 22094 36430 22146
rect 36482 22094 36484 22146
rect 36428 21026 36484 22094
rect 36540 21700 36596 24220
rect 36876 23380 36932 25004
rect 36988 24834 37044 24846
rect 36988 24782 36990 24834
rect 37042 24782 37044 24834
rect 36988 24052 37044 24782
rect 37100 24722 37156 25004
rect 37100 24670 37102 24722
rect 37154 24670 37156 24722
rect 37100 24658 37156 24670
rect 36988 23996 37268 24052
rect 37212 23940 37268 23996
rect 37436 23940 37492 25340
rect 37548 24946 37604 25452
rect 37548 24894 37550 24946
rect 37602 24894 37604 24946
rect 37548 24882 37604 24894
rect 37660 25282 37716 25294
rect 37660 25230 37662 25282
rect 37714 25230 37716 25282
rect 37660 24722 37716 25230
rect 38108 24948 38164 26852
rect 38108 24882 38164 24892
rect 38220 25620 38276 25630
rect 38220 24946 38276 25564
rect 38332 25508 38388 26852
rect 39564 26850 39620 27804
rect 39788 27858 39844 27870
rect 39788 27806 39790 27858
rect 39842 27806 39844 27858
rect 39564 26798 39566 26850
rect 39618 26798 39620 26850
rect 39564 26628 39620 26798
rect 39564 26562 39620 26572
rect 39676 27746 39732 27758
rect 39676 27694 39678 27746
rect 39730 27694 39732 27746
rect 38444 26516 38500 26526
rect 38444 26422 38500 26460
rect 39452 26404 39508 26414
rect 39676 26404 39732 27694
rect 39788 27748 39844 27806
rect 39788 27682 39844 27692
rect 39900 27858 39956 27870
rect 39900 27806 39902 27858
rect 39954 27806 39956 27858
rect 39900 27298 39956 27806
rect 39900 27246 39902 27298
rect 39954 27246 39956 27298
rect 39900 27234 39956 27246
rect 40012 27076 40068 27086
rect 40012 26982 40068 27020
rect 40236 26628 40292 29596
rect 40348 29428 40404 29438
rect 40460 29428 40516 30270
rect 40796 30210 40852 31836
rect 42028 31892 42084 32620
rect 42140 31892 42196 31902
rect 42028 31890 42196 31892
rect 42028 31838 42142 31890
rect 42194 31838 42196 31890
rect 42028 31836 42196 31838
rect 41580 31826 41636 31836
rect 42140 31826 42196 31836
rect 41804 31780 41860 31790
rect 41020 31220 41076 31230
rect 41804 31220 41860 31724
rect 41020 31218 41524 31220
rect 41020 31166 41022 31218
rect 41074 31166 41524 31218
rect 41020 31164 41524 31166
rect 41020 31154 41076 31164
rect 41356 30994 41412 31006
rect 41356 30942 41358 30994
rect 41410 30942 41412 30994
rect 40796 30158 40798 30210
rect 40850 30158 40852 30210
rect 40796 30146 40852 30158
rect 40908 30882 40964 30894
rect 40908 30830 40910 30882
rect 40962 30830 40964 30882
rect 40348 29426 40516 29428
rect 40348 29374 40350 29426
rect 40402 29374 40516 29426
rect 40348 29372 40516 29374
rect 40348 29362 40404 29372
rect 40348 28868 40404 28878
rect 40348 28642 40404 28812
rect 40348 28590 40350 28642
rect 40402 28590 40404 28642
rect 40348 28578 40404 28590
rect 40460 28420 40516 29372
rect 40796 29652 40852 29662
rect 40796 28532 40852 29596
rect 40908 28754 40964 30830
rect 40908 28702 40910 28754
rect 40962 28702 40964 28754
rect 40908 28690 40964 28702
rect 41020 28980 41076 28990
rect 41020 28642 41076 28924
rect 41020 28590 41022 28642
rect 41074 28590 41076 28642
rect 41020 28578 41076 28590
rect 41356 28754 41412 30942
rect 41468 30324 41524 31164
rect 41804 31126 41860 31164
rect 41580 30996 41636 31006
rect 41580 30902 41636 30940
rect 42028 30994 42084 31006
rect 42028 30942 42030 30994
rect 42082 30942 42084 30994
rect 41692 30882 41748 30894
rect 41692 30830 41694 30882
rect 41746 30830 41748 30882
rect 41580 30324 41636 30334
rect 41468 30322 41636 30324
rect 41468 30270 41582 30322
rect 41634 30270 41636 30322
rect 41468 30268 41636 30270
rect 41580 30258 41636 30268
rect 41356 28702 41358 28754
rect 41410 28702 41412 28754
rect 40796 28530 40964 28532
rect 40796 28478 40798 28530
rect 40850 28478 40964 28530
rect 40796 28476 40964 28478
rect 40796 28466 40852 28476
rect 40348 28364 40516 28420
rect 40572 28420 40628 28430
rect 40348 27188 40404 28364
rect 40572 28196 40628 28364
rect 40572 28140 40852 28196
rect 40796 27524 40852 28140
rect 40796 27458 40852 27468
rect 40460 27300 40516 27310
rect 40460 27298 40852 27300
rect 40460 27246 40462 27298
rect 40514 27246 40852 27298
rect 40460 27244 40852 27246
rect 40460 27234 40516 27244
rect 40348 27122 40404 27132
rect 40796 27074 40852 27244
rect 40796 27022 40798 27074
rect 40850 27022 40852 27074
rect 40796 27010 40852 27022
rect 40348 26964 40404 26974
rect 40348 26962 40516 26964
rect 40348 26910 40350 26962
rect 40402 26910 40516 26962
rect 40348 26908 40516 26910
rect 40348 26898 40404 26908
rect 40460 26852 40516 26908
rect 40572 26852 40628 26862
rect 40460 26796 40572 26852
rect 40572 26786 40628 26796
rect 39900 26572 40292 26628
rect 40348 26740 40404 26750
rect 39900 26514 39956 26572
rect 39900 26462 39902 26514
rect 39954 26462 39956 26514
rect 39900 26450 39956 26462
rect 40348 26514 40404 26684
rect 40348 26462 40350 26514
rect 40402 26462 40404 26514
rect 40348 26450 40404 26462
rect 39452 26402 39844 26404
rect 39452 26350 39454 26402
rect 39506 26350 39844 26402
rect 39452 26348 39844 26350
rect 39452 26338 39508 26348
rect 38780 26290 38836 26302
rect 38780 26238 38782 26290
rect 38834 26238 38836 26290
rect 38556 25620 38612 25630
rect 38332 25452 38500 25508
rect 38332 25284 38388 25294
rect 38444 25284 38500 25452
rect 38556 25506 38612 25564
rect 38556 25454 38558 25506
rect 38610 25454 38612 25506
rect 38556 25442 38612 25454
rect 38780 25508 38836 26238
rect 38780 25442 38836 25452
rect 38892 26180 38948 26190
rect 39788 26180 39844 26348
rect 40236 26180 40292 26190
rect 39788 26124 40068 26180
rect 38892 25508 38948 26124
rect 39340 26068 39396 26078
rect 39228 26066 39396 26068
rect 39228 26014 39342 26066
rect 39394 26014 39396 26066
rect 39228 26012 39396 26014
rect 38892 25506 39060 25508
rect 38892 25454 38894 25506
rect 38946 25454 39060 25506
rect 38892 25452 39060 25454
rect 38892 25442 38948 25452
rect 38780 25284 38836 25294
rect 38444 25228 38612 25284
rect 38332 25190 38388 25228
rect 38220 24894 38222 24946
rect 38274 24894 38276 24946
rect 38220 24882 38276 24894
rect 37660 24670 37662 24722
rect 37714 24670 37716 24722
rect 37660 24164 37716 24670
rect 38108 24724 38164 24734
rect 38108 24630 38164 24668
rect 38332 24722 38388 24734
rect 38332 24670 38334 24722
rect 38386 24670 38388 24722
rect 38332 24388 38388 24670
rect 37660 24098 37716 24108
rect 38108 24332 38388 24388
rect 38108 24052 38164 24332
rect 38332 24164 38388 24174
rect 38108 23996 38276 24052
rect 37548 23940 37604 23950
rect 37884 23940 37940 23950
rect 37212 23938 37380 23940
rect 37212 23886 37214 23938
rect 37266 23886 37380 23938
rect 37212 23884 37380 23886
rect 37436 23938 37940 23940
rect 37436 23886 37550 23938
rect 37602 23886 37886 23938
rect 37938 23886 37940 23938
rect 37436 23884 37940 23886
rect 37212 23874 37268 23884
rect 36988 23828 37044 23838
rect 36988 23734 37044 23772
rect 36540 21634 36596 21644
rect 36764 23378 36932 23380
rect 36764 23326 36878 23378
rect 36930 23326 36932 23378
rect 36764 23324 36932 23326
rect 36428 20974 36430 21026
rect 36482 20974 36484 21026
rect 36428 20962 36484 20974
rect 36652 20020 36708 20030
rect 36652 19906 36708 19964
rect 36652 19854 36654 19906
rect 36706 19854 36708 19906
rect 36428 19236 36484 19246
rect 36428 19234 36596 19236
rect 36428 19182 36430 19234
rect 36482 19182 36596 19234
rect 36428 19180 36596 19182
rect 36428 19170 36484 19180
rect 36316 17836 36484 17892
rect 36316 17668 36372 17678
rect 36204 17666 36372 17668
rect 36204 17614 36318 17666
rect 36370 17614 36372 17666
rect 36204 17612 36372 17614
rect 36092 17554 36148 17566
rect 36092 17502 36094 17554
rect 36146 17502 36148 17554
rect 36092 17220 36148 17502
rect 36092 17154 36148 17164
rect 35980 16930 36036 16940
rect 36092 16100 36148 16110
rect 36092 16006 36148 16044
rect 35868 14690 35924 14700
rect 36092 14642 36148 14654
rect 36092 14590 36094 14642
rect 36146 14590 36148 14642
rect 35868 14532 35924 14542
rect 35868 14438 35924 14476
rect 35644 13570 35700 13580
rect 36092 13524 36148 14590
rect 36204 14532 36260 17612
rect 36316 17602 36372 17612
rect 36428 17220 36484 17836
rect 36204 14438 36260 14476
rect 36316 17164 36484 17220
rect 35308 13468 35588 13524
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13132 35252 13188
rect 34972 12238 34974 12290
rect 35026 12238 35028 12290
rect 34972 12226 35028 12238
rect 35084 12404 35140 12414
rect 35084 12290 35140 12348
rect 35084 12238 35086 12290
rect 35138 12238 35140 12290
rect 35084 12226 35140 12238
rect 35196 12068 35252 13132
rect 35196 12002 35252 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34860 11508 34916 11518
rect 35084 11508 35140 11518
rect 34860 11506 35140 11508
rect 34860 11454 34862 11506
rect 34914 11454 35086 11506
rect 35138 11454 35140 11506
rect 34860 11452 35140 11454
rect 34860 11442 34916 11452
rect 35084 11442 35140 11452
rect 35532 11284 35588 13468
rect 36092 13458 36148 13468
rect 35756 12290 35812 12302
rect 35756 12238 35758 12290
rect 35810 12238 35812 12290
rect 35532 11218 35588 11228
rect 35644 12066 35700 12078
rect 35644 12014 35646 12066
rect 35698 12014 35700 12066
rect 35196 11170 35252 11182
rect 35196 11118 35198 11170
rect 35250 11118 35252 11170
rect 35196 10388 35252 11118
rect 35084 10332 35252 10388
rect 35532 11060 35588 11070
rect 34748 10220 35028 10276
rect 34300 9314 34356 9324
rect 34412 9548 34580 9604
rect 34748 10052 34804 10062
rect 33628 9268 33684 9278
rect 33516 9212 33628 9268
rect 33628 9174 33684 9212
rect 33180 7700 33236 7710
rect 33068 7644 33180 7700
rect 32172 7634 32228 7644
rect 33180 7606 33236 7644
rect 31276 7422 31278 7474
rect 31330 7422 31332 7474
rect 31276 7410 31332 7422
rect 31500 7586 31556 7598
rect 31500 7534 31502 7586
rect 31554 7534 31556 7586
rect 31500 7476 31556 7534
rect 32508 7588 32564 7598
rect 32508 7494 32564 7532
rect 31836 7476 31892 7486
rect 31500 7474 31892 7476
rect 31500 7422 31838 7474
rect 31890 7422 31892 7474
rect 31500 7420 31892 7422
rect 31164 5854 31166 5906
rect 31218 5854 31220 5906
rect 31164 5842 31220 5854
rect 31276 6578 31332 6590
rect 31276 6526 31278 6578
rect 31330 6526 31332 6578
rect 31276 5348 31332 6526
rect 31836 5908 31892 7420
rect 32284 7476 32340 7486
rect 32284 7382 32340 7420
rect 31948 6692 32004 6702
rect 31948 6598 32004 6636
rect 32732 6690 32788 6702
rect 32732 6638 32734 6690
rect 32786 6638 32788 6690
rect 31836 5842 31892 5852
rect 32172 6244 32228 6254
rect 31948 5796 32004 5806
rect 31612 5572 31668 5582
rect 31276 5282 31332 5292
rect 31500 5516 31612 5572
rect 30940 5030 30996 5068
rect 29820 4498 29876 4508
rect 31388 4226 31444 4238
rect 31388 4174 31390 4226
rect 31442 4174 31444 4226
rect 31388 3780 31444 4174
rect 31388 3714 31444 3724
rect 29484 3614 29486 3666
rect 29538 3614 29540 3666
rect 29484 3602 29540 3614
rect 30940 3668 30996 3678
rect 31500 3668 31556 5516
rect 31612 5506 31668 5516
rect 31724 5012 31780 5022
rect 31724 4918 31780 4956
rect 31836 4564 31892 4574
rect 31836 4470 31892 4508
rect 31948 4450 32004 5740
rect 31948 4398 31950 4450
rect 32002 4398 32004 4450
rect 31948 4386 32004 4398
rect 31612 4338 31668 4350
rect 31612 4286 31614 4338
rect 31666 4286 31668 4338
rect 31612 4228 31668 4286
rect 32172 4228 32228 6188
rect 32732 5572 32788 6638
rect 33292 6130 33348 7868
rect 33404 9042 33460 9054
rect 33404 8990 33406 9042
rect 33458 8990 33460 9042
rect 33404 8372 33460 8990
rect 33852 9044 33908 9054
rect 33852 8950 33908 8988
rect 34300 9042 34356 9054
rect 34300 8990 34302 9042
rect 34354 8990 34356 9042
rect 33404 7252 33460 8316
rect 33516 8930 33572 8942
rect 33516 8878 33518 8930
rect 33570 8878 33572 8930
rect 33516 8148 33572 8878
rect 34300 8484 34356 8990
rect 34300 8418 34356 8428
rect 33516 8082 33572 8092
rect 33740 8370 33796 8382
rect 33740 8318 33742 8370
rect 33794 8318 33796 8370
rect 33628 7586 33684 7598
rect 33628 7534 33630 7586
rect 33682 7534 33684 7586
rect 33404 7186 33460 7196
rect 33516 7476 33572 7486
rect 33292 6078 33294 6130
rect 33346 6078 33348 6130
rect 33292 6066 33348 6078
rect 33516 6130 33572 7420
rect 33628 6692 33684 7534
rect 33740 7588 33796 8318
rect 34412 8370 34468 9548
rect 34412 8318 34414 8370
rect 34466 8318 34468 8370
rect 34412 8306 34468 8318
rect 34524 9268 34580 9278
rect 34076 8260 34132 8270
rect 34076 8166 34132 8204
rect 34524 8258 34580 9212
rect 34524 8206 34526 8258
rect 34578 8206 34580 8258
rect 34524 8194 34580 8206
rect 34748 8258 34804 9996
rect 34972 9156 35028 10220
rect 35084 10052 35140 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 9996 35476 10052
rect 35420 9938 35476 9996
rect 35420 9886 35422 9938
rect 35474 9886 35476 9938
rect 35420 9874 35476 9886
rect 35532 9492 35588 11004
rect 35644 10164 35700 12014
rect 35756 10836 35812 12238
rect 35756 10770 35812 10780
rect 35868 12180 35924 12190
rect 35868 11394 35924 12124
rect 35980 12178 36036 12190
rect 35980 12126 35982 12178
rect 36034 12126 36036 12178
rect 35980 12068 36036 12126
rect 35980 12002 36036 12012
rect 36204 11956 36260 11966
rect 35868 11342 35870 11394
rect 35922 11342 35924 11394
rect 35644 10098 35700 10108
rect 35756 10612 35812 10622
rect 35532 9426 35588 9436
rect 35756 9156 35812 10556
rect 35868 10500 35924 11342
rect 35980 11732 36036 11742
rect 35980 11284 36036 11676
rect 36204 11394 36260 11900
rect 36204 11342 36206 11394
rect 36258 11342 36260 11394
rect 36204 11330 36260 11342
rect 35980 11190 36036 11228
rect 36316 10724 36372 17164
rect 36540 16884 36596 19180
rect 36652 18676 36708 19854
rect 36652 18610 36708 18620
rect 36540 16818 36596 16828
rect 36652 17220 36708 17230
rect 36428 15988 36484 15998
rect 36652 15988 36708 17164
rect 36428 15986 36708 15988
rect 36428 15934 36430 15986
rect 36482 15934 36708 15986
rect 36428 15932 36708 15934
rect 36428 15922 36484 15932
rect 36764 15148 36820 23324
rect 36876 23314 36932 23324
rect 37324 23044 37380 23884
rect 37548 23874 37604 23884
rect 37884 23874 37940 23884
rect 37436 23714 37492 23726
rect 37436 23662 37438 23714
rect 37490 23662 37492 23714
rect 37436 23268 37492 23662
rect 37436 23202 37492 23212
rect 37884 23716 37940 23726
rect 37772 23044 37828 23054
rect 37324 22988 37716 23044
rect 37324 22260 37380 22270
rect 37324 22166 37380 22204
rect 36988 22148 37044 22158
rect 36988 22054 37044 22092
rect 37436 21474 37492 22988
rect 37660 22370 37716 22988
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 37660 22306 37716 22318
rect 37436 21422 37438 21474
rect 37490 21422 37492 21474
rect 37436 21410 37492 21422
rect 37772 21810 37828 22988
rect 37884 22260 37940 23660
rect 37996 23714 38052 23726
rect 37996 23662 37998 23714
rect 38050 23662 38052 23714
rect 37996 23156 38052 23662
rect 38108 23716 38164 23726
rect 38108 23622 38164 23660
rect 38220 23380 38276 23996
rect 38332 23826 38388 24108
rect 38332 23774 38334 23826
rect 38386 23774 38388 23826
rect 38332 23762 38388 23774
rect 38444 23716 38500 23726
rect 38332 23380 38388 23390
rect 38220 23324 38332 23380
rect 38332 23314 38388 23324
rect 38220 23156 38276 23166
rect 38444 23156 38500 23660
rect 38556 23380 38612 25228
rect 38780 24612 38836 25228
rect 38892 25282 38948 25294
rect 38892 25230 38894 25282
rect 38946 25230 38948 25282
rect 38892 24836 38948 25230
rect 39004 25284 39060 25452
rect 39228 25506 39284 26012
rect 39340 26002 39396 26012
rect 39676 25508 39732 25518
rect 39228 25454 39230 25506
rect 39282 25454 39284 25506
rect 39228 25442 39284 25454
rect 39564 25506 39732 25508
rect 39564 25454 39678 25506
rect 39730 25454 39732 25506
rect 39564 25452 39732 25454
rect 39004 25218 39060 25228
rect 38892 24780 39396 24836
rect 38780 24546 38836 24556
rect 39004 24612 39060 24622
rect 39004 24518 39060 24556
rect 39228 24500 39284 24510
rect 39116 24498 39284 24500
rect 39116 24446 39230 24498
rect 39282 24446 39284 24498
rect 39116 24444 39284 24446
rect 39116 23828 39172 24444
rect 39228 24434 39284 24444
rect 39340 23940 39396 24780
rect 39452 24724 39508 24734
rect 39452 24630 39508 24668
rect 39564 24050 39620 25452
rect 39676 25442 39732 25452
rect 39564 23998 39566 24050
rect 39618 23998 39620 24050
rect 39564 23986 39620 23998
rect 39676 25284 39732 25294
rect 39900 25284 39956 25294
rect 39452 23940 39508 23950
rect 39340 23938 39508 23940
rect 39340 23886 39454 23938
rect 39506 23886 39508 23938
rect 39340 23884 39508 23886
rect 39452 23874 39508 23884
rect 39676 23938 39732 25228
rect 39676 23886 39678 23938
rect 39730 23886 39732 23938
rect 39676 23874 39732 23886
rect 39788 25282 39956 25284
rect 39788 25230 39902 25282
rect 39954 25230 39956 25282
rect 39788 25228 39956 25230
rect 39116 23772 39396 23828
rect 38556 23324 38724 23380
rect 37996 23154 38276 23156
rect 37996 23102 38222 23154
rect 38274 23102 38276 23154
rect 37996 23100 38276 23102
rect 38220 23090 38276 23100
rect 38332 23100 38500 23156
rect 38556 23156 38612 23166
rect 37996 22932 38052 22942
rect 37996 22484 38052 22876
rect 38108 22932 38164 22942
rect 38332 22932 38388 23100
rect 38556 23062 38612 23100
rect 38108 22930 38388 22932
rect 38108 22878 38110 22930
rect 38162 22878 38388 22930
rect 38108 22876 38388 22878
rect 38444 22930 38500 22942
rect 38668 22932 38724 23324
rect 39116 23268 39172 23278
rect 39116 23174 39172 23212
rect 38444 22878 38446 22930
rect 38498 22878 38500 22930
rect 38108 22866 38164 22876
rect 37996 22428 38164 22484
rect 37996 22260 38052 22270
rect 37884 22258 38052 22260
rect 37884 22206 37998 22258
rect 38050 22206 38052 22258
rect 37884 22204 38052 22206
rect 37996 22194 38052 22204
rect 38108 22036 38164 22428
rect 37772 21758 37774 21810
rect 37826 21758 37828 21810
rect 36988 21028 37044 21038
rect 36988 20690 37044 20972
rect 37324 20804 37380 20814
rect 37772 20804 37828 21758
rect 37996 21980 38164 22036
rect 38444 22036 38500 22878
rect 37324 20802 37828 20804
rect 37324 20750 37326 20802
rect 37378 20750 37774 20802
rect 37826 20750 37828 20802
rect 37324 20748 37828 20750
rect 37324 20738 37380 20748
rect 37772 20738 37828 20748
rect 37884 21252 37940 21262
rect 36988 20638 36990 20690
rect 37042 20638 37044 20690
rect 36988 20626 37044 20638
rect 37100 19908 37156 19918
rect 37100 19814 37156 19852
rect 37548 19906 37604 19918
rect 37548 19854 37550 19906
rect 37602 19854 37604 19906
rect 37548 19684 37604 19854
rect 37884 19906 37940 21196
rect 37996 20692 38052 21980
rect 38444 21970 38500 21980
rect 38556 22876 38724 22932
rect 39004 23154 39060 23166
rect 39004 23102 39006 23154
rect 39058 23102 39060 23154
rect 38556 21812 38612 22876
rect 38892 22148 38948 22158
rect 38892 22054 38948 22092
rect 38220 21756 38612 21812
rect 38892 21812 38948 21822
rect 39004 21812 39060 23102
rect 39228 23156 39284 23166
rect 39340 23156 39396 23772
rect 39452 23156 39508 23166
rect 39340 23154 39508 23156
rect 39340 23102 39454 23154
rect 39506 23102 39508 23154
rect 39340 23100 39508 23102
rect 39228 23062 39284 23100
rect 39452 23090 39508 23100
rect 39788 22708 39844 25228
rect 39900 25218 39956 25228
rect 39900 25060 39956 25070
rect 39900 24834 39956 25004
rect 39900 24782 39902 24834
rect 39954 24782 39956 24834
rect 39900 24770 39956 24782
rect 40012 24834 40068 26124
rect 40236 26086 40292 26124
rect 40236 25620 40292 25630
rect 40012 24782 40014 24834
rect 40066 24782 40068 24834
rect 40012 24770 40068 24782
rect 40124 25394 40180 25406
rect 40124 25342 40126 25394
rect 40178 25342 40180 25394
rect 40124 24836 40180 25342
rect 40124 24770 40180 24780
rect 40236 24722 40292 25564
rect 40796 25620 40852 25630
rect 40796 25526 40852 25564
rect 40236 24670 40238 24722
rect 40290 24670 40292 24722
rect 40236 24658 40292 24670
rect 40348 25394 40404 25406
rect 40908 25396 40964 28476
rect 41244 27970 41300 27982
rect 41244 27918 41246 27970
rect 41298 27918 41300 27970
rect 41020 27858 41076 27870
rect 41020 27806 41022 27858
rect 41074 27806 41076 27858
rect 41020 27748 41076 27806
rect 41244 27860 41300 27918
rect 41244 27794 41300 27804
rect 41020 27682 41076 27692
rect 41020 27076 41076 27086
rect 41020 26982 41076 27020
rect 41244 27076 41300 27086
rect 41244 26982 41300 27020
rect 41356 27074 41412 28702
rect 41692 28756 41748 30830
rect 41916 28980 41972 28990
rect 42028 28980 42084 30942
rect 42252 30212 42308 33292
rect 42364 31780 42420 35308
rect 42700 34802 42756 37212
rect 42812 36482 42868 36494
rect 42812 36430 42814 36482
rect 42866 36430 42868 36482
rect 42812 36370 42868 36430
rect 42812 36318 42814 36370
rect 42866 36318 42868 36370
rect 42812 36306 42868 36318
rect 42924 35698 42980 37772
rect 43036 37762 43092 37772
rect 43260 37826 43316 37838
rect 43260 37774 43262 37826
rect 43314 37774 43316 37826
rect 43260 37492 43316 37774
rect 43260 37426 43316 37436
rect 43372 37156 43428 37166
rect 43596 37156 43652 38612
rect 43036 36258 43092 36270
rect 43036 36206 43038 36258
rect 43090 36206 43092 36258
rect 43036 35924 43092 36206
rect 43036 35858 43092 35868
rect 42924 35646 42926 35698
rect 42978 35646 42980 35698
rect 42924 35634 42980 35646
rect 43372 35698 43428 37100
rect 43484 37100 43652 37156
rect 43708 38050 43764 38062
rect 43708 37998 43710 38050
rect 43762 37998 43764 38050
rect 43484 37044 43540 37100
rect 43484 36596 43540 36988
rect 43708 36820 43764 37998
rect 43932 37156 43988 38780
rect 44156 38770 44212 38780
rect 44044 37938 44100 37950
rect 44044 37886 44046 37938
rect 44098 37886 44100 37938
rect 44044 37604 44100 37886
rect 44156 37940 44212 37950
rect 44156 37846 44212 37884
rect 44380 37828 44436 37838
rect 44380 37734 44436 37772
rect 44044 37538 44100 37548
rect 43932 37090 43988 37100
rect 43708 36754 43764 36764
rect 43596 36596 43652 36606
rect 43484 36594 43652 36596
rect 43484 36542 43598 36594
rect 43650 36542 43652 36594
rect 43484 36540 43652 36542
rect 43596 36530 43652 36540
rect 43932 36482 43988 36494
rect 43932 36430 43934 36482
rect 43986 36430 43988 36482
rect 43820 36372 43876 36382
rect 43372 35646 43374 35698
rect 43426 35646 43428 35698
rect 43372 35634 43428 35646
rect 43708 36370 43876 36372
rect 43708 36318 43822 36370
rect 43874 36318 43876 36370
rect 43708 36316 43876 36318
rect 43148 35140 43204 35150
rect 43148 35046 43204 35084
rect 43708 35140 43764 36316
rect 43820 36306 43876 36316
rect 43932 35140 43988 36430
rect 44492 36036 44548 42476
rect 44940 42420 44996 42430
rect 44604 42308 44660 42318
rect 44604 42084 44660 42252
rect 44604 42018 44660 42028
rect 44716 41972 44772 41982
rect 44716 41878 44772 41916
rect 44828 41188 44884 41198
rect 44828 41094 44884 41132
rect 44940 41186 44996 42364
rect 44940 41134 44942 41186
rect 44994 41134 44996 41186
rect 44716 41076 44772 41086
rect 44604 40628 44660 40638
rect 44604 38668 44660 40572
rect 44716 40402 44772 41020
rect 44940 40964 44996 41134
rect 44716 40350 44718 40402
rect 44770 40350 44772 40402
rect 44716 40338 44772 40350
rect 44828 40908 44996 40964
rect 45052 41188 45108 42588
rect 45164 42196 45220 44270
rect 45612 44100 45668 44110
rect 45612 44006 45668 44044
rect 45948 44098 46004 44110
rect 45948 44046 45950 44098
rect 46002 44046 46004 44098
rect 45948 43652 46004 44046
rect 45948 43586 46004 43596
rect 46172 43426 46228 43438
rect 46172 43374 46174 43426
rect 46226 43374 46228 43426
rect 45276 42868 45332 42878
rect 45276 42754 45332 42812
rect 45276 42702 45278 42754
rect 45330 42702 45332 42754
rect 45276 42690 45332 42702
rect 45388 42642 45444 42654
rect 45388 42590 45390 42642
rect 45442 42590 45444 42642
rect 45388 42196 45444 42590
rect 45220 42140 45444 42196
rect 45500 42642 45556 42654
rect 45500 42590 45502 42642
rect 45554 42590 45556 42642
rect 45500 42196 45556 42590
rect 46060 42642 46116 42654
rect 46060 42590 46062 42642
rect 46114 42590 46116 42642
rect 45164 42130 45220 42140
rect 45500 42130 45556 42140
rect 45948 42530 46004 42542
rect 45948 42478 45950 42530
rect 46002 42478 46004 42530
rect 45388 41636 45444 41646
rect 45164 41412 45220 41422
rect 45164 41318 45220 41356
rect 45276 41188 45332 41198
rect 45052 41186 45332 41188
rect 45052 41134 45278 41186
rect 45330 41134 45332 41186
rect 45052 41132 45332 41134
rect 44828 39618 44884 40908
rect 44828 39566 44830 39618
rect 44882 39566 44884 39618
rect 44828 39554 44884 39566
rect 44940 40740 44996 40750
rect 44940 38946 44996 40684
rect 45052 40402 45108 41132
rect 45276 41122 45332 41132
rect 45052 40350 45054 40402
rect 45106 40350 45108 40402
rect 45052 40338 45108 40350
rect 45164 40404 45220 40414
rect 45164 40310 45220 40348
rect 45388 40402 45444 41580
rect 45836 41300 45892 41310
rect 45836 41206 45892 41244
rect 45948 41188 46004 42478
rect 46060 42532 46116 42590
rect 46172 42644 46228 43374
rect 46172 42588 46564 42644
rect 46116 42476 46452 42532
rect 46060 42438 46116 42476
rect 45948 41122 46004 41132
rect 46284 42308 46340 42318
rect 45612 41076 45668 41086
rect 45388 40350 45390 40402
rect 45442 40350 45444 40402
rect 45388 40338 45444 40350
rect 45500 41020 45612 41076
rect 45052 39620 45108 39630
rect 45052 39060 45108 39564
rect 45164 39396 45220 39406
rect 45164 39302 45220 39340
rect 45052 39058 45332 39060
rect 45052 39006 45054 39058
rect 45106 39006 45332 39058
rect 45052 39004 45332 39006
rect 45052 38994 45108 39004
rect 44940 38894 44942 38946
rect 44994 38894 44996 38946
rect 44940 38882 44996 38894
rect 45164 38836 45220 38846
rect 45164 38742 45220 38780
rect 44604 38612 44884 38668
rect 44716 38500 44772 38510
rect 44716 36148 44772 38444
rect 44828 36596 44884 38612
rect 44940 38164 44996 38174
rect 44940 38070 44996 38108
rect 45052 38052 45108 38062
rect 45052 37958 45108 37996
rect 45276 38050 45332 39004
rect 45500 38836 45556 41020
rect 45612 41010 45668 41020
rect 45724 41074 45780 41086
rect 45724 41022 45726 41074
rect 45778 41022 45780 41074
rect 45612 40628 45668 40638
rect 45612 40534 45668 40572
rect 45724 40404 45780 41022
rect 45948 40964 46004 40974
rect 45948 40870 46004 40908
rect 45836 40740 45892 40750
rect 45836 40514 45892 40684
rect 45836 40462 45838 40514
rect 45890 40462 45892 40514
rect 45836 40450 45892 40462
rect 45724 40338 45780 40348
rect 45948 40402 46004 40414
rect 45948 40350 45950 40402
rect 46002 40350 46004 40402
rect 45612 39618 45668 39630
rect 45612 39566 45614 39618
rect 45666 39566 45668 39618
rect 45612 39060 45668 39566
rect 45948 39396 46004 40350
rect 46172 39396 46228 39406
rect 46004 39340 46116 39396
rect 45948 39330 46004 39340
rect 45612 38994 45668 39004
rect 45948 38948 46004 38958
rect 45724 38946 46004 38948
rect 45724 38894 45950 38946
rect 46002 38894 46004 38946
rect 45724 38892 46004 38894
rect 45612 38836 45668 38846
rect 45500 38834 45668 38836
rect 45500 38782 45614 38834
rect 45666 38782 45668 38834
rect 45500 38780 45668 38782
rect 45612 38770 45668 38780
rect 45724 38668 45780 38892
rect 45948 38882 46004 38892
rect 45500 38612 45780 38668
rect 45276 37998 45278 38050
rect 45330 37998 45332 38050
rect 45276 37986 45332 37998
rect 45388 38050 45444 38062
rect 45388 37998 45390 38050
rect 45442 37998 45444 38050
rect 44940 37826 44996 37838
rect 44940 37774 44942 37826
rect 44994 37774 44996 37826
rect 44940 36820 44996 37774
rect 45388 37044 45444 37998
rect 44940 36754 44996 36764
rect 45164 36988 45444 37044
rect 44828 36540 45108 36596
rect 44828 36372 44884 36382
rect 44828 36278 44884 36316
rect 44940 36260 44996 36270
rect 44940 36148 44996 36204
rect 44716 36092 44996 36148
rect 44492 35980 44996 36036
rect 44044 35588 44100 35598
rect 44044 35586 44772 35588
rect 44044 35534 44046 35586
rect 44098 35534 44772 35586
rect 44044 35532 44772 35534
rect 44044 35522 44100 35532
rect 43708 35074 43764 35084
rect 43820 35084 43988 35140
rect 43820 35028 43876 35084
rect 43708 34914 43764 34926
rect 43708 34862 43710 34914
rect 43762 34862 43764 34914
rect 42700 34750 42702 34802
rect 42754 34750 42756 34802
rect 42700 34738 42756 34750
rect 43372 34802 43428 34814
rect 43372 34750 43374 34802
rect 43426 34750 43428 34802
rect 43372 34692 43428 34750
rect 43372 34626 43428 34636
rect 43484 34802 43540 34814
rect 43484 34750 43486 34802
rect 43538 34750 43540 34802
rect 43484 34244 43540 34750
rect 43708 34356 43764 34862
rect 43708 34290 43764 34300
rect 43484 34178 43540 34188
rect 43820 34018 43876 34972
rect 43820 33966 43822 34018
rect 43874 33966 43876 34018
rect 43820 33954 43876 33966
rect 43932 34914 43988 34926
rect 43932 34862 43934 34914
rect 43986 34862 43988 34914
rect 43932 33796 43988 34862
rect 44716 34580 44772 35532
rect 44940 35138 44996 35980
rect 45052 35364 45108 36540
rect 45164 36482 45220 36988
rect 45500 36596 45556 38612
rect 45948 38388 46004 38398
rect 45948 38162 46004 38332
rect 45948 38110 45950 38162
rect 46002 38110 46004 38162
rect 45948 38098 46004 38110
rect 45836 37938 45892 37950
rect 45836 37886 45838 37938
rect 45890 37886 45892 37938
rect 45836 37716 45892 37886
rect 46060 37938 46116 39340
rect 46172 39302 46228 39340
rect 46060 37886 46062 37938
rect 46114 37886 46116 37938
rect 46060 37874 46116 37886
rect 46284 37716 46340 42252
rect 45836 37660 46340 37716
rect 45500 36594 46116 36596
rect 45500 36542 45502 36594
rect 45554 36542 46116 36594
rect 45500 36540 46116 36542
rect 45500 36530 45556 36540
rect 45164 36430 45166 36482
rect 45218 36430 45220 36482
rect 45164 36418 45220 36430
rect 45276 36260 45332 36270
rect 45052 35308 45220 35364
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44940 35074 44996 35086
rect 44828 34804 44884 34814
rect 44828 34710 44884 34748
rect 45052 34802 45108 34814
rect 45052 34750 45054 34802
rect 45106 34750 45108 34802
rect 45052 34692 45108 34750
rect 44716 34524 44996 34580
rect 44828 34356 44884 34366
rect 44828 34262 44884 34300
rect 44268 34242 44324 34254
rect 44268 34190 44270 34242
rect 44322 34190 44324 34242
rect 43932 33730 43988 33740
rect 44156 34130 44212 34142
rect 44156 34078 44158 34130
rect 44210 34078 44212 34130
rect 42476 33572 42532 33582
rect 42476 32900 42532 33516
rect 42812 33348 42868 33358
rect 42812 33254 42868 33292
rect 42476 32562 42532 32844
rect 44156 32788 44212 34078
rect 44156 32722 44212 32732
rect 42476 32510 42478 32562
rect 42530 32510 42532 32562
rect 42476 32340 42532 32510
rect 43372 32564 43428 32574
rect 43372 32562 43652 32564
rect 43372 32510 43374 32562
rect 43426 32510 43652 32562
rect 43372 32508 43652 32510
rect 43372 32498 43428 32508
rect 42476 32274 42532 32284
rect 42812 32450 42868 32462
rect 42812 32398 42814 32450
rect 42866 32398 42868 32450
rect 42812 32228 42868 32398
rect 42476 31780 42532 31790
rect 42364 31778 42532 31780
rect 42364 31726 42478 31778
rect 42530 31726 42532 31778
rect 42364 31724 42532 31726
rect 42364 31108 42420 31724
rect 42476 31714 42532 31724
rect 42588 31556 42644 31566
rect 42588 31218 42644 31500
rect 42588 31166 42590 31218
rect 42642 31166 42644 31218
rect 42588 31154 42644 31166
rect 42364 31014 42420 31052
rect 42252 29426 42308 30156
rect 42252 29374 42254 29426
rect 42306 29374 42308 29426
rect 42252 29362 42308 29374
rect 42588 30100 42644 30110
rect 41972 28924 42084 28980
rect 42476 28980 42532 28990
rect 41916 28914 41972 28924
rect 41692 28690 41748 28700
rect 42364 28868 42420 28878
rect 42252 28644 42308 28654
rect 42140 27860 42196 27870
rect 42140 27766 42196 27804
rect 41916 27746 41972 27758
rect 41916 27694 41918 27746
rect 41970 27694 41972 27746
rect 41916 27636 41972 27694
rect 41916 27570 41972 27580
rect 41804 27188 41860 27198
rect 41804 27076 41860 27132
rect 41356 27022 41358 27074
rect 41410 27022 41412 27074
rect 41356 26908 41412 27022
rect 41692 27020 41972 27076
rect 41132 26850 41188 26862
rect 41356 26852 41524 26908
rect 41132 26798 41134 26850
rect 41186 26798 41188 26850
rect 41132 25620 41188 26798
rect 41468 26740 41524 26852
rect 41468 26674 41524 26684
rect 41580 26852 41636 26862
rect 41132 25554 41188 25564
rect 41468 26180 41524 26190
rect 40348 25342 40350 25394
rect 40402 25342 40404 25394
rect 40124 24612 40180 24622
rect 40012 24556 40124 24612
rect 40012 23716 40068 24556
rect 40124 24546 40180 24556
rect 40348 24162 40404 25342
rect 40796 25340 40964 25396
rect 41468 25506 41524 26124
rect 41468 25454 41470 25506
rect 41522 25454 41524 25506
rect 40684 25284 40740 25294
rect 40684 25190 40740 25228
rect 40348 24110 40350 24162
rect 40402 24110 40404 24162
rect 40348 24098 40404 24110
rect 40460 24724 40516 24734
rect 40460 24050 40516 24668
rect 40460 23998 40462 24050
rect 40514 23998 40516 24050
rect 40124 23940 40180 23950
rect 40124 23846 40180 23884
rect 40460 23828 40516 23998
rect 40460 23762 40516 23772
rect 40012 23660 40180 23716
rect 39900 22932 39956 22942
rect 39900 22930 40068 22932
rect 39900 22878 39902 22930
rect 39954 22878 40068 22930
rect 39900 22876 40068 22878
rect 39900 22866 39956 22876
rect 39788 22652 39956 22708
rect 39228 22484 39284 22494
rect 39228 22390 39284 22428
rect 39340 22370 39396 22382
rect 39340 22318 39342 22370
rect 39394 22318 39396 22370
rect 38892 21810 39284 21812
rect 38892 21758 38894 21810
rect 38946 21758 39284 21810
rect 38892 21756 39284 21758
rect 38108 21700 38164 21710
rect 38108 20804 38164 21644
rect 38108 20738 38164 20748
rect 37996 20598 38052 20636
rect 38220 20356 38276 21756
rect 38892 21746 38948 21756
rect 38556 21586 38612 21598
rect 38556 21534 38558 21586
rect 38610 21534 38612 21586
rect 38556 21140 38612 21534
rect 39228 21586 39284 21756
rect 39228 21534 39230 21586
rect 39282 21534 39284 21586
rect 39228 21522 39284 21534
rect 38556 21074 38612 21084
rect 39004 21474 39060 21486
rect 39004 21422 39006 21474
rect 39058 21422 39060 21474
rect 39004 20916 39060 21422
rect 39340 21252 39396 22318
rect 39564 22260 39620 22270
rect 39564 22258 39844 22260
rect 39564 22206 39566 22258
rect 39618 22206 39844 22258
rect 39564 22204 39844 22206
rect 39564 22194 39620 22204
rect 39676 21812 39732 21822
rect 39676 21718 39732 21756
rect 39788 21810 39844 22204
rect 39788 21758 39790 21810
rect 39842 21758 39844 21810
rect 39788 21746 39844 21758
rect 39900 21810 39956 22652
rect 40012 22370 40068 22876
rect 40012 22318 40014 22370
rect 40066 22318 40068 22370
rect 40012 22306 40068 22318
rect 39900 21758 39902 21810
rect 39954 21758 39956 21810
rect 39900 21746 39956 21758
rect 39676 21588 39732 21598
rect 39340 21186 39396 21196
rect 39564 21476 39620 21486
rect 38668 20860 39060 20916
rect 39564 20914 39620 21420
rect 39564 20862 39566 20914
rect 39618 20862 39620 20914
rect 38556 20580 38612 20590
rect 37884 19854 37886 19906
rect 37938 19854 37940 19906
rect 37884 19842 37940 19854
rect 37996 20300 38276 20356
rect 38332 20578 38612 20580
rect 38332 20526 38558 20578
rect 38610 20526 38612 20578
rect 38332 20524 38612 20526
rect 37996 19684 38052 20300
rect 38220 20020 38276 20030
rect 38332 20020 38388 20524
rect 38556 20514 38612 20524
rect 38668 20244 38724 20860
rect 39564 20850 39620 20862
rect 39676 20916 39732 21532
rect 40124 20916 40180 23660
rect 40796 23604 40852 25340
rect 41468 25284 41524 25454
rect 41580 25506 41636 26796
rect 41580 25454 41582 25506
rect 41634 25454 41636 25506
rect 41580 25442 41636 25454
rect 41692 26628 41748 27020
rect 41916 26962 41972 27020
rect 41692 25506 41748 26572
rect 41804 26906 41860 26918
rect 41804 26854 41806 26906
rect 41858 26854 41860 26906
rect 41916 26910 41918 26962
rect 41970 26910 41972 26962
rect 41916 26898 41972 26910
rect 41804 26516 41860 26854
rect 42140 26850 42196 26862
rect 42140 26798 42142 26850
rect 42194 26798 42196 26850
rect 42140 26628 42196 26798
rect 42140 26562 42196 26572
rect 41804 26450 41860 26460
rect 42252 26404 42308 28588
rect 42140 26402 42308 26404
rect 42140 26350 42254 26402
rect 42306 26350 42308 26402
rect 42140 26348 42308 26350
rect 41692 25454 41694 25506
rect 41746 25454 41748 25506
rect 41692 25442 41748 25454
rect 42028 25508 42084 25518
rect 42028 25414 42084 25452
rect 41468 25218 41524 25228
rect 40908 25172 40964 25182
rect 40908 24612 40964 25116
rect 41468 25060 41524 25070
rect 41132 24948 41188 24958
rect 41020 24836 41076 24846
rect 41020 24742 41076 24780
rect 41132 24834 41188 24892
rect 41132 24782 41134 24834
rect 41186 24782 41188 24834
rect 40908 24050 40964 24556
rect 40908 23998 40910 24050
rect 40962 23998 40964 24050
rect 40908 23986 40964 23998
rect 41020 24498 41076 24510
rect 41020 24446 41022 24498
rect 41074 24446 41076 24498
rect 41020 23716 41076 24446
rect 41132 23940 41188 24782
rect 41468 24834 41524 25004
rect 41468 24782 41470 24834
rect 41522 24782 41524 24834
rect 41468 24770 41524 24782
rect 41580 24724 41636 24734
rect 41580 24630 41636 24668
rect 41692 24500 41748 24510
rect 41580 24444 41692 24500
rect 41468 24052 41524 24062
rect 41580 24052 41636 24444
rect 41692 24434 41748 24444
rect 42140 24052 42196 26348
rect 42252 26338 42308 26348
rect 42364 25620 42420 28812
rect 42476 27074 42532 28924
rect 42588 27186 42644 30044
rect 42812 29652 42868 32172
rect 43484 32340 43540 32350
rect 42812 29586 42868 29596
rect 42924 31892 42980 31902
rect 42924 27972 42980 31836
rect 43036 31780 43092 31790
rect 43036 31686 43092 31724
rect 43372 31556 43428 31566
rect 43260 31554 43428 31556
rect 43260 31502 43374 31554
rect 43426 31502 43428 31554
rect 43260 31500 43428 31502
rect 43036 30996 43092 31006
rect 43260 30996 43316 31500
rect 43372 31490 43428 31500
rect 43036 30994 43316 30996
rect 43036 30942 43038 30994
rect 43090 30942 43316 30994
rect 43036 30940 43316 30942
rect 43484 30994 43540 32284
rect 43484 30942 43486 30994
rect 43538 30942 43540 30994
rect 43036 30548 43092 30940
rect 43484 30930 43540 30942
rect 43596 30548 43652 32508
rect 44044 32450 44100 32462
rect 44044 32398 44046 32450
rect 44098 32398 44100 32450
rect 43820 31892 43876 31902
rect 43820 31798 43876 31836
rect 43932 31556 43988 31566
rect 43932 31106 43988 31500
rect 43932 31054 43934 31106
rect 43986 31054 43988 31106
rect 43932 31042 43988 31054
rect 43596 30492 43876 30548
rect 43036 30482 43092 30492
rect 43708 30322 43764 30334
rect 43708 30270 43710 30322
rect 43762 30270 43764 30322
rect 43708 30212 43764 30270
rect 43484 30156 43764 30212
rect 43484 28868 43540 30156
rect 43820 29540 43876 30492
rect 44044 30210 44100 32398
rect 44268 30548 44324 34190
rect 44492 34132 44548 34142
rect 44492 34130 44660 34132
rect 44492 34078 44494 34130
rect 44546 34078 44660 34130
rect 44492 34076 44660 34078
rect 44492 34066 44548 34076
rect 44604 33572 44660 34076
rect 44828 33572 44884 33582
rect 44604 33570 44884 33572
rect 44604 33518 44830 33570
rect 44882 33518 44884 33570
rect 44604 33516 44884 33518
rect 44828 33506 44884 33516
rect 44940 33570 44996 34524
rect 44940 33518 44942 33570
rect 44994 33518 44996 33570
rect 44940 33506 44996 33518
rect 44940 33236 44996 33246
rect 44492 32564 44548 32574
rect 44492 31220 44548 32508
rect 44940 31892 44996 33180
rect 44940 31798 44996 31836
rect 45052 33234 45108 34636
rect 45164 34130 45220 35308
rect 45164 34078 45166 34130
rect 45218 34078 45220 34130
rect 45164 33460 45220 34078
rect 45276 34020 45332 36204
rect 45388 36260 45444 36270
rect 45388 36258 45556 36260
rect 45388 36206 45390 36258
rect 45442 36206 45556 36258
rect 45388 36204 45556 36206
rect 45388 36194 45444 36204
rect 45388 36036 45444 36046
rect 45388 34914 45444 35980
rect 45388 34862 45390 34914
rect 45442 34862 45444 34914
rect 45388 34244 45444 34862
rect 45500 34580 45556 36204
rect 45836 36258 45892 36270
rect 45836 36206 45838 36258
rect 45890 36206 45892 36258
rect 45836 35364 45892 36206
rect 46060 35588 46116 36540
rect 46172 36372 46228 36382
rect 46172 36370 46340 36372
rect 46172 36318 46174 36370
rect 46226 36318 46340 36370
rect 46172 36316 46340 36318
rect 46172 36306 46228 36316
rect 46284 35700 46340 36316
rect 46284 35634 46340 35644
rect 46172 35588 46228 35598
rect 46060 35586 46228 35588
rect 46060 35534 46174 35586
rect 46226 35534 46228 35586
rect 46060 35532 46228 35534
rect 46172 35522 46228 35532
rect 45836 35298 45892 35308
rect 45836 35140 45892 35150
rect 45892 35084 46004 35140
rect 45836 35074 45892 35084
rect 45612 34916 45668 34926
rect 45612 34914 45780 34916
rect 45612 34862 45614 34914
rect 45666 34862 45780 34914
rect 45612 34860 45780 34862
rect 45612 34850 45668 34860
rect 45500 34524 45668 34580
rect 45500 34244 45556 34254
rect 45388 34188 45500 34244
rect 45500 34178 45556 34188
rect 45612 34130 45668 34524
rect 45612 34078 45614 34130
rect 45666 34078 45668 34130
rect 45500 34020 45556 34030
rect 45276 34018 45556 34020
rect 45276 33966 45502 34018
rect 45554 33966 45556 34018
rect 45276 33964 45556 33966
rect 45500 33954 45556 33964
rect 45612 33796 45668 34078
rect 45388 33740 45668 33796
rect 45724 33796 45780 34860
rect 45388 33570 45444 33740
rect 45388 33518 45390 33570
rect 45442 33518 45444 33570
rect 45388 33506 45444 33518
rect 45612 33572 45668 33582
rect 45724 33572 45780 33740
rect 45612 33570 45780 33572
rect 45612 33518 45614 33570
rect 45666 33518 45780 33570
rect 45612 33516 45780 33518
rect 45836 34244 45892 34254
rect 45612 33506 45668 33516
rect 45164 33394 45220 33404
rect 45052 33182 45054 33234
rect 45106 33182 45108 33234
rect 44940 31220 44996 31230
rect 44492 31218 44996 31220
rect 44492 31166 44494 31218
rect 44546 31166 44942 31218
rect 44994 31166 44996 31218
rect 44492 31164 44996 31166
rect 44492 31154 44548 31164
rect 44940 31154 44996 31164
rect 44268 30482 44324 30492
rect 44380 31108 44436 31118
rect 44044 30158 44046 30210
rect 44098 30158 44100 30210
rect 44044 30146 44100 30158
rect 44156 30100 44212 30110
rect 44156 30006 44212 30044
rect 43820 29538 44212 29540
rect 43820 29486 43822 29538
rect 43874 29486 44212 29538
rect 43820 29484 44212 29486
rect 43820 29474 43876 29484
rect 43484 28802 43540 28812
rect 43484 28644 43540 28654
rect 43484 28550 43540 28588
rect 44156 28642 44212 29484
rect 44156 28590 44158 28642
rect 44210 28590 44212 28642
rect 43372 28532 43428 28542
rect 42924 27916 43204 27972
rect 42700 27748 42756 27758
rect 42700 27746 43092 27748
rect 42700 27694 42702 27746
rect 42754 27694 43092 27746
rect 42700 27692 43092 27694
rect 42700 27682 42756 27692
rect 42588 27134 42590 27186
rect 42642 27134 42644 27186
rect 42588 27122 42644 27134
rect 42924 27524 42980 27534
rect 42476 27022 42478 27074
rect 42530 27022 42532 27074
rect 42476 27010 42532 27022
rect 42924 27074 42980 27468
rect 42924 27022 42926 27074
rect 42978 27022 42980 27074
rect 42924 27010 42980 27022
rect 42700 26962 42756 26974
rect 42700 26910 42702 26962
rect 42754 26910 42756 26962
rect 42700 26628 42756 26910
rect 42700 25620 42756 26572
rect 43036 25732 43092 27692
rect 43148 27524 43204 27916
rect 43260 27748 43316 27758
rect 43260 27654 43316 27692
rect 43148 27468 43316 27524
rect 43036 25666 43092 25676
rect 43148 27074 43204 27086
rect 43148 27022 43150 27074
rect 43202 27022 43204 27074
rect 43148 26852 43204 27022
rect 42364 25564 42644 25620
rect 42588 25396 42644 25564
rect 42700 25554 42756 25564
rect 43148 25508 43204 26796
rect 43260 26628 43316 27468
rect 43260 26562 43316 26572
rect 43036 25452 43204 25508
rect 43260 25508 43316 25518
rect 42588 25340 42756 25396
rect 42364 25284 42420 25294
rect 42364 25282 42532 25284
rect 42364 25230 42366 25282
rect 42418 25230 42532 25282
rect 42364 25228 42532 25230
rect 42364 25218 42420 25228
rect 42364 24836 42420 24846
rect 41468 24050 41636 24052
rect 41468 23998 41470 24050
rect 41522 23998 41636 24050
rect 41468 23996 41636 23998
rect 42028 23996 42196 24052
rect 42252 24724 42308 24734
rect 41468 23986 41524 23996
rect 41132 23874 41188 23884
rect 41020 23650 41076 23660
rect 41468 23828 41524 23838
rect 40460 23548 40852 23604
rect 40236 23492 40292 23502
rect 40236 23266 40292 23436
rect 40348 23380 40404 23390
rect 40348 23286 40404 23324
rect 40236 23214 40238 23266
rect 40290 23214 40292 23266
rect 40236 23202 40292 23214
rect 40236 21812 40292 21822
rect 40236 21718 40292 21756
rect 40348 21476 40404 21486
rect 40348 21382 40404 21420
rect 40460 21140 40516 23548
rect 41356 23380 41412 23390
rect 41356 23286 41412 23324
rect 41020 23154 41076 23166
rect 41020 23102 41022 23154
rect 41074 23102 41076 23154
rect 41020 22594 41076 23102
rect 41020 22542 41022 22594
rect 41074 22542 41076 22594
rect 41020 22530 41076 22542
rect 41132 23154 41188 23166
rect 41132 23102 41134 23154
rect 41186 23102 41188 23154
rect 40908 22258 40964 22270
rect 40908 22206 40910 22258
rect 40962 22206 40964 22258
rect 40908 21588 40964 22206
rect 41132 21700 41188 23102
rect 41244 23156 41300 23166
rect 41468 23156 41524 23772
rect 41804 23716 41860 23726
rect 41804 23622 41860 23660
rect 41580 23380 41636 23390
rect 41580 23266 41636 23324
rect 41580 23214 41582 23266
rect 41634 23214 41636 23266
rect 41580 23202 41636 23214
rect 41244 23154 41524 23156
rect 41244 23102 41246 23154
rect 41298 23102 41524 23154
rect 41244 23100 41524 23102
rect 42028 23156 42084 23996
rect 42252 23938 42308 24668
rect 42364 24388 42420 24780
rect 42476 24724 42532 25228
rect 42700 24836 42756 25340
rect 42812 25394 42868 25406
rect 42812 25342 42814 25394
rect 42866 25342 42868 25394
rect 42812 25060 42868 25342
rect 42812 24994 42868 25004
rect 42700 24780 42868 24836
rect 42476 24610 42532 24668
rect 42476 24558 42478 24610
rect 42530 24558 42532 24610
rect 42476 24546 42532 24558
rect 42364 24332 42532 24388
rect 42476 24050 42532 24332
rect 42476 23998 42478 24050
rect 42530 23998 42532 24050
rect 42476 23986 42532 23998
rect 42252 23886 42254 23938
rect 42306 23886 42308 23938
rect 42252 23874 42308 23886
rect 42364 23940 42420 23950
rect 42364 23846 42420 23884
rect 42812 23938 42868 24780
rect 42924 24612 42980 24622
rect 42924 24518 42980 24556
rect 43036 24388 43092 25452
rect 43260 25414 43316 25452
rect 43148 25282 43204 25294
rect 43148 25230 43150 25282
rect 43202 25230 43204 25282
rect 43148 24948 43204 25230
rect 43148 24882 43204 24892
rect 43260 25060 43316 25070
rect 42812 23886 42814 23938
rect 42866 23886 42868 23938
rect 42140 23828 42196 23838
rect 42140 23604 42196 23772
rect 42588 23716 42644 23726
rect 42812 23716 42868 23886
rect 42924 24332 43092 24388
rect 43148 24724 43204 24734
rect 42924 23940 42980 24332
rect 42924 23874 42980 23884
rect 43148 23938 43204 24668
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 42588 23622 42644 23660
rect 42700 23660 42868 23716
rect 42140 23548 42420 23604
rect 41244 23090 41300 23100
rect 42028 23090 42084 23100
rect 42252 23380 42308 23390
rect 42252 23266 42308 23324
rect 42252 23214 42254 23266
rect 42306 23214 42308 23266
rect 42252 22372 42308 23214
rect 42364 23266 42420 23548
rect 42700 23492 42756 23660
rect 42700 23426 42756 23436
rect 42364 23214 42366 23266
rect 42418 23214 42420 23266
rect 42364 23202 42420 23214
rect 42476 23268 42532 23278
rect 43148 23268 43204 23886
rect 42476 23266 43204 23268
rect 42476 23214 42478 23266
rect 42530 23214 43204 23266
rect 42476 23212 43204 23214
rect 43260 23828 43316 25004
rect 43372 24722 43428 28476
rect 44156 28532 44212 28590
rect 44156 28466 44212 28476
rect 43932 27300 43988 27310
rect 43820 27244 43932 27300
rect 43820 27186 43876 27244
rect 43932 27234 43988 27244
rect 43820 27134 43822 27186
rect 43874 27134 43876 27186
rect 43820 27122 43876 27134
rect 44044 27076 44100 27086
rect 44044 26982 44100 27020
rect 44380 27076 44436 31052
rect 44940 30212 44996 30222
rect 44940 30118 44996 30156
rect 44940 28756 44996 28766
rect 44940 28662 44996 28700
rect 44828 28644 44884 28654
rect 44828 28550 44884 28588
rect 45052 28532 45108 33182
rect 45388 31892 45444 31902
rect 45388 31798 45444 31836
rect 45724 31780 45780 31790
rect 45388 30882 45444 30894
rect 45388 30830 45390 30882
rect 45442 30830 45444 30882
rect 45388 30212 45444 30830
rect 45444 30156 45556 30212
rect 45388 30118 45444 30156
rect 45388 29652 45444 29662
rect 45388 28754 45444 29596
rect 45388 28702 45390 28754
rect 45442 28702 45444 28754
rect 45388 28690 45444 28702
rect 44940 28476 45108 28532
rect 44828 27860 44884 27870
rect 44716 27300 44772 27310
rect 44716 27206 44772 27244
rect 43372 24670 43374 24722
rect 43426 24670 43428 24722
rect 43372 24658 43428 24670
rect 43484 26850 43540 26862
rect 43484 26798 43486 26850
rect 43538 26798 43540 26850
rect 43372 24164 43428 24174
rect 43484 24164 43540 26798
rect 44268 25506 44324 25518
rect 44268 25454 44270 25506
rect 44322 25454 44324 25506
rect 44156 25282 44212 25294
rect 44156 25230 44158 25282
rect 44210 25230 44212 25282
rect 44044 24612 44100 24622
rect 43372 24162 43540 24164
rect 43372 24110 43374 24162
rect 43426 24110 43540 24162
rect 43372 24108 43540 24110
rect 43708 24610 44100 24612
rect 43708 24558 44046 24610
rect 44098 24558 44100 24610
rect 43708 24556 44100 24558
rect 43708 24162 43764 24556
rect 44044 24546 44100 24556
rect 43708 24110 43710 24162
rect 43762 24110 43764 24162
rect 43372 24098 43428 24108
rect 43708 24098 43764 24110
rect 44156 24164 44212 25230
rect 44268 25284 44324 25454
rect 44268 25218 44324 25228
rect 44156 24098 44212 24108
rect 42476 23202 42532 23212
rect 42252 22306 42308 22316
rect 42364 22932 42420 22942
rect 42364 22594 42420 22876
rect 42364 22542 42366 22594
rect 42418 22542 42420 22594
rect 41804 22260 41860 22270
rect 41804 22166 41860 22204
rect 42140 22146 42196 22158
rect 42140 22094 42142 22146
rect 42194 22094 42196 22146
rect 41132 21644 41412 21700
rect 40908 21522 40964 21532
rect 41244 21364 41300 21374
rect 40460 21074 40516 21084
rect 40572 21362 41300 21364
rect 40572 21310 41246 21362
rect 41298 21310 41300 21362
rect 40572 21308 41300 21310
rect 39676 20802 39732 20860
rect 39676 20750 39678 20802
rect 39730 20750 39732 20802
rect 39676 20738 39732 20750
rect 39788 20860 40180 20916
rect 40348 20916 40404 20926
rect 38780 20692 38836 20702
rect 38780 20598 38836 20636
rect 38892 20580 38948 20590
rect 38892 20578 39060 20580
rect 38892 20526 38894 20578
rect 38946 20526 39060 20578
rect 38892 20524 39060 20526
rect 38892 20514 38948 20524
rect 38892 20244 38948 20254
rect 38668 20242 38948 20244
rect 38668 20190 38894 20242
rect 38946 20190 38948 20242
rect 38668 20188 38948 20190
rect 38892 20178 38948 20188
rect 38444 20132 38500 20142
rect 38556 20132 38612 20142
rect 38444 20130 38556 20132
rect 38444 20078 38446 20130
rect 38498 20078 38556 20130
rect 38444 20076 38556 20078
rect 38612 20076 38724 20132
rect 38444 20066 38500 20076
rect 38556 20038 38612 20076
rect 38276 19964 38388 20020
rect 38220 19954 38276 19964
rect 38220 19796 38276 19806
rect 38220 19794 38388 19796
rect 38220 19742 38222 19794
rect 38274 19742 38388 19794
rect 38220 19740 38388 19742
rect 38220 19730 38276 19740
rect 37548 19628 38052 19684
rect 37772 19460 37828 19470
rect 37548 19236 37604 19246
rect 37212 19122 37268 19134
rect 37212 19070 37214 19122
rect 37266 19070 37268 19122
rect 36876 19012 36932 19022
rect 36876 19010 37044 19012
rect 36876 18958 36878 19010
rect 36930 18958 37044 19010
rect 36876 18956 37044 18958
rect 36876 18946 36932 18956
rect 36988 16772 37044 18956
rect 37100 19010 37156 19022
rect 37100 18958 37102 19010
rect 37154 18958 37156 19010
rect 37100 17444 37156 18958
rect 37212 18676 37268 19070
rect 37212 18610 37268 18620
rect 37100 17378 37156 17388
rect 37212 17556 37268 17566
rect 36988 16706 37044 16716
rect 37212 17108 37268 17500
rect 37212 16210 37268 17052
rect 37212 16158 37214 16210
rect 37266 16158 37268 16210
rect 37212 16146 37268 16158
rect 37436 17554 37492 17566
rect 37436 17502 37438 17554
rect 37490 17502 37492 17554
rect 37436 16884 37492 17502
rect 37436 16098 37492 16828
rect 37548 16770 37604 19180
rect 37548 16718 37550 16770
rect 37602 16718 37604 16770
rect 37548 16706 37604 16718
rect 37436 16046 37438 16098
rect 37490 16046 37492 16098
rect 37436 16034 37492 16046
rect 37772 15314 37828 19404
rect 37884 19010 37940 19022
rect 37884 18958 37886 19010
rect 37938 18958 37940 19010
rect 37884 17892 37940 18958
rect 37996 18452 38052 19628
rect 37996 18386 38052 18396
rect 38220 19010 38276 19022
rect 38220 18958 38222 19010
rect 38274 18958 38276 19010
rect 37884 17826 37940 17836
rect 38220 17668 38276 18958
rect 38332 18900 38388 19740
rect 38668 19346 38724 20076
rect 39004 20130 39060 20524
rect 39340 20578 39396 20590
rect 39340 20526 39342 20578
rect 39394 20526 39396 20578
rect 39004 20078 39006 20130
rect 39058 20078 39060 20130
rect 38668 19294 38670 19346
rect 38722 19294 38724 19346
rect 38668 19282 38724 19294
rect 38780 20020 38836 20030
rect 38780 19348 38836 19964
rect 39004 19908 39060 20078
rect 39116 20132 39172 20142
rect 39116 20038 39172 20076
rect 39340 20132 39396 20526
rect 39340 20066 39396 20076
rect 39452 20578 39508 20590
rect 39452 20526 39454 20578
rect 39506 20526 39508 20578
rect 39452 19908 39508 20526
rect 39788 20188 39844 20860
rect 40348 20822 40404 20860
rect 39900 20690 39956 20702
rect 39900 20638 39902 20690
rect 39954 20638 39956 20690
rect 39900 20580 39956 20638
rect 40236 20580 40292 20590
rect 39900 20578 40292 20580
rect 39900 20526 40238 20578
rect 40290 20526 40292 20578
rect 39900 20524 40292 20526
rect 40236 20514 40292 20524
rect 39788 20132 40180 20188
rect 39564 20020 39620 20030
rect 40012 20020 40068 20030
rect 39564 20018 40068 20020
rect 39564 19966 39566 20018
rect 39618 19966 40014 20018
rect 40066 19966 40068 20018
rect 39564 19964 40068 19966
rect 39564 19954 39620 19964
rect 40012 19954 40068 19964
rect 39004 19852 39508 19908
rect 39900 19794 39956 19806
rect 39900 19742 39902 19794
rect 39954 19742 39956 19794
rect 38780 19282 38836 19292
rect 39116 19348 39172 19358
rect 39004 19236 39060 19246
rect 39004 19142 39060 19180
rect 38332 18834 38388 18844
rect 38668 19010 38724 19022
rect 38668 18958 38670 19010
rect 38722 18958 38724 19010
rect 38668 18676 38724 18958
rect 38444 18452 38500 18462
rect 38220 17612 38388 17668
rect 38332 17108 38388 17612
rect 38332 17014 38388 17052
rect 38444 17106 38500 18396
rect 38668 18004 38724 18620
rect 38780 19010 38836 19022
rect 38780 18958 38782 19010
rect 38834 18958 38836 19010
rect 38780 18228 38836 18958
rect 39116 18676 39172 19292
rect 39676 19348 39732 19358
rect 39676 19254 39732 19292
rect 39564 19236 39620 19246
rect 38892 18620 39172 18676
rect 39228 19122 39284 19134
rect 39228 19070 39230 19122
rect 39282 19070 39284 19122
rect 39228 18676 39284 19070
rect 38892 18562 38948 18620
rect 39228 18610 39284 18620
rect 39340 18900 39396 18910
rect 38892 18510 38894 18562
rect 38946 18510 38948 18562
rect 38892 18498 38948 18510
rect 38780 18162 38836 18172
rect 38668 17948 39060 18004
rect 38444 17054 38446 17106
rect 38498 17054 38500 17106
rect 38444 17042 38500 17054
rect 38668 17220 38724 17230
rect 38668 17106 38724 17164
rect 38668 17054 38670 17106
rect 38722 17054 38724 17106
rect 38668 17042 38724 17054
rect 38220 16996 38276 17006
rect 39004 16996 39060 17948
rect 39340 17106 39396 18844
rect 39564 18562 39620 19180
rect 39788 18676 39844 18686
rect 39788 18582 39844 18620
rect 39564 18510 39566 18562
rect 39618 18510 39620 18562
rect 39564 18498 39620 18510
rect 39900 18338 39956 19742
rect 39900 18286 39902 18338
rect 39954 18286 39956 18338
rect 39900 18274 39956 18286
rect 39340 17054 39342 17106
rect 39394 17054 39396 17106
rect 39340 17042 39396 17054
rect 39452 18228 39508 18238
rect 39452 17106 39508 18172
rect 39452 17054 39454 17106
rect 39506 17054 39508 17106
rect 39452 17042 39508 17054
rect 39228 16996 39284 17006
rect 39004 16994 39284 16996
rect 39004 16942 39230 16994
rect 39282 16942 39284 16994
rect 39004 16940 39284 16942
rect 38220 16210 38276 16940
rect 39228 16930 39284 16940
rect 39900 16996 39956 17006
rect 39900 16902 39956 16940
rect 38556 16884 38612 16894
rect 38556 16790 38612 16828
rect 38892 16882 38948 16894
rect 38892 16830 38894 16882
rect 38946 16830 38948 16882
rect 38892 16324 38948 16830
rect 40012 16884 40068 16894
rect 40012 16790 40068 16828
rect 38220 16158 38222 16210
rect 38274 16158 38276 16210
rect 38220 16146 38276 16158
rect 38780 16268 38892 16324
rect 37772 15262 37774 15314
rect 37826 15262 37828 15314
rect 37772 15148 37828 15262
rect 38668 15428 38724 15438
rect 38668 15314 38724 15372
rect 38668 15262 38670 15314
rect 38722 15262 38724 15314
rect 38668 15250 38724 15262
rect 36764 15092 37268 15148
rect 36764 14756 36820 14766
rect 36428 14306 36484 14318
rect 36428 14254 36430 14306
rect 36482 14254 36484 14306
rect 36428 13076 36484 14254
rect 36428 12982 36484 13020
rect 36652 12292 36708 12330
rect 36652 12226 36708 12236
rect 36428 12180 36484 12190
rect 36428 12086 36484 12124
rect 36652 12068 36708 12078
rect 36540 10948 36596 10958
rect 36428 10836 36484 10846
rect 36428 10742 36484 10780
rect 36540 10834 36596 10892
rect 36540 10782 36542 10834
rect 36594 10782 36596 10834
rect 36316 10658 36372 10668
rect 36540 10612 36596 10782
rect 36652 10722 36708 12012
rect 36764 11620 36820 14700
rect 37212 14530 37268 15092
rect 37212 14478 37214 14530
rect 37266 14478 37268 14530
rect 37212 14420 37268 14478
rect 37212 14354 37268 14364
rect 37436 15092 37828 15148
rect 36988 14308 37044 14318
rect 36988 14214 37044 14252
rect 36876 12962 36932 12974
rect 37212 12964 37268 12974
rect 36876 12910 36878 12962
rect 36930 12910 36932 12962
rect 36876 11956 36932 12910
rect 36876 11890 36932 11900
rect 36988 12962 37268 12964
rect 36988 12910 37214 12962
rect 37266 12910 37268 12962
rect 36988 12908 37268 12910
rect 36764 11564 36932 11620
rect 36652 10670 36654 10722
rect 36706 10670 36708 10722
rect 36652 10658 36708 10670
rect 36876 10724 36932 11564
rect 36988 10948 37044 12908
rect 37212 12898 37268 12908
rect 37212 12738 37268 12750
rect 37212 12686 37214 12738
rect 37266 12686 37268 12738
rect 37212 11732 37268 12686
rect 37324 12178 37380 12190
rect 37324 12126 37326 12178
rect 37378 12126 37380 12178
rect 37324 11844 37380 12126
rect 37324 11778 37380 11788
rect 37212 11666 37268 11676
rect 37436 11620 37492 15092
rect 38332 14642 38388 14654
rect 38332 14590 38334 14642
rect 38386 14590 38388 14642
rect 37548 14532 37604 14542
rect 37548 14418 37604 14476
rect 37996 14532 38052 14542
rect 38332 14532 38388 14590
rect 37996 14530 38388 14532
rect 37996 14478 37998 14530
rect 38050 14478 38388 14530
rect 37996 14476 38388 14478
rect 37996 14466 38052 14476
rect 37548 14366 37550 14418
rect 37602 14366 37604 14418
rect 37548 13634 37604 14366
rect 37548 13582 37550 13634
rect 37602 13582 37604 13634
rect 37548 13570 37604 13582
rect 37884 14418 37940 14430
rect 37884 14366 37886 14418
rect 37938 14366 37940 14418
rect 37884 13076 37940 14366
rect 37996 13634 38052 13646
rect 37996 13582 37998 13634
rect 38050 13582 38052 13634
rect 37996 13524 38052 13582
rect 37996 13458 38052 13468
rect 37884 12964 37940 13020
rect 38332 13074 38388 14476
rect 38332 13022 38334 13074
rect 38386 13022 38388 13074
rect 38332 13010 38388 13022
rect 38444 13746 38500 13758
rect 38444 13694 38446 13746
rect 38498 13694 38500 13746
rect 38444 13186 38500 13694
rect 38444 13134 38446 13186
rect 38498 13134 38500 13186
rect 37996 12964 38052 12974
rect 37884 12962 38052 12964
rect 37884 12910 37998 12962
rect 38050 12910 38052 12962
rect 37884 12908 38052 12910
rect 37996 12898 38052 12908
rect 37548 12850 37604 12862
rect 37548 12798 37550 12850
rect 37602 12798 37604 12850
rect 37548 12292 37604 12798
rect 37548 11620 37604 12236
rect 37884 12738 37940 12750
rect 37884 12686 37886 12738
rect 37938 12686 37940 12738
rect 37660 11844 37716 11854
rect 37884 11844 37940 12686
rect 38444 12180 38500 13134
rect 38780 13076 38836 16268
rect 38892 16258 38948 16268
rect 39788 15540 39844 15550
rect 39788 15446 39844 15484
rect 40124 15204 40180 20132
rect 40236 20018 40292 20030
rect 40236 19966 40238 20018
rect 40290 19966 40292 20018
rect 40236 18900 40292 19966
rect 40572 19460 40628 21308
rect 41244 21298 41300 21308
rect 41020 20916 41076 20926
rect 41356 20916 41412 21644
rect 41804 21474 41860 21486
rect 41804 21422 41806 21474
rect 41858 21422 41860 21474
rect 41580 21364 41636 21374
rect 41580 21270 41636 21308
rect 41020 20914 41300 20916
rect 41020 20862 41022 20914
rect 41074 20862 41300 20914
rect 41020 20860 41300 20862
rect 41020 20850 41076 20860
rect 40908 20804 40964 20814
rect 40684 20690 40740 20702
rect 40684 20638 40686 20690
rect 40738 20638 40740 20690
rect 40684 20188 40740 20638
rect 40908 20690 40964 20748
rect 40908 20638 40910 20690
rect 40962 20638 40964 20690
rect 40908 20626 40964 20638
rect 41244 20188 41300 20860
rect 41356 20822 41412 20860
rect 41804 20692 41860 21422
rect 42140 21474 42196 22094
rect 42252 22148 42308 22158
rect 42252 22054 42308 22092
rect 42364 21586 42420 22542
rect 42812 22484 42868 23212
rect 43260 23044 43316 23772
rect 43036 23042 43316 23044
rect 43036 22990 43262 23042
rect 43314 22990 43316 23042
rect 43036 22988 43316 22990
rect 42924 22932 42980 22942
rect 42924 22838 42980 22876
rect 42812 22428 42980 22484
rect 42700 22372 42756 22382
rect 42756 22316 42868 22372
rect 42700 22278 42756 22316
rect 42812 22036 42868 22316
rect 42924 22148 42980 22428
rect 43036 22370 43092 22988
rect 43260 22978 43316 22988
rect 43372 23940 43428 23950
rect 43148 22484 43204 22494
rect 43148 22390 43204 22428
rect 43036 22318 43038 22370
rect 43090 22318 43092 22370
rect 43036 22306 43092 22318
rect 43260 22258 43316 22270
rect 43260 22206 43262 22258
rect 43314 22206 43316 22258
rect 43260 22148 43316 22206
rect 42924 22092 43316 22148
rect 42812 21980 43316 22036
rect 42364 21534 42366 21586
rect 42418 21534 42420 21586
rect 42364 21522 42420 21534
rect 42140 21422 42142 21474
rect 42194 21422 42196 21474
rect 42140 20916 42196 21422
rect 43260 21474 43316 21980
rect 43260 21422 43262 21474
rect 43314 21422 43316 21474
rect 43260 21410 43316 21422
rect 42700 21364 42756 21374
rect 42700 21270 42756 21308
rect 42140 20850 42196 20860
rect 42476 21140 42532 21150
rect 40684 20132 41076 20188
rect 41244 20132 41748 20188
rect 40908 20018 40964 20030
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40796 19460 40852 19470
rect 40572 19404 40796 19460
rect 40236 18834 40292 18844
rect 40460 19234 40516 19246
rect 40460 19182 40462 19234
rect 40514 19182 40516 19234
rect 40460 18676 40516 19182
rect 40796 19234 40852 19404
rect 40796 19182 40798 19234
rect 40850 19182 40852 19234
rect 40796 19170 40852 19182
rect 40908 19348 40964 19966
rect 40908 18676 40964 19292
rect 41020 19346 41076 20132
rect 41020 19294 41022 19346
rect 41074 19294 41076 19346
rect 41020 19282 41076 19294
rect 41356 19348 41412 19358
rect 41356 19254 41412 19292
rect 40460 18610 40516 18620
rect 40796 18620 40964 18676
rect 40236 18338 40292 18350
rect 40236 18286 40238 18338
rect 40290 18286 40292 18338
rect 40236 16772 40292 18286
rect 40236 16706 40292 16716
rect 40348 18226 40404 18238
rect 40348 18174 40350 18226
rect 40402 18174 40404 18226
rect 40348 16548 40404 18174
rect 40796 17780 40852 18620
rect 40796 17666 40852 17724
rect 40796 17614 40798 17666
rect 40850 17614 40852 17666
rect 40796 17602 40852 17614
rect 40908 18450 40964 18462
rect 40908 18398 40910 18450
rect 40962 18398 40964 18450
rect 40348 16482 40404 16492
rect 40348 16324 40404 16334
rect 40348 16210 40404 16268
rect 40348 16158 40350 16210
rect 40402 16158 40404 16210
rect 40348 16146 40404 16158
rect 40796 16100 40852 16110
rect 40908 16100 40964 18398
rect 41692 18450 41748 20132
rect 41804 19348 41860 20636
rect 41804 19282 41860 19292
rect 41692 18398 41694 18450
rect 41746 18398 41748 18450
rect 41692 18386 41748 18398
rect 41356 17668 41412 17678
rect 41132 17108 41188 17118
rect 41132 16882 41188 17052
rect 41356 17106 41412 17612
rect 41356 17054 41358 17106
rect 41410 17054 41412 17106
rect 41356 17042 41412 17054
rect 41580 17220 41636 17230
rect 41580 17106 41636 17164
rect 41580 17054 41582 17106
rect 41634 17054 41636 17106
rect 41580 17042 41636 17054
rect 42252 17108 42308 17118
rect 41132 16830 41134 16882
rect 41186 16830 41188 16882
rect 41132 16818 41188 16830
rect 41804 16882 41860 16894
rect 41804 16830 41806 16882
rect 41858 16830 41860 16882
rect 41468 16772 41524 16782
rect 41468 16678 41524 16716
rect 41468 16548 41524 16558
rect 41468 16210 41524 16492
rect 41468 16158 41470 16210
rect 41522 16158 41524 16210
rect 41468 16146 41524 16158
rect 41804 16100 41860 16830
rect 42252 16882 42308 17052
rect 42476 17106 42532 21084
rect 43372 19908 43428 23884
rect 43596 23938 43652 23950
rect 43596 23886 43598 23938
rect 43650 23886 43652 23938
rect 43596 20804 43652 23886
rect 44156 23826 44212 23838
rect 44156 23774 44158 23826
rect 44210 23774 44212 23826
rect 44044 23716 44100 23726
rect 44044 23622 44100 23660
rect 44156 23380 44212 23774
rect 44380 23604 44436 27020
rect 44828 26962 44884 27804
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44828 26898 44884 26910
rect 44828 25732 44884 25742
rect 44828 25638 44884 25676
rect 44940 25172 44996 28476
rect 45388 27748 45444 27758
rect 45164 27746 45444 27748
rect 45164 27694 45390 27746
rect 45442 27694 45444 27746
rect 45164 27692 45444 27694
rect 45052 27188 45108 27198
rect 45052 27074 45108 27132
rect 45052 27022 45054 27074
rect 45106 27022 45108 27074
rect 45052 27010 45108 27022
rect 45164 25730 45220 27692
rect 45388 27682 45444 27692
rect 45276 26962 45332 26974
rect 45276 26910 45278 26962
rect 45330 26910 45332 26962
rect 45276 26516 45332 26910
rect 45276 26450 45332 26460
rect 45500 26290 45556 30156
rect 45724 28644 45780 31724
rect 45836 31218 45892 34188
rect 45948 33572 46004 35084
rect 46172 35028 46228 35038
rect 46172 34934 46228 34972
rect 46396 34804 46452 42476
rect 46172 34748 46452 34804
rect 46508 38836 46564 42588
rect 46060 34690 46116 34702
rect 46060 34638 46062 34690
rect 46114 34638 46116 34690
rect 46060 34356 46116 34638
rect 46060 34290 46116 34300
rect 46172 34242 46228 34748
rect 46172 34190 46174 34242
rect 46226 34190 46228 34242
rect 46172 34178 46228 34190
rect 46060 33572 46116 33582
rect 45948 33570 46116 33572
rect 45948 33518 46062 33570
rect 46114 33518 46116 33570
rect 45948 33516 46116 33518
rect 46060 33506 46116 33516
rect 46172 33460 46228 33470
rect 46172 33366 46228 33404
rect 46508 32676 46564 38780
rect 46844 40180 46900 40190
rect 46844 39396 46900 40124
rect 46060 32620 46564 32676
rect 46620 35700 46676 35710
rect 45948 31556 46004 31566
rect 45948 31462 46004 31500
rect 45836 31166 45838 31218
rect 45890 31166 45892 31218
rect 45836 31154 45892 31166
rect 45948 31108 46004 31118
rect 46060 31108 46116 32620
rect 46172 32452 46228 32462
rect 46172 32450 46340 32452
rect 46172 32398 46174 32450
rect 46226 32398 46340 32450
rect 46172 32396 46340 32398
rect 46172 32386 46228 32396
rect 45948 31106 46116 31108
rect 45948 31054 45950 31106
rect 46002 31054 46116 31106
rect 45948 31052 46116 31054
rect 45948 31042 46004 31052
rect 46172 30996 46228 31006
rect 45836 30548 45892 30558
rect 45836 30098 45892 30492
rect 46172 30212 46228 30940
rect 45836 30046 45838 30098
rect 45890 30046 45892 30098
rect 45836 30034 45892 30046
rect 45948 30210 46228 30212
rect 45948 30158 46174 30210
rect 46226 30158 46228 30210
rect 45948 30156 46228 30158
rect 45836 28644 45892 28654
rect 45724 28642 45892 28644
rect 45724 28590 45838 28642
rect 45890 28590 45892 28642
rect 45724 28588 45892 28590
rect 45836 28420 45892 28588
rect 45836 28354 45892 28364
rect 45948 28196 46004 30156
rect 46172 30146 46228 30156
rect 45836 28140 46004 28196
rect 46060 28532 46116 28542
rect 45612 27076 45668 27086
rect 45612 26982 45668 27020
rect 45500 26238 45502 26290
rect 45554 26238 45556 26290
rect 45500 26226 45556 26238
rect 45836 25956 45892 28140
rect 46060 27858 46116 28476
rect 46060 27806 46062 27858
rect 46114 27806 46116 27858
rect 46060 27794 46116 27806
rect 46060 27076 46116 27086
rect 45164 25678 45166 25730
rect 45218 25678 45220 25730
rect 45164 25666 45220 25678
rect 45724 25900 45892 25956
rect 45948 27074 46116 27076
rect 45948 27022 46062 27074
rect 46114 27022 46116 27074
rect 45948 27020 46116 27022
rect 45948 26292 46004 27020
rect 46060 27010 46116 27020
rect 46284 26908 46340 32396
rect 46060 26852 46116 26862
rect 46172 26852 46340 26908
rect 46396 31556 46452 31566
rect 46116 26796 46228 26852
rect 46060 26516 46116 26796
rect 46284 26740 46340 26750
rect 46060 26460 46228 26516
rect 45612 25620 45668 25630
rect 45612 25526 45668 25564
rect 44940 25106 44996 25116
rect 45052 25282 45108 25294
rect 45052 25230 45054 25282
rect 45106 25230 45108 25282
rect 44828 24612 44884 24622
rect 44828 24162 44884 24556
rect 44828 24110 44830 24162
rect 44882 24110 44884 24162
rect 44828 24098 44884 24110
rect 45052 23828 45108 25230
rect 45164 24052 45220 24062
rect 45164 24050 45332 24052
rect 45164 23998 45166 24050
rect 45218 23998 45332 24050
rect 45164 23996 45332 23998
rect 45164 23986 45220 23996
rect 44380 23538 44436 23548
rect 44940 23826 45108 23828
rect 44940 23774 45054 23826
rect 45106 23774 45108 23826
rect 44940 23772 45108 23774
rect 44156 23314 44212 23324
rect 43820 22932 43876 22942
rect 43820 22594 43876 22876
rect 43820 22542 43822 22594
rect 43874 22542 43876 22594
rect 43820 22530 43876 22542
rect 43708 22484 43764 22494
rect 43708 22390 43764 22428
rect 44044 22370 44100 22382
rect 44044 22318 44046 22370
rect 44098 22318 44100 22370
rect 44044 21028 44100 22318
rect 44156 22258 44212 22270
rect 44156 22206 44158 22258
rect 44210 22206 44212 22258
rect 44156 21700 44212 22206
rect 44156 21634 44212 21644
rect 44268 21588 44324 21598
rect 44044 20962 44100 20972
rect 44156 21476 44212 21486
rect 43596 20738 43652 20748
rect 43484 20692 43540 20702
rect 43484 20598 43540 20636
rect 43260 19852 43372 19908
rect 42588 18676 42644 18686
rect 42588 17890 42644 18620
rect 42588 17838 42590 17890
rect 42642 17838 42644 17890
rect 42588 17826 42644 17838
rect 42700 18452 42756 18462
rect 42700 17778 42756 18396
rect 42700 17726 42702 17778
rect 42754 17726 42756 17778
rect 42700 17714 42756 17726
rect 43036 17666 43092 17678
rect 43036 17614 43038 17666
rect 43090 17614 43092 17666
rect 42476 17054 42478 17106
rect 42530 17054 42532 17106
rect 42476 17042 42532 17054
rect 42700 17220 42756 17230
rect 42700 17106 42756 17164
rect 42700 17054 42702 17106
rect 42754 17054 42756 17106
rect 42700 17042 42756 17054
rect 43036 17108 43092 17614
rect 43260 17666 43316 19852
rect 43372 19842 43428 19852
rect 44156 20468 44212 21420
rect 43484 19124 43540 19134
rect 43484 19030 43540 19068
rect 44156 18562 44212 20412
rect 44268 20802 44324 21532
rect 44940 21476 44996 23772
rect 45052 23762 45108 23772
rect 45052 23604 45108 23614
rect 45052 22482 45108 23548
rect 45276 23268 45332 23996
rect 45388 23268 45444 23278
rect 45276 23266 45444 23268
rect 45276 23214 45390 23266
rect 45442 23214 45444 23266
rect 45276 23212 45444 23214
rect 45388 23202 45444 23212
rect 45052 22430 45054 22482
rect 45106 22430 45108 22482
rect 45052 22418 45108 22430
rect 45612 22484 45668 22494
rect 45724 22484 45780 25900
rect 45836 24052 45892 24062
rect 45948 24052 46004 26236
rect 46172 25618 46228 26460
rect 46172 25566 46174 25618
rect 46226 25566 46228 25618
rect 46172 25554 46228 25566
rect 46060 25508 46116 25518
rect 46060 25414 46116 25452
rect 46060 25284 46116 25294
rect 46060 24612 46116 25228
rect 46172 24612 46228 24622
rect 46060 24610 46228 24612
rect 46060 24558 46174 24610
rect 46226 24558 46228 24610
rect 46060 24556 46228 24558
rect 46172 24546 46228 24556
rect 46060 24164 46116 24174
rect 46060 24070 46116 24108
rect 45836 24050 46004 24052
rect 45836 23998 45838 24050
rect 45890 23998 46004 24050
rect 45836 23996 46004 23998
rect 46172 24052 46228 24062
rect 46284 24052 46340 26684
rect 46172 24050 46340 24052
rect 46172 23998 46174 24050
rect 46226 23998 46340 24050
rect 46172 23996 46340 23998
rect 45836 23986 45892 23996
rect 46172 23986 46228 23996
rect 46396 23828 46452 31500
rect 45612 22482 45780 22484
rect 45612 22430 45614 22482
rect 45666 22430 45780 22482
rect 45612 22428 45780 22430
rect 45836 23772 46452 23828
rect 46508 28420 46564 28430
rect 45612 22418 45668 22428
rect 45836 22258 45892 23772
rect 46060 23156 46116 23166
rect 46060 23062 46116 23100
rect 45836 22206 45838 22258
rect 45890 22206 45892 22258
rect 45836 22194 45892 22206
rect 46172 22260 46228 22270
rect 46228 22204 46340 22260
rect 46172 22166 46228 22204
rect 45276 22148 45332 22158
rect 44940 21410 44996 21420
rect 45052 21924 45108 21934
rect 44268 20750 44270 20802
rect 44322 20750 44324 20802
rect 44268 19236 44324 20750
rect 44940 21028 44996 21038
rect 44828 20692 44884 20702
rect 44828 20598 44884 20636
rect 44716 19906 44772 19918
rect 44716 19854 44718 19906
rect 44770 19854 44772 19906
rect 44716 19236 44772 19854
rect 44268 19234 44772 19236
rect 44268 19182 44270 19234
rect 44322 19182 44772 19234
rect 44268 19180 44772 19182
rect 44268 19170 44324 19180
rect 44156 18510 44158 18562
rect 44210 18510 44212 18562
rect 44156 18498 44212 18510
rect 43820 18452 43876 18462
rect 43820 18338 43876 18396
rect 43820 18286 43822 18338
rect 43874 18286 43876 18338
rect 43820 18274 43876 18286
rect 44380 18450 44436 18462
rect 44380 18398 44382 18450
rect 44434 18398 44436 18450
rect 44380 18228 44436 18398
rect 44604 18340 44660 18350
rect 44380 18162 44436 18172
rect 44492 18338 44660 18340
rect 44492 18286 44606 18338
rect 44658 18286 44660 18338
rect 44492 18284 44660 18286
rect 43372 17780 43428 17790
rect 43372 17778 43652 17780
rect 43372 17726 43374 17778
rect 43426 17726 43652 17778
rect 43372 17724 43652 17726
rect 43372 17714 43428 17724
rect 43260 17614 43262 17666
rect 43314 17614 43316 17666
rect 43260 17602 43316 17614
rect 43484 17442 43540 17454
rect 43484 17390 43486 17442
rect 43538 17390 43540 17442
rect 43484 17332 43540 17390
rect 43484 17266 43540 17276
rect 43036 17042 43092 17052
rect 43372 17220 43428 17230
rect 42252 16830 42254 16882
rect 42306 16830 42308 16882
rect 42252 16818 42308 16830
rect 42924 16882 42980 16894
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42588 16772 42644 16782
rect 42588 16678 42644 16716
rect 40796 16098 41188 16100
rect 40796 16046 40798 16098
rect 40850 16046 41188 16098
rect 40796 16044 41188 16046
rect 40796 16034 40852 16044
rect 41132 15426 41188 16044
rect 41804 16034 41860 16044
rect 42924 15988 42980 16830
rect 43372 16882 43428 17164
rect 43372 16830 43374 16882
rect 43426 16830 43428 16882
rect 43372 16818 43428 16830
rect 43596 16436 43652 17724
rect 44492 17668 44548 18284
rect 44604 18274 44660 18284
rect 44044 17612 44548 17668
rect 43596 16370 43652 16380
rect 43708 17554 43764 17566
rect 43708 17502 43710 17554
rect 43762 17502 43764 17554
rect 42924 15540 42980 15932
rect 43596 16210 43652 16222
rect 43596 16158 43598 16210
rect 43650 16158 43652 16210
rect 43596 16100 43652 16158
rect 42924 15484 43316 15540
rect 41132 15374 41134 15426
rect 41186 15374 41188 15426
rect 40236 15204 40292 15214
rect 40124 15202 40292 15204
rect 40124 15150 40238 15202
rect 40290 15150 40292 15202
rect 40124 15148 40292 15150
rect 38892 15090 38948 15102
rect 38892 15038 38894 15090
rect 38946 15038 38948 15090
rect 38892 13858 38948 15038
rect 38892 13806 38894 13858
rect 38946 13806 38948 13858
rect 38892 13794 38948 13806
rect 39228 15090 39284 15102
rect 39228 15038 39230 15090
rect 39282 15038 39284 15090
rect 39228 13858 39284 15038
rect 40236 14532 40292 15148
rect 39564 14420 39620 14430
rect 39564 13970 39620 14364
rect 39564 13918 39566 13970
rect 39618 13918 39620 13970
rect 39564 13906 39620 13918
rect 40236 13972 40292 14476
rect 41132 15204 41188 15374
rect 42812 15428 42868 15438
rect 41132 14530 41188 15148
rect 42700 15316 42756 15326
rect 42700 14642 42756 15260
rect 42700 14590 42702 14642
rect 42754 14590 42756 14642
rect 42700 14578 42756 14590
rect 41132 14478 41134 14530
rect 41186 14478 41188 14530
rect 41132 14466 41188 14478
rect 40460 14420 40516 14430
rect 40460 14326 40516 14364
rect 41692 14418 41748 14430
rect 41692 14366 41694 14418
rect 41746 14366 41748 14418
rect 41692 14308 41748 14366
rect 42700 14420 42756 14430
rect 41692 14242 41748 14252
rect 41804 14306 41860 14318
rect 41804 14254 41806 14306
rect 41858 14254 41860 14306
rect 41804 13972 41860 14254
rect 42028 14308 42084 14318
rect 42028 14306 42532 14308
rect 42028 14254 42030 14306
rect 42082 14254 42532 14306
rect 42028 14252 42532 14254
rect 42028 14242 42084 14252
rect 40236 13906 40292 13916
rect 41244 13916 41860 13972
rect 39228 13806 39230 13858
rect 39282 13806 39284 13858
rect 39228 13794 39284 13806
rect 40348 13860 40404 13870
rect 41244 13860 41300 13916
rect 40348 13858 41300 13860
rect 40348 13806 40350 13858
rect 40402 13806 41246 13858
rect 41298 13806 41300 13858
rect 40348 13804 41300 13806
rect 40348 13794 40404 13804
rect 41244 13794 41300 13804
rect 40012 13748 40068 13758
rect 39900 13746 40068 13748
rect 39900 13694 40014 13746
rect 40066 13694 40068 13746
rect 39900 13692 40068 13694
rect 39900 13188 39956 13692
rect 40012 13682 40068 13692
rect 41132 13636 41188 13646
rect 39340 13132 39956 13188
rect 40012 13412 40068 13422
rect 38780 13074 39172 13076
rect 38780 13022 38782 13074
rect 38834 13022 39172 13074
rect 38780 13020 39172 13022
rect 38780 13010 38836 13020
rect 38892 12740 38948 12750
rect 38892 12738 39060 12740
rect 38892 12686 38894 12738
rect 38946 12686 39060 12738
rect 38892 12684 39060 12686
rect 38892 12674 38948 12684
rect 38444 12124 38724 12180
rect 37716 11788 37940 11844
rect 38108 12066 38164 12078
rect 38108 12014 38110 12066
rect 38162 12014 38164 12066
rect 38108 11788 38164 12014
rect 38220 11956 38276 11966
rect 38220 11954 38612 11956
rect 38220 11902 38222 11954
rect 38274 11902 38612 11954
rect 38220 11900 38612 11902
rect 38220 11890 38276 11900
rect 37660 11778 37716 11788
rect 37996 11732 38164 11788
rect 38220 11732 38276 11742
rect 37660 11620 37716 11630
rect 37548 11564 37660 11620
rect 37436 11554 37492 11564
rect 37660 11554 37716 11564
rect 37100 11508 37156 11518
rect 37100 11506 37380 11508
rect 37100 11454 37102 11506
rect 37154 11454 37380 11506
rect 37100 11452 37380 11454
rect 37100 11442 37156 11452
rect 37324 11396 37380 11452
rect 37772 11506 37828 11518
rect 37772 11454 37774 11506
rect 37826 11454 37828 11506
rect 37660 11396 37716 11434
rect 37772 11396 37828 11454
rect 37324 11340 37660 11396
rect 37716 11340 37828 11396
rect 37660 11330 37716 11340
rect 36988 10882 37044 10892
rect 37100 11284 37156 11294
rect 37884 11284 37940 11294
rect 36876 10668 37044 10724
rect 36540 10546 36596 10556
rect 36764 10610 36820 10622
rect 36764 10558 36766 10610
rect 36818 10558 36820 10610
rect 35980 10500 36036 10510
rect 35868 10498 36372 10500
rect 35868 10446 35982 10498
rect 36034 10446 36372 10498
rect 35868 10444 36372 10446
rect 35980 10434 36036 10444
rect 36316 10388 36372 10444
rect 36764 10388 36820 10558
rect 36316 10332 36820 10388
rect 34972 9100 35140 9156
rect 34972 8932 35028 8942
rect 34748 8206 34750 8258
rect 34802 8206 34804 8258
rect 34748 8194 34804 8206
rect 34860 8930 35028 8932
rect 34860 8878 34974 8930
rect 35026 8878 35028 8930
rect 34860 8876 35028 8878
rect 33964 8148 34020 8158
rect 33964 8036 34020 8092
rect 33964 7980 34244 8036
rect 34076 7812 34132 7822
rect 34076 7698 34132 7756
rect 34076 7646 34078 7698
rect 34130 7646 34132 7698
rect 34076 7634 34132 7646
rect 33964 7588 34020 7598
rect 33740 7532 33964 7588
rect 33964 7494 34020 7532
rect 34188 7476 34244 7980
rect 34300 8034 34356 8046
rect 34300 7982 34302 8034
rect 34354 7982 34356 8034
rect 34300 7700 34356 7982
rect 34860 7924 34916 8876
rect 34972 8866 35028 8876
rect 35084 8820 35140 9100
rect 35756 9090 35812 9100
rect 36092 9826 36148 9838
rect 36092 9774 36094 9826
rect 36146 9774 36148 9826
rect 35084 8484 35140 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35532 8484 35588 8494
rect 35084 8428 35364 8484
rect 34300 7634 34356 7644
rect 34524 7868 34916 7924
rect 35084 8260 35140 8270
rect 35084 8146 35140 8204
rect 35308 8258 35364 8428
rect 35308 8206 35310 8258
rect 35362 8206 35364 8258
rect 35308 8194 35364 8206
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 35084 7924 35140 8094
rect 34524 7698 34580 7868
rect 35084 7858 35140 7868
rect 34524 7646 34526 7698
rect 34578 7646 34580 7698
rect 34524 7634 34580 7646
rect 35084 7700 35140 7710
rect 34412 7476 34468 7486
rect 34188 7474 34468 7476
rect 34188 7422 34414 7474
rect 34466 7422 34468 7474
rect 34188 7420 34468 7422
rect 34412 7410 34468 7420
rect 34524 7364 34580 7374
rect 34412 7252 34468 7262
rect 33964 6916 34020 6926
rect 33628 6626 33684 6636
rect 33852 6804 33908 6814
rect 33740 6466 33796 6478
rect 33740 6414 33742 6466
rect 33794 6414 33796 6466
rect 33740 6244 33796 6414
rect 33740 6178 33796 6188
rect 33516 6078 33518 6130
rect 33570 6078 33572 6130
rect 33180 5908 33236 5918
rect 33180 5814 33236 5852
rect 32732 5506 32788 5516
rect 33404 5794 33460 5806
rect 33404 5742 33406 5794
rect 33458 5742 33460 5794
rect 33404 5348 33460 5742
rect 32396 5292 33460 5348
rect 32284 5012 32340 5022
rect 32284 4562 32340 4956
rect 32284 4510 32286 4562
rect 32338 4510 32340 4562
rect 32284 4498 32340 4510
rect 32396 4450 32452 5292
rect 32396 4398 32398 4450
rect 32450 4398 32452 4450
rect 32396 4386 32452 4398
rect 33068 5124 33124 5134
rect 33068 4338 33124 5068
rect 33516 5012 33572 6078
rect 33740 6020 33796 6030
rect 33852 6020 33908 6748
rect 33740 6018 33908 6020
rect 33740 5966 33742 6018
rect 33794 5966 33908 6018
rect 33740 5964 33908 5966
rect 33740 5954 33796 5964
rect 33852 5234 33908 5964
rect 33852 5182 33854 5234
rect 33906 5182 33908 5234
rect 33852 5170 33908 5182
rect 33516 4946 33572 4956
rect 33852 4452 33908 4462
rect 33964 4452 34020 6860
rect 34300 5908 34356 5918
rect 34300 5348 34356 5852
rect 34300 5122 34356 5292
rect 34300 5070 34302 5122
rect 34354 5070 34356 5122
rect 34300 5058 34356 5070
rect 34412 5122 34468 7196
rect 34524 5234 34580 7308
rect 34860 7362 34916 7374
rect 34860 7310 34862 7362
rect 34914 7310 34916 7362
rect 34524 5182 34526 5234
rect 34578 5182 34580 5234
rect 34524 5170 34580 5182
rect 34636 5796 34692 5806
rect 34412 5070 34414 5122
rect 34466 5070 34468 5122
rect 34412 5058 34468 5070
rect 34636 5124 34692 5740
rect 34860 5236 34916 7310
rect 35084 6916 35140 7644
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6860 35364 6916
rect 35308 5908 35364 6860
rect 35308 5842 35364 5852
rect 35420 5796 35476 5806
rect 35532 5796 35588 8428
rect 36092 8484 36148 9774
rect 36092 8418 36148 8428
rect 36988 8258 37044 10668
rect 37100 10610 37156 11228
rect 37772 11228 37884 11284
rect 37212 11170 37268 11182
rect 37660 11172 37716 11182
rect 37212 11118 37214 11170
rect 37266 11118 37268 11170
rect 37212 10948 37268 11118
rect 37436 11170 37716 11172
rect 37436 11118 37662 11170
rect 37714 11118 37716 11170
rect 37436 11116 37716 11118
rect 37212 10882 37268 10892
rect 37324 11060 37380 11070
rect 37100 10558 37102 10610
rect 37154 10558 37156 10610
rect 37100 10546 37156 10558
rect 37100 9604 37156 9614
rect 37100 9510 37156 9548
rect 37100 9044 37156 9054
rect 37100 8930 37156 8988
rect 37100 8878 37102 8930
rect 37154 8878 37156 8930
rect 37100 8866 37156 8878
rect 36988 8206 36990 8258
rect 37042 8206 37044 8258
rect 36988 8194 37044 8206
rect 37212 8260 37268 8270
rect 37212 8166 37268 8204
rect 36092 8146 36148 8158
rect 36092 8094 36094 8146
rect 36146 8094 36148 8146
rect 36092 6804 36148 8094
rect 36204 8036 36260 8046
rect 36204 8034 36372 8036
rect 36204 7982 36206 8034
rect 36258 7982 36372 8034
rect 36204 7980 36372 7982
rect 36204 7970 36260 7980
rect 36092 6738 36148 6748
rect 36204 6692 36260 6702
rect 36204 6598 36260 6636
rect 35476 5740 35588 5796
rect 35644 6578 35700 6590
rect 35644 6526 35646 6578
rect 35698 6526 35700 6578
rect 35420 5730 35476 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34860 5170 34916 5180
rect 35196 5348 35252 5358
rect 34636 5058 34692 5068
rect 34748 5122 34804 5134
rect 34748 5070 34750 5122
rect 34802 5070 34804 5122
rect 34524 5012 34580 5022
rect 34524 4900 34580 4956
rect 34636 4900 34692 4910
rect 34524 4898 34692 4900
rect 34524 4846 34638 4898
rect 34690 4846 34692 4898
rect 34524 4844 34692 4846
rect 34636 4834 34692 4844
rect 33852 4450 34020 4452
rect 33852 4398 33854 4450
rect 33906 4398 34020 4450
rect 33852 4396 34020 4398
rect 33852 4386 33908 4396
rect 33068 4286 33070 4338
rect 33122 4286 33124 4338
rect 33068 4274 33124 4286
rect 34748 4228 34804 5070
rect 35196 5122 35252 5292
rect 35420 5236 35476 5246
rect 35644 5236 35700 6526
rect 36092 6580 36148 6590
rect 35420 5234 35700 5236
rect 35420 5182 35422 5234
rect 35474 5182 35700 5234
rect 35420 5180 35700 5182
rect 35756 6466 35812 6478
rect 35756 6414 35758 6466
rect 35810 6414 35812 6466
rect 35420 5170 35476 5180
rect 35196 5070 35198 5122
rect 35250 5070 35252 5122
rect 35196 5058 35252 5070
rect 35644 5012 35700 5022
rect 35644 4918 35700 4956
rect 35420 4900 35476 4910
rect 35420 4806 35476 4844
rect 35756 4452 35812 6414
rect 35980 5348 36036 5358
rect 35868 5012 35924 5022
rect 35868 4918 35924 4956
rect 35980 4452 36036 5292
rect 35756 4386 35812 4396
rect 35868 4396 36036 4452
rect 32172 4172 32564 4228
rect 31612 4162 31668 4172
rect 31612 3668 31668 3678
rect 31500 3666 31668 3668
rect 31500 3614 31614 3666
rect 31666 3614 31668 3666
rect 31500 3612 31668 3614
rect 28700 3502 28702 3554
rect 28754 3502 28756 3554
rect 28700 3490 28756 3502
rect 26348 3390 26350 3442
rect 26402 3390 26404 3442
rect 26348 3378 26404 3390
rect 27804 3444 27860 3454
rect 26012 3278 26014 3330
rect 26066 3278 26068 3330
rect 26012 3266 26068 3278
rect 26236 3332 26292 3342
rect 26236 800 26292 3276
rect 27020 3332 27076 3342
rect 27020 3238 27076 3276
rect 27804 800 27860 3388
rect 29372 3444 29428 3454
rect 29372 800 29428 3388
rect 30940 800 30996 3612
rect 31612 3602 31668 3612
rect 32172 3556 32228 3566
rect 32172 3462 32228 3500
rect 32508 800 32564 4172
rect 34748 4162 34804 4172
rect 34076 4116 34132 4126
rect 33740 3444 33796 3482
rect 33740 3378 33796 3388
rect 34076 800 34132 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35868 3780 35924 4396
rect 35980 4228 36036 4238
rect 35980 4004 36036 4172
rect 35980 3938 36036 3948
rect 35420 3724 35924 3780
rect 35980 3780 36036 3790
rect 35196 3556 35252 3566
rect 35196 3462 35252 3500
rect 35420 3442 35476 3724
rect 35980 3554 36036 3724
rect 35980 3502 35982 3554
rect 36034 3502 36036 3554
rect 35980 3490 36036 3502
rect 35420 3390 35422 3442
rect 35474 3390 35476 3442
rect 35420 3378 35476 3390
rect 36092 980 36148 6524
rect 36316 6132 36372 7980
rect 37100 8034 37156 8046
rect 37100 7982 37102 8034
rect 37154 7982 37156 8034
rect 36988 7588 37044 7598
rect 37100 7588 37156 7982
rect 36988 7586 37156 7588
rect 36988 7534 36990 7586
rect 37042 7534 37156 7586
rect 36988 7532 37156 7534
rect 36988 7522 37044 7532
rect 37324 7476 37380 11004
rect 37436 10722 37492 11116
rect 37660 11106 37716 11116
rect 37772 11170 37828 11228
rect 37884 11218 37940 11228
rect 37772 11118 37774 11170
rect 37826 11118 37828 11170
rect 37436 10670 37438 10722
rect 37490 10670 37492 10722
rect 37436 10052 37492 10670
rect 37436 9986 37492 9996
rect 37548 10612 37604 10622
rect 37436 9604 37492 9614
rect 37436 8258 37492 9548
rect 37548 9042 37604 10556
rect 37772 10610 37828 11118
rect 37772 10558 37774 10610
rect 37826 10558 37828 10610
rect 37772 10546 37828 10558
rect 37996 11170 38052 11732
rect 38220 11394 38276 11676
rect 38220 11342 38222 11394
rect 38274 11342 38276 11394
rect 38220 11330 38276 11342
rect 38332 11396 38388 11406
rect 37996 11118 37998 11170
rect 38050 11118 38052 11170
rect 37660 10500 37716 10510
rect 37660 10406 37716 10444
rect 37996 10276 38052 11118
rect 38220 11172 38276 11182
rect 38220 10722 38276 11116
rect 38332 10834 38388 11340
rect 38556 11394 38612 11900
rect 38556 11342 38558 11394
rect 38610 11342 38612 11394
rect 38556 11330 38612 11342
rect 38668 11284 38724 12124
rect 38780 11506 38836 11518
rect 38780 11454 38782 11506
rect 38834 11454 38836 11506
rect 38780 11396 38836 11454
rect 38780 11330 38836 11340
rect 39004 11394 39060 12684
rect 39116 12402 39172 13020
rect 39340 12850 39396 13132
rect 39340 12798 39342 12850
rect 39394 12798 39396 12850
rect 39116 12350 39118 12402
rect 39170 12350 39172 12402
rect 39116 12338 39172 12350
rect 39228 12738 39284 12750
rect 39228 12686 39230 12738
rect 39282 12686 39284 12738
rect 39228 11732 39284 12686
rect 39228 11666 39284 11676
rect 39004 11342 39006 11394
rect 39058 11342 39060 11394
rect 39004 11330 39060 11342
rect 39116 11620 39172 11630
rect 39116 11394 39172 11564
rect 39116 11342 39118 11394
rect 39170 11342 39172 11394
rect 39116 11330 39172 11342
rect 38668 11218 38724 11228
rect 38780 11170 38836 11182
rect 38780 11118 38782 11170
rect 38834 11118 38836 11170
rect 38780 11060 38836 11118
rect 38780 10994 38836 11004
rect 39340 11060 39396 12798
rect 39452 12964 39508 12974
rect 39452 12178 39508 12908
rect 39900 12850 39956 12862
rect 39900 12798 39902 12850
rect 39954 12798 39956 12850
rect 39788 12740 39844 12750
rect 39788 12646 39844 12684
rect 39452 12126 39454 12178
rect 39506 12126 39508 12178
rect 39452 12114 39508 12126
rect 39676 12066 39732 12078
rect 39676 12014 39678 12066
rect 39730 12014 39732 12066
rect 39452 11396 39508 11406
rect 39452 11302 39508 11340
rect 39340 10994 39396 11004
rect 38332 10782 38334 10834
rect 38386 10782 38388 10834
rect 38332 10770 38388 10782
rect 39452 10836 39508 10846
rect 39452 10742 39508 10780
rect 39228 10724 39284 10734
rect 38220 10670 38222 10722
rect 38274 10670 38276 10722
rect 38220 10658 38276 10670
rect 38780 10722 39284 10724
rect 38780 10670 39230 10722
rect 39282 10670 39284 10722
rect 38780 10668 39284 10670
rect 38332 10388 38388 10398
rect 37548 8990 37550 9042
rect 37602 8990 37604 9042
rect 37548 8978 37604 8990
rect 37772 10220 38052 10276
rect 38108 10386 38388 10388
rect 38108 10334 38334 10386
rect 38386 10334 38388 10386
rect 38108 10332 38388 10334
rect 37772 9044 37828 10220
rect 37884 9604 37940 9614
rect 37884 9510 37940 9548
rect 37772 8978 37828 8988
rect 37996 9044 38052 9054
rect 38108 9044 38164 10332
rect 38332 10322 38388 10332
rect 38332 9714 38388 9726
rect 38332 9662 38334 9714
rect 38386 9662 38388 9714
rect 37996 9042 38164 9044
rect 37996 8990 37998 9042
rect 38050 8990 38164 9042
rect 37996 8988 38164 8990
rect 38220 9602 38276 9614
rect 38220 9550 38222 9602
rect 38274 9550 38276 9602
rect 37996 8978 38052 8988
rect 37436 8206 37438 8258
rect 37490 8206 37492 8258
rect 37436 7700 37492 8206
rect 37660 8932 37716 8942
rect 38220 8932 38276 9550
rect 38332 9044 38388 9662
rect 38332 8978 38388 8988
rect 38668 9714 38724 9726
rect 38668 9662 38670 9714
rect 38722 9662 38724 9714
rect 37660 8258 37716 8876
rect 38108 8876 38276 8932
rect 37772 8820 37828 8830
rect 38108 8820 38164 8876
rect 38444 8820 38500 8830
rect 37772 8818 38164 8820
rect 37772 8766 37774 8818
rect 37826 8766 38164 8818
rect 37772 8764 38164 8766
rect 38332 8818 38500 8820
rect 38332 8766 38446 8818
rect 38498 8766 38500 8818
rect 38332 8764 38500 8766
rect 37772 8754 37828 8764
rect 37660 8206 37662 8258
rect 37714 8206 37716 8258
rect 37660 8194 37716 8206
rect 37884 8596 37940 8606
rect 37436 7634 37492 7644
rect 37324 7410 37380 7420
rect 37660 7474 37716 7486
rect 37660 7422 37662 7474
rect 37714 7422 37716 7474
rect 36428 6916 36484 6926
rect 36428 6578 36484 6860
rect 36428 6526 36430 6578
rect 36482 6526 36484 6578
rect 36428 6514 36484 6526
rect 36316 6066 36372 6076
rect 37212 6468 37268 6478
rect 36204 5796 36260 5806
rect 36204 5124 36260 5740
rect 36316 5236 36372 5246
rect 36316 5142 36372 5180
rect 36204 4340 36260 5068
rect 36988 5124 37044 5134
rect 36988 5030 37044 5068
rect 36428 4898 36484 4910
rect 36428 4846 36430 4898
rect 36482 4846 36484 4898
rect 36316 4340 36372 4350
rect 36204 4338 36372 4340
rect 36204 4286 36318 4338
rect 36370 4286 36372 4338
rect 36204 4284 36372 4286
rect 36316 4274 36372 4284
rect 36428 3444 36484 4846
rect 37100 4452 37156 4462
rect 37100 4358 37156 4396
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 36428 3378 36484 3388
rect 35644 924 36148 980
rect 35644 800 35700 924
rect 37212 800 37268 6412
rect 37660 5124 37716 7422
rect 37772 6580 37828 6590
rect 37772 6486 37828 6524
rect 37884 5460 37940 8540
rect 37996 8258 38052 8270
rect 37996 8206 37998 8258
rect 38050 8206 38052 8258
rect 37996 7028 38052 8206
rect 38332 8260 38388 8764
rect 38444 8754 38500 8764
rect 38668 8370 38724 9662
rect 38668 8318 38670 8370
rect 38722 8318 38724 8370
rect 38668 8306 38724 8318
rect 38556 8260 38612 8270
rect 38332 8258 38612 8260
rect 38332 8206 38558 8258
rect 38610 8206 38612 8258
rect 38332 8204 38612 8206
rect 38556 8194 38612 8204
rect 38780 8260 38836 10668
rect 39228 10658 39284 10668
rect 39564 10612 39620 10622
rect 39564 10518 39620 10556
rect 38892 10498 38948 10510
rect 38892 10446 38894 10498
rect 38946 10446 38948 10498
rect 38892 10052 38948 10446
rect 39004 10388 39060 10398
rect 39004 10386 39172 10388
rect 39004 10334 39006 10386
rect 39058 10334 39172 10386
rect 39004 10332 39172 10334
rect 39004 10322 39060 10332
rect 38892 9986 38948 9996
rect 39004 10164 39060 10174
rect 38892 9828 38948 9866
rect 38892 9762 38948 9772
rect 39004 9714 39060 10108
rect 39004 9662 39006 9714
rect 39058 9662 39060 9714
rect 39004 9650 39060 9662
rect 39004 9492 39060 9502
rect 38892 8484 38948 8494
rect 38892 8390 38948 8428
rect 38780 8166 38836 8204
rect 38556 7924 38612 7934
rect 38556 7698 38612 7868
rect 39004 7812 39060 9436
rect 39116 9380 39172 10332
rect 39452 9940 39508 9950
rect 39452 9826 39508 9884
rect 39452 9774 39454 9826
rect 39506 9774 39508 9826
rect 39452 9762 39508 9774
rect 39676 9716 39732 12014
rect 39900 11396 39956 12798
rect 40012 12178 40068 13356
rect 40684 12964 40740 12974
rect 40684 12870 40740 12908
rect 41132 12962 41188 13580
rect 41132 12910 41134 12962
rect 41186 12910 41188 12962
rect 41132 12898 41188 12910
rect 41356 12962 41412 13916
rect 41916 13860 41972 13870
rect 41468 13748 41524 13758
rect 41468 13654 41524 13692
rect 41804 13748 41860 13758
rect 41692 13636 41748 13646
rect 41580 13580 41692 13636
rect 41580 12964 41636 13580
rect 41692 13570 41748 13580
rect 41804 13634 41860 13692
rect 41804 13582 41806 13634
rect 41858 13582 41860 13634
rect 41804 13570 41860 13582
rect 41356 12910 41358 12962
rect 41410 12910 41412 12962
rect 40348 12850 40404 12862
rect 40348 12798 40350 12850
rect 40402 12798 40404 12850
rect 40236 12738 40292 12750
rect 40236 12686 40238 12738
rect 40290 12686 40292 12738
rect 40012 12126 40014 12178
rect 40066 12126 40068 12178
rect 40012 12114 40068 12126
rect 40124 12292 40180 12302
rect 40236 12292 40292 12686
rect 40124 12290 40292 12292
rect 40124 12238 40126 12290
rect 40178 12238 40292 12290
rect 40124 12236 40292 12238
rect 40124 11508 40180 12236
rect 40348 12180 40404 12798
rect 40796 12850 40852 12862
rect 40796 12798 40798 12850
rect 40850 12798 40852 12850
rect 40796 12404 40852 12798
rect 40796 12348 41300 12404
rect 41132 12180 41188 12190
rect 40348 12178 41188 12180
rect 40348 12126 41134 12178
rect 41186 12126 41188 12178
rect 40348 12124 41188 12126
rect 40684 11508 40740 11518
rect 40124 11442 40180 11452
rect 40572 11506 40740 11508
rect 40572 11454 40686 11506
rect 40738 11454 40740 11506
rect 40572 11452 40740 11454
rect 39676 9650 39732 9660
rect 39788 11340 39956 11396
rect 40236 11396 40292 11406
rect 39564 9604 39620 9614
rect 39116 9324 39284 9380
rect 39116 9154 39172 9166
rect 39116 9102 39118 9154
rect 39170 9102 39172 9154
rect 39116 9044 39172 9102
rect 39116 8978 39172 8988
rect 39004 7746 39060 7756
rect 38556 7646 38558 7698
rect 38610 7646 38612 7698
rect 38556 7634 38612 7646
rect 39228 7588 39284 9324
rect 39340 9268 39396 9278
rect 39340 9174 39396 9212
rect 39564 9266 39620 9548
rect 39564 9214 39566 9266
rect 39618 9214 39620 9266
rect 39564 9202 39620 9214
rect 39788 9268 39844 11340
rect 40124 11284 40180 11294
rect 40236 11284 40292 11340
rect 40124 11282 40292 11284
rect 40124 11230 40126 11282
rect 40178 11230 40292 11282
rect 40124 11228 40292 11230
rect 40124 11218 40180 11228
rect 39900 11170 39956 11182
rect 39900 11118 39902 11170
rect 39954 11118 39956 11170
rect 39900 10948 39956 11118
rect 40012 11170 40068 11182
rect 40012 11118 40014 11170
rect 40066 11118 40068 11170
rect 40012 10948 40068 11118
rect 40012 10892 40180 10948
rect 39900 10882 39956 10892
rect 40012 10722 40068 10734
rect 40012 10670 40014 10722
rect 40066 10670 40068 10722
rect 39900 10386 39956 10398
rect 39900 10334 39902 10386
rect 39954 10334 39956 10386
rect 39900 9828 39956 10334
rect 40012 10052 40068 10670
rect 40012 9986 40068 9996
rect 39900 9762 39956 9772
rect 40012 9826 40068 9838
rect 40012 9774 40014 9826
rect 40066 9774 40068 9826
rect 40012 9716 40068 9774
rect 40124 9828 40180 10892
rect 40348 10612 40404 10622
rect 40124 9762 40180 9772
rect 40236 10386 40292 10398
rect 40236 10334 40238 10386
rect 40290 10334 40292 10386
rect 40012 9650 40068 9660
rect 39900 9268 39956 9278
rect 40236 9268 40292 10334
rect 40348 9604 40404 10556
rect 40460 9828 40516 9838
rect 40460 9734 40516 9772
rect 40348 9548 40516 9604
rect 39788 9266 40068 9268
rect 39788 9214 39902 9266
rect 39954 9214 40068 9266
rect 39788 9212 40068 9214
rect 39900 9202 39956 9212
rect 39452 8932 39508 8942
rect 39788 8932 39844 8942
rect 39452 8930 39732 8932
rect 39452 8878 39454 8930
rect 39506 8878 39732 8930
rect 39452 8876 39732 8878
rect 39452 8866 39508 8876
rect 39676 8596 39732 8876
rect 39788 8838 39844 8876
rect 40012 8932 40068 9212
rect 40236 9202 40292 9212
rect 40012 8866 40068 8876
rect 40124 9042 40180 9054
rect 40124 8990 40126 9042
rect 40178 8990 40180 9042
rect 40124 8820 40180 8990
rect 40124 8754 40180 8764
rect 40348 9042 40404 9054
rect 40348 8990 40350 9042
rect 40402 8990 40404 9042
rect 39676 8540 40292 8596
rect 40124 8370 40180 8382
rect 40124 8318 40126 8370
rect 40178 8318 40180 8370
rect 39228 7522 39284 7532
rect 39676 8260 39732 8270
rect 39676 7586 39732 8204
rect 40012 8258 40068 8270
rect 40012 8206 40014 8258
rect 40066 8206 40068 8258
rect 39676 7534 39678 7586
rect 39730 7534 39732 7586
rect 39676 7522 39732 7534
rect 39788 7924 39844 7934
rect 37996 6962 38052 6972
rect 38332 7474 38388 7486
rect 38332 7422 38334 7474
rect 38386 7422 38388 7474
rect 37884 5394 37940 5404
rect 37772 5348 37828 5358
rect 37772 5234 37828 5292
rect 37772 5182 37774 5234
rect 37826 5182 37828 5234
rect 37772 5170 37828 5182
rect 37660 5058 37716 5068
rect 38332 4788 38388 7422
rect 38332 4722 38388 4732
rect 38444 7474 38500 7486
rect 38444 7422 38446 7474
rect 38498 7422 38500 7474
rect 38444 7028 38500 7422
rect 38668 7476 38724 7486
rect 38668 7474 38836 7476
rect 38668 7422 38670 7474
rect 38722 7422 38836 7474
rect 38668 7420 38836 7422
rect 38668 7410 38724 7420
rect 38444 3444 38500 6972
rect 38780 4900 38836 7420
rect 38892 7474 38948 7486
rect 38892 7422 38894 7474
rect 38946 7422 38948 7474
rect 38892 7028 38948 7422
rect 39564 7476 39620 7486
rect 39340 7364 39396 7374
rect 39340 7270 39396 7308
rect 39228 7252 39284 7262
rect 39228 7158 39284 7196
rect 38892 6962 38948 6972
rect 39452 6690 39508 6702
rect 39452 6638 39454 6690
rect 39506 6638 39508 6690
rect 39452 6356 39508 6638
rect 39228 6300 39452 6356
rect 39228 5796 39284 6300
rect 39452 6290 39508 6300
rect 39452 6020 39508 6030
rect 39228 5730 39284 5740
rect 39340 5964 39452 6020
rect 38780 4834 38836 4844
rect 39228 4900 39284 4910
rect 38892 4788 38948 4798
rect 38892 4004 38948 4732
rect 38892 3778 38948 3948
rect 39228 4226 39284 4844
rect 39228 4174 39230 4226
rect 39282 4174 39284 4226
rect 39228 4004 39284 4174
rect 39228 3938 39284 3948
rect 38892 3726 38894 3778
rect 38946 3726 38948 3778
rect 38892 3714 38948 3726
rect 39228 3780 39284 3790
rect 39340 3780 39396 5964
rect 39452 5954 39508 5964
rect 39564 5906 39620 7420
rect 39788 6916 39844 7868
rect 40012 7698 40068 8206
rect 40012 7646 40014 7698
rect 40066 7646 40068 7698
rect 40012 7634 40068 7646
rect 39900 7588 39956 7598
rect 39900 7494 39956 7532
rect 39788 6860 39956 6916
rect 39564 5854 39566 5906
rect 39618 5854 39620 5906
rect 39564 5842 39620 5854
rect 39788 6692 39844 6702
rect 39788 5236 39844 6636
rect 39900 5908 39956 6860
rect 40012 6578 40068 6590
rect 40012 6526 40014 6578
rect 40066 6526 40068 6578
rect 40012 6132 40068 6526
rect 40124 6356 40180 8318
rect 40236 7586 40292 8540
rect 40236 7534 40238 7586
rect 40290 7534 40292 7586
rect 40236 7522 40292 7534
rect 40348 7028 40404 8990
rect 40460 7140 40516 9548
rect 40572 7364 40628 11452
rect 40684 11442 40740 11452
rect 41020 11282 41076 11294
rect 41020 11230 41022 11282
rect 41074 11230 41076 11282
rect 40796 11170 40852 11182
rect 40796 11118 40798 11170
rect 40850 11118 40852 11170
rect 40796 10836 40852 11118
rect 41020 11172 41076 11230
rect 41020 11106 41076 11116
rect 40796 10770 40852 10780
rect 41132 10612 41188 12124
rect 41244 12178 41300 12348
rect 41356 12290 41412 12910
rect 41356 12238 41358 12290
rect 41410 12238 41412 12290
rect 41356 12226 41412 12238
rect 41468 12908 41636 12964
rect 41244 12126 41246 12178
rect 41298 12126 41300 12178
rect 41244 11732 41300 12126
rect 41244 11666 41300 11676
rect 41356 11508 41412 11518
rect 41356 11414 41412 11452
rect 41468 10834 41524 12908
rect 41580 12738 41636 12750
rect 41580 12686 41582 12738
rect 41634 12686 41636 12738
rect 41580 11844 41636 12686
rect 41580 11778 41636 11788
rect 41692 12738 41748 12750
rect 41692 12686 41694 12738
rect 41746 12686 41748 12738
rect 41580 11620 41636 11630
rect 41692 11620 41748 12686
rect 41804 12180 41860 12190
rect 41916 12180 41972 13804
rect 42476 13858 42532 14252
rect 42476 13806 42478 13858
rect 42530 13806 42532 13858
rect 42140 13746 42196 13758
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 13524 42196 13694
rect 42364 13748 42420 13758
rect 42364 13654 42420 13692
rect 42476 13524 42532 13806
rect 42140 13458 42196 13468
rect 42364 13468 42532 13524
rect 42588 14306 42644 14318
rect 42588 14254 42590 14306
rect 42642 14254 42644 14306
rect 42364 13074 42420 13468
rect 42364 13022 42366 13074
rect 42418 13022 42420 13074
rect 42364 13010 42420 13022
rect 42476 12964 42532 12974
rect 42476 12870 42532 12908
rect 42364 12292 42420 12302
rect 41804 12178 41972 12180
rect 41804 12126 41806 12178
rect 41858 12126 41972 12178
rect 41804 12124 41972 12126
rect 42252 12290 42420 12292
rect 42252 12238 42366 12290
rect 42418 12238 42420 12290
rect 42252 12236 42420 12238
rect 41804 12114 41860 12124
rect 42028 11954 42084 11966
rect 42028 11902 42030 11954
rect 42082 11902 42084 11954
rect 41916 11732 41972 11742
rect 41580 11618 41748 11620
rect 41580 11566 41582 11618
rect 41634 11566 41748 11618
rect 41580 11564 41748 11566
rect 41804 11676 41916 11732
rect 41580 11554 41636 11564
rect 41468 10782 41470 10834
rect 41522 10782 41524 10834
rect 41468 10770 41524 10782
rect 41244 10612 41300 10622
rect 41132 10610 41300 10612
rect 41132 10558 41246 10610
rect 41298 10558 41300 10610
rect 41132 10556 41300 10558
rect 40796 9826 40852 9838
rect 40796 9774 40798 9826
rect 40850 9774 40852 9826
rect 40796 9716 40852 9774
rect 40796 9650 40852 9660
rect 41020 9826 41076 9838
rect 41020 9774 41022 9826
rect 41074 9774 41076 9826
rect 40684 9604 40740 9614
rect 40684 9510 40740 9548
rect 40908 9156 40964 9166
rect 40684 9154 40964 9156
rect 40684 9102 40910 9154
rect 40962 9102 40964 9154
rect 40684 9100 40964 9102
rect 40684 8148 40740 9100
rect 40908 9090 40964 9100
rect 40908 8820 40964 8830
rect 40908 8370 40964 8764
rect 41020 8708 41076 9774
rect 41132 9492 41188 9502
rect 41132 9266 41188 9436
rect 41132 9214 41134 9266
rect 41186 9214 41188 9266
rect 41132 9202 41188 9214
rect 41020 8652 41188 8708
rect 41020 8484 41076 8494
rect 41132 8484 41188 8652
rect 41020 8482 41188 8484
rect 41020 8430 41022 8482
rect 41074 8430 41188 8482
rect 41020 8428 41188 8430
rect 41020 8418 41076 8428
rect 40908 8318 40910 8370
rect 40962 8318 40964 8370
rect 40908 8306 40964 8318
rect 41244 8372 41300 10556
rect 41692 9828 41748 9838
rect 41804 9828 41860 11676
rect 41916 11666 41972 11676
rect 41916 11396 41972 11406
rect 41916 11302 41972 11340
rect 42028 11172 42084 11902
rect 42028 11106 42084 11116
rect 42140 10612 42196 10622
rect 42028 10498 42084 10510
rect 42028 10446 42030 10498
rect 42082 10446 42084 10498
rect 42028 9940 42084 10446
rect 42028 9874 42084 9884
rect 42140 9938 42196 10556
rect 42252 10276 42308 12236
rect 42364 12226 42420 12236
rect 42364 11394 42420 11406
rect 42364 11342 42366 11394
rect 42418 11342 42420 11394
rect 42364 11172 42420 11342
rect 42476 11396 42532 11406
rect 42476 11302 42532 11340
rect 42364 11106 42420 11116
rect 42252 10210 42308 10220
rect 42364 10836 42420 10846
rect 42364 10722 42420 10780
rect 42364 10670 42366 10722
rect 42418 10670 42420 10722
rect 42140 9886 42142 9938
rect 42194 9886 42196 9938
rect 42140 9874 42196 9886
rect 41692 9826 41860 9828
rect 41692 9774 41694 9826
rect 41746 9774 41860 9826
rect 41692 9772 41860 9774
rect 42364 9828 42420 10670
rect 42588 10612 42644 14254
rect 42700 12852 42756 14364
rect 42812 13076 42868 15372
rect 42924 14420 42980 14430
rect 42924 13970 42980 14364
rect 43148 14418 43204 14430
rect 43148 14366 43150 14418
rect 43202 14366 43204 14418
rect 42924 13918 42926 13970
rect 42978 13918 42980 13970
rect 42924 13906 42980 13918
rect 43036 14306 43092 14318
rect 43036 14254 43038 14306
rect 43090 14254 43092 14306
rect 43036 13636 43092 14254
rect 43036 13570 43092 13580
rect 43148 13412 43204 14366
rect 43260 13634 43316 15484
rect 43260 13582 43262 13634
rect 43314 13582 43316 13634
rect 43260 13570 43316 13582
rect 43372 15316 43428 15326
rect 43148 13346 43204 13356
rect 42812 13010 42868 13020
rect 43148 12964 43204 12974
rect 43148 12870 43204 12908
rect 42700 12796 42980 12852
rect 42812 12290 42868 12302
rect 42812 12238 42814 12290
rect 42866 12238 42868 12290
rect 42700 11394 42756 11406
rect 42700 11342 42702 11394
rect 42754 11342 42756 11394
rect 42700 11284 42756 11342
rect 42700 11218 42756 11228
rect 42588 10518 42644 10556
rect 42812 10052 42868 12238
rect 42924 11618 42980 12796
rect 43260 12068 43316 12078
rect 43372 12068 43428 15260
rect 43596 13412 43652 16044
rect 43708 15316 43764 17502
rect 44044 16994 44100 17612
rect 44044 16942 44046 16994
rect 44098 16942 44100 16994
rect 44044 16930 44100 16942
rect 44156 17442 44212 17454
rect 44156 17390 44158 17442
rect 44210 17390 44212 17442
rect 44044 15988 44100 15998
rect 44044 15894 44100 15932
rect 43708 15250 43764 15260
rect 43932 15874 43988 15886
rect 43932 15822 43934 15874
rect 43986 15822 43988 15874
rect 43932 15148 43988 15822
rect 44156 15540 44212 17390
rect 44716 17220 44772 19180
rect 44940 19234 44996 20972
rect 45052 20020 45108 21868
rect 45164 21364 45220 21374
rect 45164 21026 45220 21308
rect 45164 20974 45166 21026
rect 45218 20974 45220 21026
rect 45164 20188 45220 20974
rect 45276 21026 45332 22092
rect 46172 22036 46228 22046
rect 45948 21980 46172 22036
rect 45388 21700 45444 21710
rect 45388 21606 45444 21644
rect 45276 20974 45278 21026
rect 45330 20974 45332 21026
rect 45276 20962 45332 20974
rect 45948 20914 46004 21980
rect 46172 21970 46228 21980
rect 46060 21588 46116 21598
rect 46060 21494 46116 21532
rect 46284 21588 46340 22204
rect 46284 21522 46340 21532
rect 45948 20862 45950 20914
rect 46002 20862 46004 20914
rect 45948 20850 46004 20862
rect 45164 20132 45780 20188
rect 45052 19964 45220 20020
rect 45164 19684 45220 19964
rect 45164 19628 45444 19684
rect 45276 19460 45332 19470
rect 44940 19182 44942 19234
rect 44994 19182 44996 19234
rect 44940 19170 44996 19182
rect 45164 19236 45220 19246
rect 45164 19142 45220 19180
rect 44828 19124 44884 19134
rect 44828 19030 44884 19068
rect 44940 18564 44996 18574
rect 44828 18562 44996 18564
rect 44828 18510 44942 18562
rect 44994 18510 44996 18562
rect 44828 18508 44996 18510
rect 44828 18450 44884 18508
rect 44940 18498 44996 18508
rect 45164 18562 45220 18574
rect 45164 18510 45166 18562
rect 45218 18510 45220 18562
rect 44828 18398 44830 18450
rect 44882 18398 44884 18450
rect 44828 18386 44884 18398
rect 45164 18452 45220 18510
rect 45276 18562 45332 19404
rect 45276 18510 45278 18562
rect 45330 18510 45332 18562
rect 45276 18498 45332 18510
rect 45164 18386 45220 18396
rect 44940 18340 44996 18350
rect 44940 17780 44996 18284
rect 45388 18116 45444 19628
rect 45724 19458 45780 20132
rect 45724 19406 45726 19458
rect 45778 19406 45780 19458
rect 45724 19394 45780 19406
rect 45948 19348 46004 19358
rect 45836 19236 45892 19246
rect 45836 19142 45892 19180
rect 45948 19122 46004 19292
rect 45948 19070 45950 19122
rect 46002 19070 46004 19122
rect 45948 19058 46004 19070
rect 45724 18338 45780 18350
rect 46172 18340 46228 18350
rect 45724 18286 45726 18338
rect 45778 18286 45780 18338
rect 45612 18228 45668 18238
rect 45612 18134 45668 18172
rect 45388 18050 45444 18060
rect 44940 17686 44996 17724
rect 45388 17780 45444 17790
rect 45388 17686 45444 17724
rect 44828 17220 44884 17230
rect 44716 17164 44828 17220
rect 44828 17154 44884 17164
rect 44828 16772 44884 16782
rect 44828 16210 44884 16716
rect 45724 16322 45780 18286
rect 45948 18284 46172 18340
rect 45836 17444 45892 17454
rect 45836 17350 45892 17388
rect 45724 16270 45726 16322
rect 45778 16270 45780 16322
rect 45724 16258 45780 16270
rect 44828 16158 44830 16210
rect 44882 16158 44884 16210
rect 44828 16146 44884 16158
rect 45276 16212 45332 16222
rect 45276 16118 45332 16156
rect 45836 16212 45892 16222
rect 45948 16212 46004 18284
rect 46172 18246 46228 18284
rect 46172 18116 46228 18126
rect 46172 17556 46228 18060
rect 46508 17780 46564 28364
rect 46620 24500 46676 35644
rect 46620 24434 46676 24444
rect 46844 22036 46900 39340
rect 46844 21970 46900 21980
rect 46508 17714 46564 17724
rect 46172 17554 46340 17556
rect 46172 17502 46174 17554
rect 46226 17502 46340 17554
rect 46172 17500 46340 17502
rect 46172 17490 46228 17500
rect 45836 16210 46004 16212
rect 45836 16158 45838 16210
rect 45890 16158 46004 16210
rect 45836 16156 46004 16158
rect 46060 17220 46116 17230
rect 44940 15876 44996 15886
rect 45388 15876 45444 15886
rect 44940 15874 45332 15876
rect 44940 15822 44942 15874
rect 44994 15822 45332 15874
rect 44940 15820 45332 15822
rect 44940 15810 44996 15820
rect 44156 15474 44212 15484
rect 43820 15092 43988 15148
rect 45276 15148 45332 15820
rect 45388 15874 45556 15876
rect 45388 15822 45390 15874
rect 45442 15822 45556 15874
rect 45388 15820 45556 15822
rect 45388 15810 45444 15820
rect 45276 15092 45444 15148
rect 43708 14420 43764 14430
rect 43708 14326 43764 14364
rect 43596 13346 43652 13356
rect 43484 13076 43540 13086
rect 43484 12962 43540 13020
rect 43484 12910 43486 12962
rect 43538 12910 43540 12962
rect 43484 12180 43540 12910
rect 43708 12964 43764 12974
rect 43708 12870 43764 12908
rect 43484 12114 43540 12124
rect 43260 12066 43428 12068
rect 43260 12014 43262 12066
rect 43314 12014 43428 12066
rect 43260 12012 43428 12014
rect 43260 12002 43316 12012
rect 43820 11732 43876 15092
rect 43820 11666 43876 11676
rect 43932 14476 44212 14532
rect 42924 11566 42926 11618
rect 42978 11566 42980 11618
rect 42924 11554 42980 11566
rect 43372 11620 43428 11630
rect 43036 11396 43092 11406
rect 43036 11302 43092 11340
rect 42812 9986 42868 9996
rect 42924 11172 42980 11182
rect 42924 10050 42980 11116
rect 43260 11060 43316 11070
rect 43260 10498 43316 11004
rect 43260 10446 43262 10498
rect 43314 10446 43316 10498
rect 43260 10434 43316 10446
rect 42924 9998 42926 10050
rect 42978 9998 42980 10050
rect 42924 9986 42980 9998
rect 42700 9828 42756 9838
rect 42364 9826 42756 9828
rect 42364 9774 42366 9826
rect 42418 9774 42702 9826
rect 42754 9774 42756 9826
rect 42364 9772 42756 9774
rect 41356 9492 41412 9502
rect 41356 9266 41412 9436
rect 41356 9214 41358 9266
rect 41410 9214 41412 9266
rect 41356 9202 41412 9214
rect 41468 9268 41524 9278
rect 41692 9268 41748 9772
rect 42364 9762 42420 9772
rect 41468 9266 41748 9268
rect 41468 9214 41470 9266
rect 41522 9214 41748 9266
rect 41468 9212 41748 9214
rect 41804 9602 41860 9614
rect 41804 9550 41806 9602
rect 41858 9550 41860 9602
rect 41804 9268 41860 9550
rect 41468 9202 41524 9212
rect 41804 9202 41860 9212
rect 41916 9604 41972 9614
rect 41468 9044 41524 9054
rect 41356 8988 41468 9044
rect 41916 9044 41972 9548
rect 42252 9044 42308 9054
rect 41916 9042 42308 9044
rect 41916 8990 42254 9042
rect 42306 8990 42308 9042
rect 41916 8988 42308 8990
rect 41356 8930 41412 8988
rect 41468 8978 41524 8988
rect 41356 8878 41358 8930
rect 41410 8878 41412 8930
rect 41356 8866 41412 8878
rect 41356 8372 41412 8382
rect 41244 8370 41412 8372
rect 41244 8318 41358 8370
rect 41410 8318 41412 8370
rect 41244 8316 41412 8318
rect 41356 8306 41412 8316
rect 41244 8148 41300 8158
rect 40684 8092 40964 8148
rect 40572 7298 40628 7308
rect 40908 7140 40964 8092
rect 41300 8092 41412 8148
rect 41244 8082 41300 8092
rect 41132 7924 41188 7934
rect 41020 7140 41076 7150
rect 40460 7084 40852 7140
rect 40908 7084 41020 7140
rect 40348 6972 40628 7028
rect 40460 6804 40516 6814
rect 40460 6690 40516 6748
rect 40460 6638 40462 6690
rect 40514 6638 40516 6690
rect 40460 6626 40516 6638
rect 40236 6578 40292 6590
rect 40236 6526 40238 6578
rect 40290 6526 40292 6578
rect 40236 6468 40292 6526
rect 40236 6412 40516 6468
rect 40124 6300 40292 6356
rect 40012 6076 40180 6132
rect 40012 5908 40068 5918
rect 39900 5906 40068 5908
rect 39900 5854 40014 5906
rect 40066 5854 40068 5906
rect 39900 5852 40068 5854
rect 40012 5842 40068 5852
rect 40124 5908 40180 6076
rect 40236 6130 40292 6300
rect 40460 6244 40516 6412
rect 40460 6178 40516 6188
rect 40236 6078 40238 6130
rect 40290 6078 40292 6130
rect 40236 6066 40292 6078
rect 40572 6132 40628 6972
rect 40684 6690 40740 6702
rect 40684 6638 40686 6690
rect 40738 6638 40740 6690
rect 40684 6468 40740 6638
rect 40684 6402 40740 6412
rect 40796 6466 40852 7084
rect 41020 7074 41076 7084
rect 40908 6692 40964 6702
rect 40908 6598 40964 6636
rect 40796 6414 40798 6466
rect 40850 6414 40852 6466
rect 40796 6402 40852 6414
rect 41020 6580 41076 6590
rect 41020 6356 41076 6524
rect 40908 6300 41076 6356
rect 40572 6076 40852 6132
rect 40348 6020 40404 6030
rect 40348 5926 40404 5964
rect 39900 5236 39956 5246
rect 39788 5234 39956 5236
rect 39788 5182 39902 5234
rect 39954 5182 39956 5234
rect 39788 5180 39956 5182
rect 39900 5170 39956 5180
rect 40124 5012 40180 5852
rect 40796 5796 40852 6076
rect 40908 6020 40964 6300
rect 41020 6132 41076 6142
rect 41020 6038 41076 6076
rect 41132 6130 41188 7868
rect 41356 6916 41412 8092
rect 41132 6078 41134 6130
rect 41186 6078 41188 6130
rect 41132 6066 41188 6078
rect 41244 6132 41300 6142
rect 41356 6132 41412 6860
rect 41244 6130 41412 6132
rect 41244 6078 41246 6130
rect 41298 6078 41412 6130
rect 41244 6076 41412 6078
rect 41468 7812 41524 7822
rect 40908 5954 40964 5964
rect 41244 5796 41300 6076
rect 41468 5906 41524 7756
rect 41692 7140 41748 7150
rect 41468 5854 41470 5906
rect 41522 5854 41524 5906
rect 41468 5842 41524 5854
rect 41580 6692 41636 6702
rect 39900 4956 40180 5012
rect 40572 5348 40628 5358
rect 39228 3778 39396 3780
rect 39228 3726 39230 3778
rect 39282 3726 39396 3778
rect 39228 3724 39396 3726
rect 39564 4114 39620 4126
rect 39564 4062 39566 4114
rect 39618 4062 39620 4114
rect 39228 3714 39284 3724
rect 38444 3378 38500 3388
rect 38780 3668 38836 3678
rect 38780 800 38836 3612
rect 39564 3556 39620 4062
rect 39900 3668 39956 4956
rect 40460 4900 40516 4910
rect 40124 4898 40516 4900
rect 40124 4846 40462 4898
rect 40514 4846 40516 4898
rect 40124 4844 40516 4846
rect 40124 4450 40180 4844
rect 40460 4834 40516 4844
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 4386 40180 4398
rect 40012 4338 40068 4350
rect 40012 4286 40014 4338
rect 40066 4286 40068 4338
rect 40012 4228 40068 4286
rect 40348 4340 40404 4350
rect 40572 4340 40628 5292
rect 40796 5348 40852 5740
rect 41020 5740 41300 5796
rect 40796 5346 40964 5348
rect 40796 5294 40798 5346
rect 40850 5294 40964 5346
rect 40796 5292 40964 5294
rect 40796 5282 40852 5292
rect 40348 4338 40628 4340
rect 40348 4286 40350 4338
rect 40402 4286 40628 4338
rect 40348 4284 40628 4286
rect 40796 4338 40852 4350
rect 40796 4286 40798 4338
rect 40850 4286 40852 4338
rect 40348 4274 40404 4284
rect 40012 4162 40068 4172
rect 40796 4228 40852 4286
rect 40908 4340 40964 5292
rect 41020 5234 41076 5740
rect 41020 5182 41022 5234
rect 41074 5182 41076 5234
rect 41020 4562 41076 5182
rect 41356 5236 41412 5246
rect 41580 5236 41636 6636
rect 41692 5908 41748 7084
rect 42028 7028 42084 7038
rect 41916 6690 41972 6702
rect 41916 6638 41918 6690
rect 41970 6638 41972 6690
rect 41916 6132 41972 6638
rect 41916 6066 41972 6076
rect 41692 5814 41748 5852
rect 41356 5234 41636 5236
rect 41356 5182 41358 5234
rect 41410 5182 41636 5234
rect 41356 5180 41636 5182
rect 41356 5170 41412 5180
rect 41020 4510 41022 4562
rect 41074 4510 41076 4562
rect 41020 4498 41076 4510
rect 41916 4900 41972 4910
rect 41132 4340 41188 4350
rect 40908 4338 41188 4340
rect 40908 4286 41134 4338
rect 41186 4286 41188 4338
rect 40908 4284 41188 4286
rect 41132 4274 41188 4284
rect 40796 4162 40852 4172
rect 41580 4228 41636 4238
rect 41580 4134 41636 4172
rect 40348 3892 40404 3902
rect 40124 3668 40180 3678
rect 39900 3666 40180 3668
rect 39900 3614 40126 3666
rect 40178 3614 40180 3666
rect 39900 3612 40180 3614
rect 40124 3602 40180 3612
rect 39564 3490 39620 3500
rect 39116 3444 39172 3454
rect 39116 3350 39172 3388
rect 40348 800 40404 3836
rect 41916 800 41972 4844
rect 42028 4338 42084 6972
rect 42140 6580 42196 6590
rect 42140 6486 42196 6524
rect 42252 6244 42308 8988
rect 42252 6018 42308 6188
rect 42252 5966 42254 6018
rect 42306 5966 42308 6018
rect 42252 5954 42308 5966
rect 42364 6916 42420 6926
rect 42364 6468 42420 6860
rect 42364 6018 42420 6412
rect 42364 5966 42366 6018
rect 42418 5966 42420 6018
rect 42364 5954 42420 5966
rect 42140 5908 42196 5918
rect 42140 5814 42196 5852
rect 42028 4286 42030 4338
rect 42082 4286 42084 4338
rect 42028 4274 42084 4286
rect 42252 5012 42308 5022
rect 42252 3666 42308 4956
rect 42476 4452 42532 4462
rect 42476 4358 42532 4396
rect 42588 4228 42644 9772
rect 42700 9762 42756 9772
rect 43260 9716 43316 9726
rect 42924 9714 43316 9716
rect 42924 9662 43262 9714
rect 43314 9662 43316 9714
rect 42924 9660 43316 9662
rect 42924 9156 42980 9660
rect 43260 9650 43316 9660
rect 42812 9100 42980 9156
rect 43036 9156 43092 9166
rect 42812 9042 42868 9100
rect 42812 8990 42814 9042
rect 42866 8990 42868 9042
rect 42812 6916 42868 8990
rect 42924 8930 42980 8942
rect 42924 8878 42926 8930
rect 42978 8878 42980 8930
rect 42924 8260 42980 8878
rect 42924 8194 42980 8204
rect 42812 6850 42868 6860
rect 42812 6692 42868 6702
rect 42812 6598 42868 6636
rect 42924 6580 42980 6590
rect 42924 6486 42980 6524
rect 42812 5796 42868 5806
rect 42812 5702 42868 5740
rect 43036 5572 43092 9100
rect 43260 8932 43316 8942
rect 43372 8932 43428 11564
rect 43820 11396 43876 11406
rect 43820 11302 43876 11340
rect 43596 11172 43652 11182
rect 43260 8930 43428 8932
rect 43260 8878 43262 8930
rect 43314 8878 43428 8930
rect 43260 8876 43428 8878
rect 43484 11170 43652 11172
rect 43484 11118 43598 11170
rect 43650 11118 43652 11170
rect 43484 11116 43652 11118
rect 43260 8866 43316 8876
rect 43260 8484 43316 8494
rect 43260 5794 43316 8428
rect 43484 8370 43540 11116
rect 43596 11106 43652 11116
rect 43932 9828 43988 14476
rect 44044 14306 44100 14318
rect 44044 14254 44046 14306
rect 44098 14254 44100 14306
rect 44044 12964 44100 14254
rect 44156 14308 44212 14476
rect 44828 14308 44884 14318
rect 45276 14308 45332 14318
rect 44156 14306 44884 14308
rect 44156 14254 44830 14306
rect 44882 14254 44884 14306
rect 44156 14252 44884 14254
rect 44828 14242 44884 14252
rect 44940 14306 45332 14308
rect 44940 14254 45278 14306
rect 45330 14254 45332 14306
rect 44940 14252 45332 14254
rect 44044 12898 44100 12908
rect 44044 12740 44100 12750
rect 44044 12738 44884 12740
rect 44044 12686 44046 12738
rect 44098 12686 44884 12738
rect 44044 12684 44884 12686
rect 44044 12674 44100 12684
rect 44716 12404 44772 12414
rect 44380 12348 44716 12404
rect 43820 9772 43988 9828
rect 44044 11284 44100 11294
rect 43596 9604 43652 9614
rect 43596 9510 43652 9548
rect 43484 8318 43486 8370
rect 43538 8318 43540 8370
rect 43484 8306 43540 8318
rect 43484 7364 43540 7374
rect 43540 7308 43652 7364
rect 43484 7298 43540 7308
rect 43596 6914 43652 7308
rect 43596 6862 43598 6914
rect 43650 6862 43652 6914
rect 43596 6850 43652 6862
rect 43708 6916 43764 6926
rect 43708 6822 43764 6860
rect 43260 5742 43262 5794
rect 43314 5742 43316 5794
rect 43260 5730 43316 5742
rect 43036 5516 43652 5572
rect 43484 5236 43540 5246
rect 43484 5142 43540 5180
rect 43372 5124 43428 5134
rect 43036 5068 43372 5124
rect 42700 4228 42756 4238
rect 42588 4172 42700 4228
rect 42700 4162 42756 4172
rect 42812 4226 42868 4238
rect 42812 4174 42814 4226
rect 42866 4174 42868 4226
rect 42812 4004 42868 4174
rect 42812 3938 42868 3948
rect 42924 4114 42980 4126
rect 42924 4062 42926 4114
rect 42978 4062 42980 4114
rect 42924 3892 42980 4062
rect 42924 3826 42980 3836
rect 42252 3614 42254 3666
rect 42306 3614 42308 3666
rect 42252 3602 42308 3614
rect 43036 3554 43092 5068
rect 43372 5058 43428 5068
rect 43596 4900 43652 5516
rect 43372 4844 43652 4900
rect 43260 4228 43316 4238
rect 43260 4134 43316 4172
rect 43036 3502 43038 3554
rect 43090 3502 43092 3554
rect 43036 3490 43092 3502
rect 43372 2772 43428 4844
rect 43708 3556 43764 3566
rect 43708 3462 43764 3500
rect 43820 3388 43876 9772
rect 43932 9602 43988 9614
rect 43932 9550 43934 9602
rect 43986 9550 43988 9602
rect 43932 9492 43988 9550
rect 43932 8484 43988 9436
rect 43932 8418 43988 8428
rect 44044 8260 44100 11228
rect 44268 8372 44324 8382
rect 44268 8260 44324 8316
rect 43932 8204 44100 8260
rect 44156 8258 44324 8260
rect 44156 8206 44270 8258
rect 44322 8206 44324 8258
rect 44156 8204 44324 8206
rect 43932 7028 43988 8204
rect 43932 6914 43988 6972
rect 43932 6862 43934 6914
rect 43986 6862 43988 6914
rect 43932 6850 43988 6862
rect 44044 7700 44100 7710
rect 44044 6916 44100 7644
rect 44156 7588 44212 8204
rect 44268 8194 44324 8204
rect 44156 7586 44324 7588
rect 44156 7534 44158 7586
rect 44210 7534 44324 7586
rect 44156 7532 44324 7534
rect 44156 7522 44212 7532
rect 44156 6916 44212 6926
rect 44044 6860 44156 6916
rect 44156 6822 44212 6860
rect 44044 6468 44100 6478
rect 44044 6374 44100 6412
rect 44268 5124 44324 7532
rect 44268 5030 44324 5068
rect 44380 5012 44436 12348
rect 44716 12338 44772 12348
rect 44492 12180 44548 12190
rect 44492 11788 44548 12124
rect 44492 11732 44772 11788
rect 44716 8372 44772 11732
rect 44828 11394 44884 12684
rect 44828 11342 44830 11394
rect 44882 11342 44884 11394
rect 44828 11330 44884 11342
rect 44828 9604 44884 9614
rect 44828 9510 44884 9548
rect 44828 8372 44884 8382
rect 44716 8370 44884 8372
rect 44716 8318 44830 8370
rect 44882 8318 44884 8370
rect 44716 8316 44884 8318
rect 44828 8306 44884 8316
rect 44940 8036 44996 14252
rect 45276 14242 45332 14252
rect 45388 13858 45444 15092
rect 45388 13806 45390 13858
rect 45442 13806 45444 13858
rect 45388 13794 45444 13806
rect 45500 13636 45556 15820
rect 45836 15314 45892 16156
rect 45836 15262 45838 15314
rect 45890 15262 45892 15314
rect 45836 15250 45892 15262
rect 45948 15204 46004 15214
rect 45388 13580 45556 13636
rect 45724 14306 45780 14318
rect 45724 14254 45726 14306
rect 45778 14254 45780 14306
rect 45276 12964 45332 12974
rect 45164 12738 45220 12750
rect 45164 12686 45166 12738
rect 45218 12686 45220 12738
rect 45164 12404 45220 12686
rect 45164 12338 45220 12348
rect 45276 12068 45332 12908
rect 45388 12290 45444 13580
rect 45500 12852 45556 12862
rect 45500 12850 45668 12852
rect 45500 12798 45502 12850
rect 45554 12798 45668 12850
rect 45500 12796 45668 12798
rect 45500 12786 45556 12796
rect 45388 12238 45390 12290
rect 45442 12238 45444 12290
rect 45388 12226 45444 12238
rect 45276 12012 45444 12068
rect 45164 11172 45220 11182
rect 45164 11170 45332 11172
rect 45164 11118 45166 11170
rect 45218 11118 45332 11170
rect 45164 11116 45332 11118
rect 45164 11106 45220 11116
rect 45164 9714 45220 9726
rect 45164 9662 45166 9714
rect 45218 9662 45220 9714
rect 45052 8260 45108 8270
rect 45052 8166 45108 8204
rect 44828 7980 44996 8036
rect 44716 7476 44772 7486
rect 44716 7382 44772 7420
rect 44828 5572 44884 7980
rect 44940 6802 44996 6814
rect 44940 6750 44942 6802
rect 44994 6750 44996 6802
rect 44940 5796 44996 6750
rect 45052 6804 45108 6814
rect 45052 6710 45108 6748
rect 45164 5908 45220 9662
rect 45276 9156 45332 11116
rect 45388 10722 45444 12012
rect 45388 10670 45390 10722
rect 45442 10670 45444 10722
rect 45388 10658 45444 10670
rect 45388 9156 45444 9166
rect 45276 9154 45444 9156
rect 45276 9102 45390 9154
rect 45442 9102 45444 9154
rect 45276 9100 45444 9102
rect 45388 9090 45444 9100
rect 45388 8260 45444 8270
rect 45388 8166 45444 8204
rect 45276 7028 45332 7038
rect 45276 6914 45332 6972
rect 45276 6862 45278 6914
rect 45330 6862 45332 6914
rect 45276 6850 45332 6862
rect 45500 6916 45556 6926
rect 45500 6822 45556 6860
rect 45612 6690 45668 12796
rect 45724 8372 45780 14254
rect 45836 13188 45892 13198
rect 45836 12850 45892 13132
rect 45836 12798 45838 12850
rect 45890 12798 45892 12850
rect 45836 12786 45892 12798
rect 45948 12180 46004 15148
rect 46060 13746 46116 17164
rect 46284 16884 46340 17500
rect 46284 16818 46340 16828
rect 46172 16770 46228 16782
rect 46172 16718 46174 16770
rect 46226 16718 46228 16770
rect 46172 16322 46228 16718
rect 46172 16270 46174 16322
rect 46226 16270 46228 16322
rect 46172 16258 46228 16270
rect 46060 13694 46062 13746
rect 46114 13694 46116 13746
rect 46060 13682 46116 13694
rect 46060 12962 46116 12974
rect 46060 12910 46062 12962
rect 46114 12910 46116 12962
rect 46060 12516 46116 12910
rect 46060 12450 46116 12460
rect 46060 12180 46116 12190
rect 45948 12178 46116 12180
rect 45948 12126 46062 12178
rect 46114 12126 46116 12178
rect 45948 12124 46116 12126
rect 46060 12114 46116 12124
rect 45836 11170 45892 11182
rect 45836 11118 45838 11170
rect 45890 11118 45892 11170
rect 45836 10724 45892 11118
rect 46172 11172 46228 11182
rect 46172 11170 46340 11172
rect 46172 11118 46174 11170
rect 46226 11118 46340 11170
rect 46172 11116 46340 11118
rect 46172 11106 46228 11116
rect 45836 10658 45892 10668
rect 46060 10610 46116 10622
rect 46060 10558 46062 10610
rect 46114 10558 46116 10610
rect 45836 9604 45892 9614
rect 45836 9510 45892 9548
rect 46060 9042 46116 10558
rect 46172 9714 46228 9726
rect 46172 9662 46174 9714
rect 46226 9662 46228 9714
rect 46172 9156 46228 9662
rect 46172 9090 46228 9100
rect 46060 8990 46062 9042
rect 46114 8990 46116 9042
rect 46060 8372 46116 8990
rect 45724 8316 45892 8372
rect 45612 6638 45614 6690
rect 45666 6638 45668 6690
rect 45612 6626 45668 6638
rect 45724 8034 45780 8046
rect 45724 7982 45726 8034
rect 45778 7982 45780 8034
rect 45724 6468 45780 7982
rect 45388 6412 45780 6468
rect 45388 6018 45444 6412
rect 45388 5966 45390 6018
rect 45442 5966 45444 6018
rect 45388 5954 45444 5966
rect 45164 5852 45332 5908
rect 45276 5796 45332 5852
rect 45276 5740 45444 5796
rect 44940 5730 44996 5740
rect 44380 4946 44436 4956
rect 44716 5516 44884 5572
rect 44604 4116 44660 4126
rect 44604 3778 44660 4060
rect 44604 3726 44606 3778
rect 44658 3726 44660 3778
rect 44604 3714 44660 3726
rect 44716 3388 44772 5516
rect 44828 5348 44884 5358
rect 44828 5234 44884 5292
rect 45388 5346 45444 5740
rect 45388 5294 45390 5346
rect 45442 5294 45444 5346
rect 45388 5282 45444 5294
rect 44828 5182 44830 5234
rect 44882 5182 44884 5234
rect 44828 5170 44884 5182
rect 45052 5122 45108 5134
rect 45052 5070 45054 5122
rect 45106 5070 45108 5122
rect 45052 4452 45108 5070
rect 45724 4900 45780 4910
rect 45500 4898 45780 4900
rect 45500 4846 45726 4898
rect 45778 4846 45780 4898
rect 45500 4844 45780 4846
rect 45052 4386 45108 4396
rect 45388 4452 45444 4462
rect 45500 4452 45556 4844
rect 45724 4834 45780 4844
rect 45836 4900 45892 8316
rect 46116 8316 46228 8372
rect 46060 8306 46116 8316
rect 45948 8260 46004 8270
rect 45948 8166 46004 8204
rect 45948 6468 46004 6478
rect 45948 5122 46004 6412
rect 46060 6466 46116 6478
rect 46060 6414 46062 6466
rect 46114 6414 46116 6466
rect 46060 6356 46116 6414
rect 46060 6290 46116 6300
rect 45948 5070 45950 5122
rect 46002 5070 46004 5122
rect 45948 5058 46004 5070
rect 46172 5906 46228 8316
rect 46284 8036 46340 11116
rect 46284 7970 46340 7980
rect 46172 5854 46174 5906
rect 46226 5854 46228 5906
rect 45836 4834 45892 4844
rect 45388 4450 45556 4452
rect 45388 4398 45390 4450
rect 45442 4398 45556 4450
rect 45388 4396 45556 4398
rect 45388 4386 45444 4396
rect 46172 4338 46228 5854
rect 46172 4286 46174 4338
rect 46226 4286 46228 4338
rect 46172 4274 46228 4286
rect 43372 2706 43428 2716
rect 43596 3332 43876 3388
rect 44492 3332 44772 3388
rect 43596 2436 43652 3332
rect 43484 2380 43652 2436
rect 43484 800 43540 2380
rect 44492 980 44548 3332
rect 44492 924 45108 980
rect 45052 800 45108 924
rect 2688 0 2800 800
rect 4256 0 4368 800
rect 5824 0 5936 800
rect 7392 0 7504 800
rect 8960 0 9072 800
rect 10528 0 10640 800
rect 12096 0 12208 800
rect 13664 0 13776 800
rect 15232 0 15344 800
rect 16800 0 16912 800
rect 18368 0 18480 800
rect 19936 0 20048 800
rect 21504 0 21616 800
rect 23072 0 23184 800
rect 24640 0 24752 800
rect 26208 0 26320 800
rect 27776 0 27888 800
rect 29344 0 29456 800
rect 30912 0 31024 800
rect 32480 0 32592 800
rect 34048 0 34160 800
rect 35616 0 35728 800
rect 37184 0 37296 800
rect 38752 0 38864 800
rect 40320 0 40432 800
rect 41888 0 42000 800
rect 43456 0 43568 800
rect 45024 0 45136 800
<< via2 >>
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 9548 43820 9604 43876
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 6076 41132 6132 41188
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 6076 39228 6132 39284
rect 2828 38946 2884 38948
rect 2828 38894 2830 38946
rect 2830 38894 2882 38946
rect 2882 38894 2884 38946
rect 2828 38892 2884 38894
rect 3500 38946 3556 38948
rect 3500 38894 3502 38946
rect 3502 38894 3554 38946
rect 3554 38894 3556 38946
rect 3500 38892 3556 38894
rect 3052 38722 3108 38724
rect 3052 38670 3054 38722
rect 3054 38670 3106 38722
rect 3106 38670 3108 38722
rect 3052 38668 3108 38670
rect 1820 37212 1876 37268
rect 1708 37154 1764 37156
rect 1708 37102 1710 37154
rect 1710 37102 1762 37154
rect 1762 37102 1764 37154
rect 1708 37100 1764 37102
rect 3388 37100 3444 37156
rect 3948 38668 4004 38724
rect 3612 38220 3668 38276
rect 3500 37884 3556 37940
rect 2828 36482 2884 36484
rect 2828 36430 2830 36482
rect 2830 36430 2882 36482
rect 2882 36430 2884 36482
rect 2828 36428 2884 36430
rect 3276 36482 3332 36484
rect 3276 36430 3278 36482
rect 3278 36430 3330 36482
rect 3330 36430 3332 36482
rect 3276 36428 3332 36430
rect 2828 34860 2884 34916
rect 2716 34130 2772 34132
rect 2716 34078 2718 34130
rect 2718 34078 2770 34130
rect 2770 34078 2772 34130
rect 2716 34076 2772 34078
rect 2156 33964 2212 34020
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4284 38220 4340 38276
rect 4172 37884 4228 37940
rect 3948 37100 4004 37156
rect 3388 36428 3444 36484
rect 3836 36258 3892 36260
rect 3836 36206 3838 36258
rect 3838 36206 3890 36258
rect 3890 36206 3892 36258
rect 3836 36204 3892 36206
rect 3836 35756 3892 35812
rect 3276 34914 3332 34916
rect 3276 34862 3278 34914
rect 3278 34862 3330 34914
rect 3330 34862 3332 34914
rect 3276 34860 3332 34862
rect 4620 37266 4676 37268
rect 4620 37214 4622 37266
rect 4622 37214 4674 37266
rect 4674 37214 4676 37266
rect 4620 37212 4676 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5068 38780 5124 38836
rect 6636 42924 6692 42980
rect 10108 43820 10164 43876
rect 6636 42588 6692 42644
rect 10108 43036 10164 43092
rect 9660 42754 9716 42756
rect 9660 42702 9662 42754
rect 9662 42702 9714 42754
rect 9714 42702 9716 42754
rect 9660 42700 9716 42702
rect 9548 42642 9604 42644
rect 9548 42590 9550 42642
rect 9550 42590 9602 42642
rect 9602 42590 9604 42642
rect 9548 42588 9604 42590
rect 9324 42028 9380 42084
rect 11900 44044 11956 44100
rect 9100 40348 9156 40404
rect 6860 39788 6916 39844
rect 7084 39394 7140 39396
rect 7084 39342 7086 39394
rect 7086 39342 7138 39394
rect 7138 39342 7140 39394
rect 7084 39340 7140 39342
rect 5180 37490 5236 37492
rect 5180 37438 5182 37490
rect 5182 37438 5234 37490
rect 5234 37438 5236 37490
rect 5180 37436 5236 37438
rect 5740 37266 5796 37268
rect 5740 37214 5742 37266
rect 5742 37214 5794 37266
rect 5794 37214 5796 37266
rect 5740 37212 5796 37214
rect 6412 38892 6468 38948
rect 4956 37042 5012 37044
rect 4956 36990 4958 37042
rect 4958 36990 5010 37042
rect 5010 36990 5012 37042
rect 4956 36988 5012 36990
rect 4732 35756 4788 35812
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 35026 4900 35028
rect 4844 34974 4846 35026
rect 4846 34974 4898 35026
rect 4898 34974 4900 35026
rect 4844 34972 4900 34974
rect 4396 34914 4452 34916
rect 4396 34862 4398 34914
rect 4398 34862 4450 34914
rect 4450 34862 4452 34914
rect 4396 34860 4452 34862
rect 4396 34242 4452 34244
rect 4396 34190 4398 34242
rect 4398 34190 4450 34242
rect 4450 34190 4452 34242
rect 4396 34188 4452 34190
rect 3052 34076 3108 34132
rect 2940 33964 2996 34020
rect 4508 34130 4564 34132
rect 4508 34078 4510 34130
rect 4510 34078 4562 34130
rect 4562 34078 4564 34130
rect 4508 34076 4564 34078
rect 3388 33964 3444 34020
rect 5852 36316 5908 36372
rect 5628 35644 5684 35700
rect 5740 35810 5796 35812
rect 5740 35758 5742 35810
rect 5742 35758 5794 35810
rect 5794 35758 5796 35810
rect 5740 35756 5796 35758
rect 5068 34860 5124 34916
rect 5292 35196 5348 35252
rect 5180 34188 5236 34244
rect 4844 33964 4900 34020
rect 5292 34130 5348 34132
rect 5292 34078 5294 34130
rect 5294 34078 5346 34130
rect 5346 34078 5348 34130
rect 5292 34076 5348 34078
rect 5964 35586 6020 35588
rect 5964 35534 5966 35586
rect 5966 35534 6018 35586
rect 6018 35534 6020 35586
rect 5964 35532 6020 35534
rect 7756 39340 7812 39396
rect 7756 38668 7812 38724
rect 8764 39394 8820 39396
rect 8764 39342 8766 39394
rect 8766 39342 8818 39394
rect 8818 39342 8820 39394
rect 8764 39340 8820 39342
rect 8652 38834 8708 38836
rect 8652 38782 8654 38834
rect 8654 38782 8706 38834
rect 8706 38782 8708 38834
rect 8652 38780 8708 38782
rect 7420 37996 7476 38052
rect 10108 41186 10164 41188
rect 10108 41134 10110 41186
rect 10110 41134 10162 41186
rect 10162 41134 10164 41186
rect 10108 41132 10164 41134
rect 8988 39340 9044 39396
rect 8988 38946 9044 38948
rect 8988 38894 8990 38946
rect 8990 38894 9042 38946
rect 9042 38894 9044 38946
rect 8988 38892 9044 38894
rect 9772 39394 9828 39396
rect 9772 39342 9774 39394
rect 9774 39342 9826 39394
rect 9826 39342 9828 39394
rect 9772 39340 9828 39342
rect 10108 39788 10164 39844
rect 10556 42028 10612 42084
rect 10332 40348 10388 40404
rect 11004 42978 11060 42980
rect 11004 42926 11006 42978
rect 11006 42926 11058 42978
rect 11058 42926 11060 42978
rect 11004 42924 11060 42926
rect 11676 42978 11732 42980
rect 11676 42926 11678 42978
rect 11678 42926 11730 42978
rect 11730 42926 11732 42978
rect 11676 42924 11732 42926
rect 10892 42754 10948 42756
rect 10892 42702 10894 42754
rect 10894 42702 10946 42754
rect 10946 42702 10948 42754
rect 10892 42700 10948 42702
rect 11452 42754 11508 42756
rect 11452 42702 11454 42754
rect 11454 42702 11506 42754
rect 11506 42702 11508 42754
rect 11452 42700 11508 42702
rect 13468 42978 13524 42980
rect 13468 42926 13470 42978
rect 13470 42926 13522 42978
rect 13522 42926 13524 42978
rect 13468 42924 13524 42926
rect 12460 42700 12516 42756
rect 10668 41132 10724 41188
rect 11788 41132 11844 41188
rect 11452 41020 11508 41076
rect 11116 39730 11172 39732
rect 11116 39678 11118 39730
rect 11118 39678 11170 39730
rect 11170 39678 11172 39730
rect 11116 39676 11172 39678
rect 11788 39842 11844 39844
rect 11788 39790 11790 39842
rect 11790 39790 11842 39842
rect 11842 39790 11844 39842
rect 11788 39788 11844 39790
rect 11676 39452 11732 39508
rect 9436 38668 9492 38724
rect 8764 37548 8820 37604
rect 9884 38444 9940 38500
rect 11900 39340 11956 39396
rect 12908 42642 12964 42644
rect 12908 42590 12910 42642
rect 12910 42590 12962 42642
rect 12962 42590 12964 42642
rect 12908 42588 12964 42590
rect 12796 41244 12852 41300
rect 13804 44098 13860 44100
rect 13804 44046 13806 44098
rect 13806 44046 13858 44098
rect 13858 44046 13860 44098
rect 13804 44044 13860 44046
rect 14588 44434 14644 44436
rect 14588 44382 14590 44434
rect 14590 44382 14642 44434
rect 14642 44382 14644 44434
rect 14588 44380 14644 44382
rect 15596 44434 15652 44436
rect 15596 44382 15598 44434
rect 15598 44382 15650 44434
rect 15650 44382 15652 44434
rect 15596 44380 15652 44382
rect 13916 42754 13972 42756
rect 13916 42702 13918 42754
rect 13918 42702 13970 42754
rect 13970 42702 13972 42754
rect 13916 42700 13972 42702
rect 13692 42588 13748 42644
rect 14028 42642 14084 42644
rect 14028 42590 14030 42642
rect 14030 42590 14082 42642
rect 14082 42590 14084 42642
rect 14028 42588 14084 42590
rect 13692 41804 13748 41860
rect 14028 41074 14084 41076
rect 14028 41022 14030 41074
rect 14030 41022 14082 41074
rect 14082 41022 14084 41074
rect 14028 41020 14084 41022
rect 12572 40290 12628 40292
rect 12572 40238 12574 40290
rect 12574 40238 12626 40290
rect 12626 40238 12628 40290
rect 12572 40236 12628 40238
rect 13468 40236 13524 40292
rect 12908 39618 12964 39620
rect 12908 39566 12910 39618
rect 12910 39566 12962 39618
rect 12962 39566 12964 39618
rect 12908 39564 12964 39566
rect 13468 39452 13524 39508
rect 13804 39506 13860 39508
rect 13804 39454 13806 39506
rect 13806 39454 13858 39506
rect 13858 39454 13860 39506
rect 13804 39452 13860 39454
rect 9996 38220 10052 38276
rect 11116 38220 11172 38276
rect 9884 38108 9940 38164
rect 8988 37490 9044 37492
rect 8988 37438 8990 37490
rect 8990 37438 9042 37490
rect 9042 37438 9044 37490
rect 8988 37436 9044 37438
rect 8204 37324 8260 37380
rect 8876 37378 8932 37380
rect 8876 37326 8878 37378
rect 8878 37326 8930 37378
rect 8930 37326 8932 37378
rect 8876 37324 8932 37326
rect 7756 36370 7812 36372
rect 7756 36318 7758 36370
rect 7758 36318 7810 36370
rect 7810 36318 7812 36370
rect 7756 36316 7812 36318
rect 6972 36204 7028 36260
rect 6748 35698 6804 35700
rect 6748 35646 6750 35698
rect 6750 35646 6802 35698
rect 6802 35646 6804 35698
rect 6748 35644 6804 35646
rect 6860 35586 6916 35588
rect 6860 35534 6862 35586
rect 6862 35534 6914 35586
rect 6914 35534 6916 35586
rect 6860 35532 6916 35534
rect 6524 35196 6580 35252
rect 6300 34860 6356 34916
rect 6524 34972 6580 35028
rect 7196 35196 7252 35252
rect 9548 37378 9604 37380
rect 9548 37326 9550 37378
rect 9550 37326 9602 37378
rect 9602 37326 9604 37378
rect 9548 37324 9604 37326
rect 8988 36258 9044 36260
rect 8988 36206 8990 36258
rect 8990 36206 9042 36258
rect 9042 36206 9044 36258
rect 8988 36204 9044 36206
rect 9324 37212 9380 37268
rect 8876 35532 8932 35588
rect 7868 35084 7924 35140
rect 8204 35196 8260 35252
rect 7756 34972 7812 35028
rect 7868 34914 7924 34916
rect 7868 34862 7870 34914
rect 7870 34862 7922 34914
rect 7922 34862 7924 34914
rect 7868 34860 7924 34862
rect 7308 34802 7364 34804
rect 7308 34750 7310 34802
rect 7310 34750 7362 34802
rect 7362 34750 7364 34802
rect 7308 34748 7364 34750
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5292 33628 5348 33684
rect 4620 33516 4676 33572
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4620 31890 4676 31892
rect 4620 31838 4622 31890
rect 4622 31838 4674 31890
rect 4674 31838 4676 31890
rect 4620 31836 4676 31838
rect 5516 31554 5572 31556
rect 5516 31502 5518 31554
rect 5518 31502 5570 31554
rect 5570 31502 5572 31554
rect 5516 31500 5572 31502
rect 6860 34242 6916 34244
rect 6860 34190 6862 34242
rect 6862 34190 6914 34242
rect 6914 34190 6916 34242
rect 6860 34188 6916 34190
rect 6412 34130 6468 34132
rect 6412 34078 6414 34130
rect 6414 34078 6466 34130
rect 6466 34078 6468 34130
rect 6412 34076 6468 34078
rect 6972 34130 7028 34132
rect 6972 34078 6974 34130
rect 6974 34078 7026 34130
rect 7026 34078 7028 34130
rect 6972 34076 7028 34078
rect 7756 34130 7812 34132
rect 7756 34078 7758 34130
rect 7758 34078 7810 34130
rect 7810 34078 7812 34130
rect 7756 34076 7812 34078
rect 8092 34076 8148 34132
rect 8764 35084 8820 35140
rect 8204 33964 8260 34020
rect 7532 33516 7588 33572
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5180 30492 5236 30548
rect 4396 30380 4452 30436
rect 2492 29932 2548 29988
rect 3164 30268 3220 30324
rect 1820 29708 1876 29764
rect 3276 30156 3332 30212
rect 1820 29260 1876 29316
rect 1708 28476 1764 28532
rect 2044 29202 2100 29204
rect 2044 29150 2046 29202
rect 2046 29150 2098 29202
rect 2098 29150 2100 29202
rect 2044 29148 2100 29150
rect 2044 28364 2100 28420
rect 1708 24892 1764 24948
rect 2604 28476 2660 28532
rect 3052 29426 3108 29428
rect 3052 29374 3054 29426
rect 3054 29374 3106 29426
rect 3106 29374 3108 29426
rect 3052 29372 3108 29374
rect 3836 30098 3892 30100
rect 3836 30046 3838 30098
rect 3838 30046 3890 30098
rect 3890 30046 3892 30098
rect 3836 30044 3892 30046
rect 4620 30268 4676 30324
rect 3724 29426 3780 29428
rect 3724 29374 3726 29426
rect 3726 29374 3778 29426
rect 3778 29374 3780 29426
rect 3724 29372 3780 29374
rect 4844 29372 4900 29428
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4956 28364 5012 28420
rect 2828 27916 2884 27972
rect 2604 27580 2660 27636
rect 2492 26572 2548 26628
rect 3500 27916 3556 27972
rect 3948 27858 4004 27860
rect 3948 27806 3950 27858
rect 3950 27806 4002 27858
rect 4002 27806 4004 27858
rect 3948 27804 4004 27806
rect 3276 27580 3332 27636
rect 4732 27634 4788 27636
rect 4732 27582 4734 27634
rect 4734 27582 4786 27634
rect 4786 27582 4788 27634
rect 4732 27580 4788 27582
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5740 31836 5796 31892
rect 5852 31388 5908 31444
rect 5740 30492 5796 30548
rect 5628 30268 5684 30324
rect 5852 30210 5908 30212
rect 5852 30158 5854 30210
rect 5854 30158 5906 30210
rect 5906 30158 5908 30210
rect 5852 30156 5908 30158
rect 5516 29484 5572 29540
rect 5740 30098 5796 30100
rect 5740 30046 5742 30098
rect 5742 30046 5794 30098
rect 5794 30046 5796 30098
rect 5740 30044 5796 30046
rect 5628 29148 5684 29204
rect 5740 28364 5796 28420
rect 5292 27970 5348 27972
rect 5292 27918 5294 27970
rect 5294 27918 5346 27970
rect 5346 27918 5348 27970
rect 5292 27916 5348 27918
rect 5516 27858 5572 27860
rect 5516 27806 5518 27858
rect 5518 27806 5570 27858
rect 5570 27806 5572 27858
rect 5516 27804 5572 27806
rect 3164 26796 3220 26852
rect 3052 26684 3108 26740
rect 3164 26514 3220 26516
rect 3164 26462 3166 26514
rect 3166 26462 3218 26514
rect 3218 26462 3220 26514
rect 3164 26460 3220 26462
rect 3836 26796 3892 26852
rect 3948 26572 4004 26628
rect 3164 25116 3220 25172
rect 3276 24946 3332 24948
rect 3276 24894 3278 24946
rect 3278 24894 3330 24946
rect 3330 24894 3332 24946
rect 3276 24892 3332 24894
rect 3948 25116 4004 25172
rect 2380 24668 2436 24724
rect 3164 24722 3220 24724
rect 3164 24670 3166 24722
rect 3166 24670 3218 24722
rect 3218 24670 3220 24722
rect 3164 24668 3220 24670
rect 4620 26514 4676 26516
rect 4620 26462 4622 26514
rect 4622 26462 4674 26514
rect 4674 26462 4676 26514
rect 4620 26460 4676 26462
rect 5852 26684 5908 26740
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4508 25676 4564 25732
rect 3836 24444 3892 24500
rect 5964 27804 6020 27860
rect 5740 26290 5796 26292
rect 5740 26238 5742 26290
rect 5742 26238 5794 26290
rect 5794 26238 5796 26290
rect 5740 26236 5796 26238
rect 5740 25676 5796 25732
rect 4956 24892 5012 24948
rect 4620 24668 4676 24724
rect 4956 24722 5012 24724
rect 4956 24670 4958 24722
rect 4958 24670 5010 24722
rect 5010 24670 5012 24722
rect 4956 24668 5012 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2492 23660 2548 23716
rect 3612 23714 3668 23716
rect 3612 23662 3614 23714
rect 3614 23662 3666 23714
rect 3666 23662 3668 23714
rect 3612 23660 3668 23662
rect 3500 23324 3556 23380
rect 4732 23714 4788 23716
rect 4732 23662 4734 23714
rect 4734 23662 4786 23714
rect 4786 23662 4788 23714
rect 4732 23660 4788 23662
rect 4396 23100 4452 23156
rect 4620 23212 4676 23268
rect 5404 24946 5460 24948
rect 5404 24894 5406 24946
rect 5406 24894 5458 24946
rect 5458 24894 5460 24946
rect 5404 24892 5460 24894
rect 5404 24498 5460 24500
rect 5404 24446 5406 24498
rect 5406 24446 5458 24498
rect 5458 24446 5460 24498
rect 5404 24444 5460 24446
rect 5740 23714 5796 23716
rect 5740 23662 5742 23714
rect 5742 23662 5794 23714
rect 5794 23662 5796 23714
rect 5740 23660 5796 23662
rect 7644 31724 7700 31780
rect 6188 31500 6244 31556
rect 6300 31388 6356 31444
rect 6188 30210 6244 30212
rect 6188 30158 6190 30210
rect 6190 30158 6242 30210
rect 6242 30158 6244 30210
rect 6188 30156 6244 30158
rect 7196 31164 7252 31220
rect 7420 31666 7476 31668
rect 7420 31614 7422 31666
rect 7422 31614 7474 31666
rect 7474 31614 7476 31666
rect 7420 31612 7476 31614
rect 8428 31778 8484 31780
rect 8428 31726 8430 31778
rect 8430 31726 8482 31778
rect 8482 31726 8484 31778
rect 8428 31724 8484 31726
rect 7756 31388 7812 31444
rect 6972 30380 7028 30436
rect 7308 30380 7364 30436
rect 6748 30268 6804 30324
rect 6636 29986 6692 29988
rect 6636 29934 6638 29986
rect 6638 29934 6690 29986
rect 6690 29934 6692 29986
rect 6636 29932 6692 29934
rect 6524 29484 6580 29540
rect 7420 30322 7476 30324
rect 7420 30270 7422 30322
rect 7422 30270 7474 30322
rect 7474 30270 7476 30322
rect 7420 30268 7476 30270
rect 7868 31052 7924 31108
rect 7868 30268 7924 30324
rect 7084 30210 7140 30212
rect 7084 30158 7086 30210
rect 7086 30158 7138 30210
rect 7138 30158 7140 30210
rect 7084 30156 7140 30158
rect 6860 29596 6916 29652
rect 6636 28754 6692 28756
rect 6636 28702 6638 28754
rect 6638 28702 6690 28754
rect 6690 28702 6692 28754
rect 6636 28700 6692 28702
rect 7308 29426 7364 29428
rect 7308 29374 7310 29426
rect 7310 29374 7362 29426
rect 7362 29374 7364 29426
rect 7308 29372 7364 29374
rect 7420 28754 7476 28756
rect 7420 28702 7422 28754
rect 7422 28702 7474 28754
rect 7474 28702 7476 28754
rect 7420 28700 7476 28702
rect 6412 28140 6468 28196
rect 6188 27916 6244 27972
rect 8092 31164 8148 31220
rect 8428 31106 8484 31108
rect 8428 31054 8430 31106
rect 8430 31054 8482 31106
rect 8482 31054 8484 31106
rect 8428 31052 8484 31054
rect 8428 30380 8484 30436
rect 8092 30044 8148 30100
rect 7756 28140 7812 28196
rect 7644 27858 7700 27860
rect 7644 27806 7646 27858
rect 7646 27806 7698 27858
rect 7698 27806 7700 27858
rect 7644 27804 7700 27806
rect 6076 24332 6132 24388
rect 6188 24722 6244 24724
rect 6188 24670 6190 24722
rect 6190 24670 6242 24722
rect 6242 24670 6244 24722
rect 6188 24668 6244 24670
rect 6076 23884 6132 23940
rect 5516 23378 5572 23380
rect 5516 23326 5518 23378
rect 5518 23326 5570 23378
rect 5570 23326 5572 23378
rect 5516 23324 5572 23326
rect 2828 22316 2884 22372
rect 2716 21644 2772 21700
rect 2492 21474 2548 21476
rect 2492 21422 2494 21474
rect 2494 21422 2546 21474
rect 2546 21422 2548 21474
rect 2492 21420 2548 21422
rect 2044 20300 2100 20356
rect 2268 20578 2324 20580
rect 2268 20526 2270 20578
rect 2270 20526 2322 20578
rect 2322 20526 2324 20578
rect 2268 20524 2324 20526
rect 3052 20690 3108 20692
rect 3052 20638 3054 20690
rect 3054 20638 3106 20690
rect 3106 20638 3108 20690
rect 3052 20636 3108 20638
rect 3276 20300 3332 20356
rect 2604 20018 2660 20020
rect 2604 19966 2606 20018
rect 2606 19966 2658 20018
rect 2658 19966 2660 20018
rect 2604 19964 2660 19966
rect 1820 18508 1876 18564
rect 2492 19068 2548 19124
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4732 22482 4788 22484
rect 4732 22430 4734 22482
rect 4734 22430 4786 22482
rect 4786 22430 4788 22482
rect 4732 22428 4788 22430
rect 4396 22370 4452 22372
rect 4396 22318 4398 22370
rect 4398 22318 4450 22370
rect 4450 22318 4452 22370
rect 4396 22316 4452 22318
rect 4060 22204 4116 22260
rect 3948 22092 4004 22148
rect 3612 21420 3668 21476
rect 3500 20690 3556 20692
rect 3500 20638 3502 20690
rect 3502 20638 3554 20690
rect 3554 20638 3556 20690
rect 3500 20636 3556 20638
rect 5516 22146 5572 22148
rect 5516 22094 5518 22146
rect 5518 22094 5570 22146
rect 5570 22094 5572 22146
rect 5516 22092 5572 22094
rect 5292 21756 5348 21812
rect 4956 21698 5012 21700
rect 4956 21646 4958 21698
rect 4958 21646 5010 21698
rect 5010 21646 5012 21698
rect 4956 21644 5012 21646
rect 5740 23266 5796 23268
rect 5740 23214 5742 23266
rect 5742 23214 5794 23266
rect 5794 23214 5796 23266
rect 5740 23212 5796 23214
rect 5852 23154 5908 23156
rect 5852 23102 5854 23154
rect 5854 23102 5906 23154
rect 5906 23102 5908 23154
rect 5852 23100 5908 23102
rect 6524 25004 6580 25060
rect 6524 24834 6580 24836
rect 6524 24782 6526 24834
rect 6526 24782 6578 24834
rect 6578 24782 6580 24834
rect 6524 24780 6580 24782
rect 7196 25116 7252 25172
rect 7084 25004 7140 25060
rect 6412 23548 6468 23604
rect 7980 27858 8036 27860
rect 7980 27806 7982 27858
rect 7982 27806 8034 27858
rect 8034 27806 8036 27858
rect 7980 27804 8036 27806
rect 10108 38050 10164 38052
rect 10108 37998 10110 38050
rect 10110 37998 10162 38050
rect 10162 37998 10164 38050
rect 10108 37996 10164 37998
rect 11564 38220 11620 38276
rect 11900 38668 11956 38724
rect 13132 39116 13188 39172
rect 11900 37884 11956 37940
rect 10892 37660 10948 37716
rect 9884 37266 9940 37268
rect 9884 37214 9886 37266
rect 9886 37214 9938 37266
rect 9938 37214 9940 37266
rect 9884 37212 9940 37214
rect 9436 35644 9492 35700
rect 9772 35586 9828 35588
rect 9772 35534 9774 35586
rect 9774 35534 9826 35586
rect 9826 35534 9828 35586
rect 9772 35532 9828 35534
rect 10108 35196 10164 35252
rect 9884 35084 9940 35140
rect 9660 35026 9716 35028
rect 9660 34974 9662 35026
rect 9662 34974 9714 35026
rect 9714 34974 9716 35026
rect 9660 34972 9716 34974
rect 9884 34354 9940 34356
rect 9884 34302 9886 34354
rect 9886 34302 9938 34354
rect 9938 34302 9940 34354
rect 9884 34300 9940 34302
rect 9996 34748 10052 34804
rect 10332 34412 10388 34468
rect 10780 34412 10836 34468
rect 10444 34354 10500 34356
rect 10444 34302 10446 34354
rect 10446 34302 10498 34354
rect 10498 34302 10500 34354
rect 10444 34300 10500 34302
rect 9660 34188 9716 34244
rect 9996 33346 10052 33348
rect 9996 33294 9998 33346
rect 9998 33294 10050 33346
rect 10050 33294 10052 33346
rect 9996 33292 10052 33294
rect 9548 32284 9604 32340
rect 9548 31612 9604 31668
rect 11788 37266 11844 37268
rect 11788 37214 11790 37266
rect 11790 37214 11842 37266
rect 11842 37214 11844 37266
rect 11788 37212 11844 37214
rect 12348 37826 12404 37828
rect 12348 37774 12350 37826
rect 12350 37774 12402 37826
rect 12402 37774 12404 37826
rect 12348 37772 12404 37774
rect 13132 38220 13188 38276
rect 12796 37938 12852 37940
rect 12796 37886 12798 37938
rect 12798 37886 12850 37938
rect 12850 37886 12852 37938
rect 12796 37884 12852 37886
rect 12684 37660 12740 37716
rect 13692 37938 13748 37940
rect 13692 37886 13694 37938
rect 13694 37886 13746 37938
rect 13746 37886 13748 37938
rect 13692 37884 13748 37886
rect 12684 37212 12740 37268
rect 11452 37042 11508 37044
rect 11452 36990 11454 37042
rect 11454 36990 11506 37042
rect 11506 36990 11508 37042
rect 11452 36988 11508 36990
rect 11116 34354 11172 34356
rect 11116 34302 11118 34354
rect 11118 34302 11170 34354
rect 11170 34302 11172 34354
rect 11116 34300 11172 34302
rect 11788 34300 11844 34356
rect 11900 34524 11956 34580
rect 12012 34412 12068 34468
rect 11452 34242 11508 34244
rect 11452 34190 11454 34242
rect 11454 34190 11506 34242
rect 11506 34190 11508 34242
rect 11452 34188 11508 34190
rect 11676 34242 11732 34244
rect 11676 34190 11678 34242
rect 11678 34190 11730 34242
rect 11730 34190 11732 34242
rect 11676 34188 11732 34190
rect 11004 34018 11060 34020
rect 11004 33966 11006 34018
rect 11006 33966 11058 34018
rect 11058 33966 11060 34018
rect 11004 33964 11060 33966
rect 11900 34076 11956 34132
rect 11788 34018 11844 34020
rect 11788 33966 11790 34018
rect 11790 33966 11842 34018
rect 11842 33966 11844 34018
rect 11788 33964 11844 33966
rect 11788 33516 11844 33572
rect 11116 32562 11172 32564
rect 11116 32510 11118 32562
rect 11118 32510 11170 32562
rect 11170 32510 11172 32562
rect 11116 32508 11172 32510
rect 10332 32396 10388 32452
rect 10444 32338 10500 32340
rect 10444 32286 10446 32338
rect 10446 32286 10498 32338
rect 10498 32286 10500 32338
rect 10444 32284 10500 32286
rect 11788 32508 11844 32564
rect 12012 33852 12068 33908
rect 11900 33292 11956 33348
rect 11564 32396 11620 32452
rect 12348 37154 12404 37156
rect 12348 37102 12350 37154
rect 12350 37102 12402 37154
rect 12402 37102 12404 37154
rect 12348 37100 12404 37102
rect 13132 36988 13188 37044
rect 12572 36316 12628 36372
rect 12684 35532 12740 35588
rect 12572 34524 12628 34580
rect 12236 31948 12292 32004
rect 10220 31612 10276 31668
rect 9100 30994 9156 30996
rect 9100 30942 9102 30994
rect 9102 30942 9154 30994
rect 9154 30942 9156 30994
rect 9100 30940 9156 30942
rect 9884 30994 9940 30996
rect 9884 30942 9886 30994
rect 9886 30942 9938 30994
rect 9938 30942 9940 30994
rect 9884 30940 9940 30942
rect 11900 31500 11956 31556
rect 10668 30940 10724 30996
rect 10332 30268 10388 30324
rect 9548 30098 9604 30100
rect 9548 30046 9550 30098
rect 9550 30046 9602 30098
rect 9602 30046 9604 30098
rect 9548 30044 9604 30046
rect 8652 29650 8708 29652
rect 8652 29598 8654 29650
rect 8654 29598 8706 29650
rect 8706 29598 8708 29650
rect 8652 29596 8708 29598
rect 8876 29538 8932 29540
rect 8876 29486 8878 29538
rect 8878 29486 8930 29538
rect 8930 29486 8932 29538
rect 8876 29484 8932 29486
rect 8540 29372 8596 29428
rect 8988 29426 9044 29428
rect 8988 29374 8990 29426
rect 8990 29374 9042 29426
rect 9042 29374 9044 29426
rect 8988 29372 9044 29374
rect 8316 28588 8372 28644
rect 8764 28140 8820 28196
rect 8540 27858 8596 27860
rect 8540 27806 8542 27858
rect 8542 27806 8594 27858
rect 8594 27806 8596 27858
rect 8540 27804 8596 27806
rect 9548 28642 9604 28644
rect 9548 28590 9550 28642
rect 9550 28590 9602 28642
rect 9602 28590 9604 28642
rect 9548 28588 9604 28590
rect 10668 29986 10724 29988
rect 10668 29934 10670 29986
rect 10670 29934 10722 29986
rect 10722 29934 10724 29986
rect 10668 29932 10724 29934
rect 10444 28252 10500 28308
rect 9660 28140 9716 28196
rect 9212 26572 9268 26628
rect 9436 26236 9492 26292
rect 8316 25564 8372 25620
rect 7756 25228 7812 25284
rect 9660 26460 9716 26516
rect 10892 30940 10948 30996
rect 10892 30268 10948 30324
rect 12572 31388 12628 31444
rect 12460 29986 12516 29988
rect 12460 29934 12462 29986
rect 12462 29934 12514 29986
rect 12514 29934 12516 29986
rect 12460 29932 12516 29934
rect 11228 29484 11284 29540
rect 11116 28754 11172 28756
rect 11116 28702 11118 28754
rect 11118 28702 11170 28754
rect 11170 28702 11172 28754
rect 11116 28700 11172 28702
rect 11564 28700 11620 28756
rect 12236 28812 12292 28868
rect 10780 28642 10836 28644
rect 10780 28590 10782 28642
rect 10782 28590 10834 28642
rect 10834 28590 10836 28642
rect 10780 28588 10836 28590
rect 11676 28530 11732 28532
rect 11676 28478 11678 28530
rect 11678 28478 11730 28530
rect 11730 28478 11732 28530
rect 11676 28476 11732 28478
rect 11564 28418 11620 28420
rect 11564 28366 11566 28418
rect 11566 28366 11618 28418
rect 11618 28366 11620 28418
rect 11564 28364 11620 28366
rect 11004 28252 11060 28308
rect 11788 28252 11844 28308
rect 10668 26460 10724 26516
rect 11676 28140 11732 28196
rect 9436 25340 9492 25396
rect 8540 25228 8596 25284
rect 9772 25228 9828 25284
rect 10780 26290 10836 26292
rect 10780 26238 10782 26290
rect 10782 26238 10834 26290
rect 10834 26238 10836 26290
rect 10780 26236 10836 26238
rect 11004 25394 11060 25396
rect 11004 25342 11006 25394
rect 11006 25342 11058 25394
rect 11058 25342 11060 25394
rect 11004 25340 11060 25342
rect 7084 24108 7140 24164
rect 7756 24108 7812 24164
rect 6524 23660 6580 23716
rect 5740 22258 5796 22260
rect 5740 22206 5742 22258
rect 5742 22206 5794 22258
rect 5794 22206 5796 22258
rect 5740 22204 5796 22206
rect 5964 22876 6020 22932
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 3948 20524 4004 20580
rect 3052 19740 3108 19796
rect 2828 19292 2884 19348
rect 3500 19292 3556 19348
rect 3388 18508 3444 18564
rect 3836 18956 3892 19012
rect 4620 20300 4676 20356
rect 4620 19852 4676 19908
rect 4508 19740 4564 19796
rect 5852 21698 5908 21700
rect 5852 21646 5854 21698
rect 5854 21646 5906 21698
rect 5906 21646 5908 21698
rect 5852 21644 5908 21646
rect 5292 19740 5348 19796
rect 5516 19964 5572 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4732 19404 4788 19460
rect 4620 19346 4676 19348
rect 4620 19294 4622 19346
rect 4622 19294 4674 19346
rect 4674 19294 4676 19346
rect 4620 19292 4676 19294
rect 4284 19068 4340 19124
rect 5740 19292 5796 19348
rect 5852 18956 5908 19012
rect 5740 18844 5796 18900
rect 5292 18508 5348 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 6300 21756 6356 21812
rect 6300 20524 6356 20580
rect 6300 19964 6356 20020
rect 6076 19404 6132 19460
rect 6188 19852 6244 19908
rect 6188 18844 6244 18900
rect 5852 18508 5908 18564
rect 6636 23996 6692 24052
rect 7308 23826 7364 23828
rect 7308 23774 7310 23826
rect 7310 23774 7362 23826
rect 7362 23774 7364 23826
rect 7308 23772 7364 23774
rect 7084 23660 7140 23716
rect 6860 23154 6916 23156
rect 6860 23102 6862 23154
rect 6862 23102 6914 23154
rect 6914 23102 6916 23154
rect 6860 23100 6916 23102
rect 7084 22930 7140 22932
rect 7084 22878 7086 22930
rect 7086 22878 7138 22930
rect 7138 22878 7140 22930
rect 7084 22876 7140 22878
rect 7756 22428 7812 22484
rect 8540 24834 8596 24836
rect 8540 24782 8542 24834
rect 8542 24782 8594 24834
rect 8594 24782 8596 24834
rect 8540 24780 8596 24782
rect 8316 24722 8372 24724
rect 8316 24670 8318 24722
rect 8318 24670 8370 24722
rect 8370 24670 8372 24722
rect 8316 24668 8372 24670
rect 8092 23996 8148 24052
rect 7980 23938 8036 23940
rect 7980 23886 7982 23938
rect 7982 23886 8034 23938
rect 8034 23886 8036 23938
rect 7980 23884 8036 23886
rect 8204 23772 8260 23828
rect 7980 23660 8036 23716
rect 8652 24050 8708 24052
rect 8652 23998 8654 24050
rect 8654 23998 8706 24050
rect 8706 23998 8708 24050
rect 8652 23996 8708 23998
rect 8204 23154 8260 23156
rect 8204 23102 8206 23154
rect 8206 23102 8258 23154
rect 8258 23102 8260 23154
rect 8204 23100 8260 23102
rect 7084 21868 7140 21924
rect 6972 21810 7028 21812
rect 6972 21758 6974 21810
rect 6974 21758 7026 21810
rect 7026 21758 7028 21810
rect 6972 21756 7028 21758
rect 7868 21810 7924 21812
rect 7868 21758 7870 21810
rect 7870 21758 7922 21810
rect 7922 21758 7924 21810
rect 7868 21756 7924 21758
rect 8316 21868 8372 21924
rect 8428 23212 8484 23268
rect 8764 23100 8820 23156
rect 9772 24722 9828 24724
rect 9772 24670 9774 24722
rect 9774 24670 9826 24722
rect 9826 24670 9828 24722
rect 9772 24668 9828 24670
rect 9772 23772 9828 23828
rect 9884 23154 9940 23156
rect 9884 23102 9886 23154
rect 9886 23102 9938 23154
rect 9938 23102 9940 23154
rect 9884 23100 9940 23102
rect 11452 24108 11508 24164
rect 10780 23826 10836 23828
rect 10780 23774 10782 23826
rect 10782 23774 10834 23826
rect 10834 23774 10836 23826
rect 10780 23772 10836 23774
rect 10556 23266 10612 23268
rect 10556 23214 10558 23266
rect 10558 23214 10610 23266
rect 10610 23214 10612 23266
rect 10556 23212 10612 23214
rect 8764 22652 8820 22708
rect 9996 22370 10052 22372
rect 9996 22318 9998 22370
rect 9998 22318 10050 22370
rect 10050 22318 10052 22370
rect 9996 22316 10052 22318
rect 8540 21756 8596 21812
rect 8092 21586 8148 21588
rect 8092 21534 8094 21586
rect 8094 21534 8146 21586
rect 8146 21534 8148 21586
rect 8092 21532 8148 21534
rect 7756 20636 7812 20692
rect 8428 21420 8484 21476
rect 8092 20076 8148 20132
rect 8204 19852 8260 19908
rect 9772 21586 9828 21588
rect 9772 21534 9774 21586
rect 9774 21534 9826 21586
rect 9826 21534 9828 21586
rect 9772 21532 9828 21534
rect 10332 23154 10388 23156
rect 10332 23102 10334 23154
rect 10334 23102 10386 23154
rect 10386 23102 10388 23154
rect 10332 23100 10388 23102
rect 9436 20690 9492 20692
rect 9436 20638 9438 20690
rect 9438 20638 9490 20690
rect 9490 20638 9492 20690
rect 9436 20636 9492 20638
rect 8876 20130 8932 20132
rect 8876 20078 8878 20130
rect 8878 20078 8930 20130
rect 8930 20078 8932 20130
rect 8876 20076 8932 20078
rect 11452 22316 11508 22372
rect 10780 21756 10836 21812
rect 10668 20636 10724 20692
rect 10108 20076 10164 20132
rect 9772 19906 9828 19908
rect 9772 19854 9774 19906
rect 9774 19854 9826 19906
rect 9826 19854 9828 19906
rect 9772 19852 9828 19854
rect 8540 19740 8596 19796
rect 4620 16770 4676 16772
rect 4620 16718 4622 16770
rect 4622 16718 4674 16770
rect 4674 16718 4676 16770
rect 4620 16716 4676 16718
rect 5516 16770 5572 16772
rect 5516 16718 5518 16770
rect 5518 16718 5570 16770
rect 5570 16718 5572 16770
rect 5516 16716 5572 16718
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2492 16268 2548 16324
rect 4732 16322 4788 16324
rect 4732 16270 4734 16322
rect 4734 16270 4786 16322
rect 4786 16270 4788 16322
rect 4732 16268 4788 16270
rect 3500 15596 3556 15652
rect 3836 15596 3892 15652
rect 4732 15596 4788 15652
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4396 14530 4452 14532
rect 4396 14478 4398 14530
rect 4398 14478 4450 14530
rect 4450 14478 4452 14530
rect 4396 14476 4452 14478
rect 5628 15708 5684 15764
rect 6076 15314 6132 15316
rect 6076 15262 6078 15314
rect 6078 15262 6130 15314
rect 6130 15262 6132 15314
rect 6076 15260 6132 15262
rect 5852 14476 5908 14532
rect 5628 14418 5684 14420
rect 5628 14366 5630 14418
rect 5630 14366 5682 14418
rect 5682 14366 5684 14418
rect 5628 14364 5684 14366
rect 7756 19234 7812 19236
rect 7756 19182 7758 19234
rect 7758 19182 7810 19234
rect 7810 19182 7812 19234
rect 7756 19180 7812 19182
rect 8652 19234 8708 19236
rect 8652 19182 8654 19234
rect 8654 19182 8706 19234
rect 8706 19182 8708 19234
rect 8652 19180 8708 19182
rect 7532 18956 7588 19012
rect 8540 19010 8596 19012
rect 8540 18958 8542 19010
rect 8542 18958 8594 19010
rect 8594 18958 8596 19010
rect 8540 18956 8596 18958
rect 10332 20524 10388 20580
rect 9100 19010 9156 19012
rect 9100 18958 9102 19010
rect 9102 18958 9154 19010
rect 9154 18958 9156 19010
rect 9100 18956 9156 18958
rect 6860 16770 6916 16772
rect 6860 16718 6862 16770
rect 6862 16718 6914 16770
rect 6914 16718 6916 16770
rect 6860 16716 6916 16718
rect 6188 14028 6244 14084
rect 3612 13692 3668 13748
rect 2268 13580 2324 13636
rect 1820 8428 1876 8484
rect 1708 6636 1764 6692
rect 3052 13020 3108 13076
rect 3276 12850 3332 12852
rect 3276 12798 3278 12850
rect 3278 12798 3330 12850
rect 3330 12798 3332 12850
rect 3276 12796 3332 12798
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5180 13746 5236 13748
rect 5180 13694 5182 13746
rect 5182 13694 5234 13746
rect 5234 13694 5236 13746
rect 5180 13692 5236 13694
rect 4508 12962 4564 12964
rect 4508 12910 4510 12962
rect 4510 12910 4562 12962
rect 4562 12910 4564 12962
rect 4508 12908 4564 12910
rect 3724 12850 3780 12852
rect 3724 12798 3726 12850
rect 3726 12798 3778 12850
rect 3778 12798 3780 12850
rect 3724 12796 3780 12798
rect 4172 12572 4228 12628
rect 5740 13020 5796 13076
rect 5852 12962 5908 12964
rect 5852 12910 5854 12962
rect 5854 12910 5906 12962
rect 5906 12910 5908 12962
rect 5852 12908 5908 12910
rect 7084 15036 7140 15092
rect 9660 16882 9716 16884
rect 9660 16830 9662 16882
rect 9662 16830 9714 16882
rect 9714 16830 9716 16882
rect 9660 16828 9716 16830
rect 10108 17052 10164 17108
rect 8876 16098 8932 16100
rect 8876 16046 8878 16098
rect 8878 16046 8930 16098
rect 8930 16046 8932 16098
rect 8876 16044 8932 16046
rect 9548 16098 9604 16100
rect 9548 16046 9550 16098
rect 9550 16046 9602 16098
rect 9602 16046 9604 16098
rect 9548 16044 9604 16046
rect 9660 15986 9716 15988
rect 9660 15934 9662 15986
rect 9662 15934 9714 15986
rect 9714 15934 9716 15986
rect 9660 15932 9716 15934
rect 9212 15874 9268 15876
rect 9212 15822 9214 15874
rect 9214 15822 9266 15874
rect 9266 15822 9268 15874
rect 9212 15820 9268 15822
rect 10108 15820 10164 15876
rect 10780 18396 10836 18452
rect 11004 20578 11060 20580
rect 11004 20526 11006 20578
rect 11006 20526 11058 20578
rect 11058 20526 11060 20578
rect 11004 20524 11060 20526
rect 11228 19404 11284 19460
rect 10780 17052 10836 17108
rect 10556 16716 10612 16772
rect 10444 15986 10500 15988
rect 10444 15934 10446 15986
rect 10446 15934 10498 15986
rect 10498 15934 10500 15986
rect 10444 15932 10500 15934
rect 10668 15874 10724 15876
rect 10668 15822 10670 15874
rect 10670 15822 10722 15874
rect 10722 15822 10724 15874
rect 10668 15820 10724 15822
rect 8876 15260 8932 15316
rect 8988 15148 9044 15204
rect 10332 15314 10388 15316
rect 10332 15262 10334 15314
rect 10334 15262 10386 15314
rect 10386 15262 10388 15314
rect 10332 15260 10388 15262
rect 8092 14700 8148 14756
rect 7756 14642 7812 14644
rect 7756 14590 7758 14642
rect 7758 14590 7810 14642
rect 7810 14590 7812 14642
rect 7756 14588 7812 14590
rect 6748 13916 6804 13972
rect 6972 14364 7028 14420
rect 7084 14252 7140 14308
rect 8428 14252 8484 14308
rect 6636 13580 6692 13636
rect 6748 13468 6804 13524
rect 7308 13522 7364 13524
rect 7308 13470 7310 13522
rect 7310 13470 7362 13522
rect 7362 13470 7364 13522
rect 7308 13468 7364 13470
rect 8876 13970 8932 13972
rect 8876 13918 8878 13970
rect 8878 13918 8930 13970
rect 8930 13918 8932 13970
rect 8876 13916 8932 13918
rect 8764 13858 8820 13860
rect 8764 13806 8766 13858
rect 8766 13806 8818 13858
rect 8818 13806 8820 13858
rect 8764 13804 8820 13806
rect 10220 15202 10276 15204
rect 10220 15150 10222 15202
rect 10222 15150 10274 15202
rect 10274 15150 10276 15202
rect 10220 15148 10276 15150
rect 9884 14476 9940 14532
rect 9548 13970 9604 13972
rect 9548 13918 9550 13970
rect 9550 13918 9602 13970
rect 9602 13918 9604 13970
rect 9548 13916 9604 13918
rect 10220 14642 10276 14644
rect 10220 14590 10222 14642
rect 10222 14590 10274 14642
rect 10274 14590 10276 14642
rect 10220 14588 10276 14590
rect 10332 14418 10388 14420
rect 10332 14366 10334 14418
rect 10334 14366 10386 14418
rect 10386 14366 10388 14418
rect 10332 14364 10388 14366
rect 11116 16828 11172 16884
rect 10892 14530 10948 14532
rect 10892 14478 10894 14530
rect 10894 14478 10946 14530
rect 10946 14478 10948 14530
rect 10892 14476 10948 14478
rect 9772 13468 9828 13524
rect 5068 12738 5124 12740
rect 5068 12686 5070 12738
rect 5070 12686 5122 12738
rect 5122 12686 5124 12738
rect 5068 12684 5124 12686
rect 2492 10780 2548 10836
rect 2828 11116 2884 11172
rect 3276 8316 3332 8372
rect 3052 8092 3108 8148
rect 2492 6860 2548 6916
rect 2604 6748 2660 6804
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4844 11394 4900 11396
rect 4844 11342 4846 11394
rect 4846 11342 4898 11394
rect 4898 11342 4900 11394
rect 4844 11340 4900 11342
rect 4508 11282 4564 11284
rect 4508 11230 4510 11282
rect 4510 11230 4562 11282
rect 4562 11230 4564 11282
rect 4508 11228 4564 11230
rect 4620 11170 4676 11172
rect 4620 11118 4622 11170
rect 4622 11118 4674 11170
rect 4674 11118 4676 11170
rect 4620 11116 4676 11118
rect 6076 12572 6132 12628
rect 6524 12684 6580 12740
rect 5516 12290 5572 12292
rect 5516 12238 5518 12290
rect 5518 12238 5570 12290
rect 5570 12238 5572 12290
rect 5516 12236 5572 12238
rect 5740 12178 5796 12180
rect 5740 12126 5742 12178
rect 5742 12126 5794 12178
rect 5794 12126 5796 12178
rect 5740 12124 5796 12126
rect 5516 11228 5572 11284
rect 5292 10780 5348 10836
rect 5964 12124 6020 12180
rect 6188 11788 6244 11844
rect 5964 11340 6020 11396
rect 7532 12684 7588 12740
rect 7084 12236 7140 12292
rect 6636 12178 6692 12180
rect 6636 12126 6638 12178
rect 6638 12126 6690 12178
rect 6690 12126 6692 12178
rect 6636 12124 6692 12126
rect 6748 11788 6804 11844
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 9660 12402 9716 12404
rect 9660 12350 9662 12402
rect 9662 12350 9714 12402
rect 9714 12350 9716 12402
rect 9660 12348 9716 12350
rect 7980 10668 8036 10724
rect 8540 10722 8596 10724
rect 8540 10670 8542 10722
rect 8542 10670 8594 10722
rect 8594 10670 8596 10722
rect 8540 10668 8596 10670
rect 9436 10444 9492 10500
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 3612 8428 3668 8484
rect 7084 9826 7140 9828
rect 7084 9774 7086 9826
rect 7086 9774 7138 9826
rect 7138 9774 7140 9826
rect 7084 9772 7140 9774
rect 7532 9602 7588 9604
rect 7532 9550 7534 9602
rect 7534 9550 7586 9602
rect 7586 9550 7588 9602
rect 7532 9548 7588 9550
rect 7756 9436 7812 9492
rect 8428 9548 8484 9604
rect 7644 9100 7700 9156
rect 3500 8370 3556 8372
rect 3500 8318 3502 8370
rect 3502 8318 3554 8370
rect 3554 8318 3556 8370
rect 3500 8316 3556 8318
rect 3612 8204 3668 8260
rect 3500 7980 3556 8036
rect 6412 8876 6468 8932
rect 9100 8988 9156 9044
rect 8428 8540 8484 8596
rect 8876 8652 8932 8708
rect 3948 8092 4004 8148
rect 2940 7532 2996 7588
rect 3836 7362 3892 7364
rect 3836 7310 3838 7362
rect 3838 7310 3890 7362
rect 3890 7310 3892 7362
rect 3836 7308 3892 7310
rect 3276 6802 3332 6804
rect 3276 6750 3278 6802
rect 3278 6750 3330 6802
rect 3330 6750 3332 6802
rect 3276 6748 3332 6750
rect 4508 8204 4564 8260
rect 4284 8146 4340 8148
rect 4284 8094 4286 8146
rect 4286 8094 4338 8146
rect 4338 8094 4340 8146
rect 4284 8092 4340 8094
rect 4620 7980 4676 8036
rect 4956 7586 5012 7588
rect 4956 7534 4958 7586
rect 4958 7534 5010 7586
rect 5010 7534 5012 7586
rect 4956 7532 5012 7534
rect 4508 7474 4564 7476
rect 4508 7422 4510 7474
rect 4510 7422 4562 7474
rect 4562 7422 4564 7474
rect 4508 7420 4564 7422
rect 5068 7362 5124 7364
rect 5068 7310 5070 7362
rect 5070 7310 5122 7362
rect 5122 7310 5124 7362
rect 5068 7308 5124 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4060 6748 4116 6804
rect 4396 6748 4452 6804
rect 2828 6636 2884 6692
rect 3612 6690 3668 6692
rect 3612 6638 3614 6690
rect 3614 6638 3666 6690
rect 3666 6638 3668 6690
rect 3612 6636 3668 6638
rect 4172 6690 4228 6692
rect 4172 6638 4174 6690
rect 4174 6638 4226 6690
rect 4226 6638 4228 6690
rect 4172 6636 4228 6638
rect 4956 6802 5012 6804
rect 4956 6750 4958 6802
rect 4958 6750 5010 6802
rect 5010 6750 5012 6802
rect 4956 6748 5012 6750
rect 8988 8428 9044 8484
rect 5628 7474 5684 7476
rect 5628 7422 5630 7474
rect 5630 7422 5682 7474
rect 5682 7422 5684 7474
rect 5628 7420 5684 7422
rect 5740 6860 5796 6916
rect 5628 6802 5684 6804
rect 5628 6750 5630 6802
rect 5630 6750 5682 6802
rect 5682 6750 5684 6802
rect 5628 6748 5684 6750
rect 5068 6690 5124 6692
rect 5068 6638 5070 6690
rect 5070 6638 5122 6690
rect 5122 6638 5124 6690
rect 5068 6636 5124 6638
rect 6188 6130 6244 6132
rect 6188 6078 6190 6130
rect 6190 6078 6242 6130
rect 6242 6078 6244 6130
rect 6188 6076 6244 6078
rect 6636 6412 6692 6468
rect 4844 5628 4900 5684
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4172 5180 4228 5236
rect 5516 5682 5572 5684
rect 5516 5630 5518 5682
rect 5518 5630 5570 5682
rect 5570 5630 5572 5682
rect 5516 5628 5572 5630
rect 5964 5628 6020 5684
rect 4956 5516 5012 5572
rect 7084 6188 7140 6244
rect 7420 6466 7476 6468
rect 7420 6414 7422 6466
rect 7422 6414 7474 6466
rect 7474 6414 7476 6466
rect 7420 6412 7476 6414
rect 7196 6076 7252 6132
rect 6636 5516 6692 5572
rect 7084 5516 7140 5572
rect 6300 5180 6356 5236
rect 5180 5122 5236 5124
rect 5180 5070 5182 5122
rect 5182 5070 5234 5122
rect 5234 5070 5236 5122
rect 5180 5068 5236 5070
rect 6076 5122 6132 5124
rect 6076 5070 6078 5122
rect 6078 5070 6130 5122
rect 6130 5070 6132 5122
rect 6076 5068 6132 5070
rect 9436 9436 9492 9492
rect 10444 13970 10500 13972
rect 10444 13918 10446 13970
rect 10446 13918 10498 13970
rect 10498 13918 10500 13970
rect 10444 13916 10500 13918
rect 11228 16716 11284 16772
rect 11564 16940 11620 16996
rect 11228 16044 11284 16100
rect 11116 13916 11172 13972
rect 11452 13970 11508 13972
rect 11452 13918 11454 13970
rect 11454 13918 11506 13970
rect 11506 13918 11508 13970
rect 11452 13916 11508 13918
rect 11564 13858 11620 13860
rect 11564 13806 11566 13858
rect 11566 13806 11618 13858
rect 11618 13806 11620 13858
rect 11564 13804 11620 13806
rect 11116 13746 11172 13748
rect 11116 13694 11118 13746
rect 11118 13694 11170 13746
rect 11170 13694 11172 13746
rect 11116 13692 11172 13694
rect 10108 12402 10164 12404
rect 10108 12350 10110 12402
rect 10110 12350 10162 12402
rect 10162 12350 10164 12402
rect 10108 12348 10164 12350
rect 11340 12348 11396 12404
rect 9548 8988 9604 9044
rect 9660 8930 9716 8932
rect 9660 8878 9662 8930
rect 9662 8878 9714 8930
rect 9714 8878 9716 8930
rect 9660 8876 9716 8878
rect 9436 8540 9492 8596
rect 10892 10610 10948 10612
rect 10892 10558 10894 10610
rect 10894 10558 10946 10610
rect 10946 10558 10948 10610
rect 10892 10556 10948 10558
rect 11004 10498 11060 10500
rect 11004 10446 11006 10498
rect 11006 10446 11058 10498
rect 11058 10446 11060 10498
rect 11004 10444 11060 10446
rect 11452 9884 11508 9940
rect 11228 9266 11284 9268
rect 11228 9214 11230 9266
rect 11230 9214 11282 9266
rect 11282 9214 11284 9266
rect 11228 9212 11284 9214
rect 10108 9154 10164 9156
rect 10108 9102 10110 9154
rect 10110 9102 10162 9154
rect 10162 9102 10164 9154
rect 10108 9100 10164 9102
rect 11788 24220 11844 24276
rect 12124 28252 12180 28308
rect 12124 27580 12180 27636
rect 12460 27858 12516 27860
rect 12460 27806 12462 27858
rect 12462 27806 12514 27858
rect 12514 27806 12516 27858
rect 12460 27804 12516 27806
rect 13020 35308 13076 35364
rect 13020 34354 13076 34356
rect 13020 34302 13022 34354
rect 13022 34302 13074 34354
rect 13074 34302 13076 34354
rect 13020 34300 13076 34302
rect 12796 33964 12852 34020
rect 12908 33122 12964 33124
rect 12908 33070 12910 33122
rect 12910 33070 12962 33122
rect 12962 33070 12964 33122
rect 12908 33068 12964 33070
rect 13020 31388 13076 31444
rect 13020 28754 13076 28756
rect 13020 28702 13022 28754
rect 13022 28702 13074 28754
rect 13074 28702 13076 28754
rect 13020 28700 13076 28702
rect 14140 39618 14196 39620
rect 14140 39566 14142 39618
rect 14142 39566 14194 39618
rect 14194 39566 14196 39618
rect 14140 39564 14196 39566
rect 14028 39340 14084 39396
rect 13916 38108 13972 38164
rect 15148 43708 15204 43764
rect 18172 44380 18228 44436
rect 17500 44322 17556 44324
rect 17500 44270 17502 44322
rect 17502 44270 17554 44322
rect 17554 44270 17556 44322
rect 17500 44268 17556 44270
rect 14364 42700 14420 42756
rect 14364 39564 14420 39620
rect 14924 41804 14980 41860
rect 15148 42754 15204 42756
rect 15148 42702 15150 42754
rect 15150 42702 15202 42754
rect 15202 42702 15204 42754
rect 15148 42700 15204 42702
rect 14700 41244 14756 41300
rect 17948 43820 18004 43876
rect 15932 43372 15988 43428
rect 15820 42754 15876 42756
rect 15820 42702 15822 42754
rect 15822 42702 15874 42754
rect 15874 42702 15876 42754
rect 15820 42700 15876 42702
rect 15484 41580 15540 41636
rect 15036 40514 15092 40516
rect 15036 40462 15038 40514
rect 15038 40462 15090 40514
rect 15090 40462 15092 40514
rect 15036 40460 15092 40462
rect 15596 41186 15652 41188
rect 15596 41134 15598 41186
rect 15598 41134 15650 41186
rect 15650 41134 15652 41186
rect 15596 41132 15652 41134
rect 15708 40514 15764 40516
rect 15708 40462 15710 40514
rect 15710 40462 15762 40514
rect 15762 40462 15764 40514
rect 15708 40460 15764 40462
rect 16268 41692 16324 41748
rect 16156 41468 16212 41524
rect 16828 43426 16884 43428
rect 16828 43374 16830 43426
rect 16830 43374 16882 43426
rect 16882 43374 16884 43426
rect 16828 43372 16884 43374
rect 16828 42028 16884 42084
rect 17276 42364 17332 42420
rect 16492 41132 16548 41188
rect 15484 39618 15540 39620
rect 15484 39566 15486 39618
rect 15486 39566 15538 39618
rect 15538 39566 15540 39618
rect 15484 39564 15540 39566
rect 14588 39452 14644 39508
rect 14476 39394 14532 39396
rect 14476 39342 14478 39394
rect 14478 39342 14530 39394
rect 14530 39342 14532 39394
rect 14476 39340 14532 39342
rect 15260 39340 15316 39396
rect 14252 37884 14308 37940
rect 14364 38668 14420 38724
rect 15148 38722 15204 38724
rect 15148 38670 15150 38722
rect 15150 38670 15202 38722
rect 15202 38670 15204 38722
rect 15148 38668 15204 38670
rect 15596 38780 15652 38836
rect 13468 36316 13524 36372
rect 14588 36204 14644 36260
rect 14700 37996 14756 38052
rect 13692 35026 13748 35028
rect 13692 34974 13694 35026
rect 13694 34974 13746 35026
rect 13746 34974 13748 35026
rect 13692 34972 13748 34974
rect 13804 34412 13860 34468
rect 17500 42082 17556 42084
rect 17500 42030 17502 42082
rect 17502 42030 17554 42082
rect 17554 42030 17556 42082
rect 17500 42028 17556 42030
rect 17388 41580 17444 41636
rect 16604 39452 16660 39508
rect 16716 39340 16772 39396
rect 16940 39564 16996 39620
rect 16156 38610 16212 38612
rect 16156 38558 16158 38610
rect 16158 38558 16210 38610
rect 16210 38558 16212 38610
rect 16156 38556 16212 38558
rect 16492 38780 16548 38836
rect 16716 37772 16772 37828
rect 16380 37154 16436 37156
rect 16380 37102 16382 37154
rect 16382 37102 16434 37154
rect 16434 37102 16436 37154
rect 16380 37100 16436 37102
rect 15596 36092 15652 36148
rect 16380 35980 16436 36036
rect 15708 35698 15764 35700
rect 15708 35646 15710 35698
rect 15710 35646 15762 35698
rect 15762 35646 15764 35698
rect 15708 35644 15764 35646
rect 15932 35308 15988 35364
rect 14700 34300 14756 34356
rect 14924 34412 14980 34468
rect 13580 34188 13636 34244
rect 13356 34130 13412 34132
rect 13356 34078 13358 34130
rect 13358 34078 13410 34130
rect 13410 34078 13412 34130
rect 13356 34076 13412 34078
rect 13468 31666 13524 31668
rect 13468 31614 13470 31666
rect 13470 31614 13522 31666
rect 13522 31614 13524 31666
rect 13468 31612 13524 31614
rect 13692 34018 13748 34020
rect 13692 33966 13694 34018
rect 13694 33966 13746 34018
rect 13746 33966 13748 34018
rect 13692 33964 13748 33966
rect 13916 33852 13972 33908
rect 14476 33852 14532 33908
rect 14252 33234 14308 33236
rect 14252 33182 14254 33234
rect 14254 33182 14306 33234
rect 14306 33182 14308 33234
rect 14252 33180 14308 33182
rect 14028 33068 14084 33124
rect 13916 31836 13972 31892
rect 13804 31554 13860 31556
rect 13804 31502 13806 31554
rect 13806 31502 13858 31554
rect 13858 31502 13860 31554
rect 13804 31500 13860 31502
rect 14812 32562 14868 32564
rect 14812 32510 14814 32562
rect 14814 32510 14866 32562
rect 14866 32510 14868 32562
rect 14812 32508 14868 32510
rect 14588 31836 14644 31892
rect 14140 31388 14196 31444
rect 15260 33964 15316 34020
rect 18396 42700 18452 42756
rect 18172 42476 18228 42532
rect 18060 41970 18116 41972
rect 18060 41918 18062 41970
rect 18062 41918 18114 41970
rect 18114 41918 18116 41970
rect 18060 41916 18116 41918
rect 17836 41356 17892 41412
rect 18060 41692 18116 41748
rect 18060 41244 18116 41300
rect 18396 41580 18452 41636
rect 18172 41132 18228 41188
rect 18396 41356 18452 41412
rect 17500 40348 17556 40404
rect 17612 40460 17668 40516
rect 17724 40178 17780 40180
rect 17724 40126 17726 40178
rect 17726 40126 17778 40178
rect 17778 40126 17780 40178
rect 17724 40124 17780 40126
rect 18060 38892 18116 38948
rect 17724 38834 17780 38836
rect 17724 38782 17726 38834
rect 17726 38782 17778 38834
rect 17778 38782 17780 38834
rect 17724 38780 17780 38782
rect 17164 38444 17220 38500
rect 17948 37996 18004 38052
rect 17500 37772 17556 37828
rect 17724 37548 17780 37604
rect 16940 37266 16996 37268
rect 16940 37214 16942 37266
rect 16942 37214 16994 37266
rect 16994 37214 16996 37266
rect 16940 37212 16996 37214
rect 17052 36652 17108 36708
rect 17388 36482 17444 36484
rect 17388 36430 17390 36482
rect 17390 36430 17442 36482
rect 17442 36430 17444 36482
rect 17388 36428 17444 36430
rect 17612 36428 17668 36484
rect 17500 36316 17556 36372
rect 16828 36092 16884 36148
rect 16940 35980 16996 36036
rect 17164 35980 17220 36036
rect 17052 35868 17108 35924
rect 16828 35810 16884 35812
rect 16828 35758 16830 35810
rect 16830 35758 16882 35810
rect 16882 35758 16884 35810
rect 16828 35756 16884 35758
rect 16940 34972 16996 35028
rect 16604 34914 16660 34916
rect 16604 34862 16606 34914
rect 16606 34862 16658 34914
rect 16658 34862 16660 34914
rect 16604 34860 16660 34862
rect 16492 34412 16548 34468
rect 17052 34300 17108 34356
rect 15372 33180 15428 33236
rect 15260 31724 15316 31780
rect 15372 31948 15428 32004
rect 14812 31388 14868 31444
rect 14588 31276 14644 31332
rect 13356 30994 13412 30996
rect 13356 30942 13358 30994
rect 13358 30942 13410 30994
rect 13410 30942 13412 30994
rect 13356 30940 13412 30942
rect 14028 30994 14084 30996
rect 14028 30942 14030 30994
rect 14030 30942 14082 30994
rect 14082 30942 14084 30994
rect 14028 30940 14084 30942
rect 13468 28418 13524 28420
rect 13468 28366 13470 28418
rect 13470 28366 13522 28418
rect 13522 28366 13524 28418
rect 13468 28364 13524 28366
rect 13580 27858 13636 27860
rect 13580 27806 13582 27858
rect 13582 27806 13634 27858
rect 13634 27806 13636 27858
rect 13580 27804 13636 27806
rect 13356 27692 13412 27748
rect 13244 27132 13300 27188
rect 14700 31106 14756 31108
rect 14700 31054 14702 31106
rect 14702 31054 14754 31106
rect 14754 31054 14756 31106
rect 14700 31052 14756 31054
rect 15260 30156 15316 30212
rect 14476 29260 14532 29316
rect 15260 29148 15316 29204
rect 14476 28700 14532 28756
rect 14700 27970 14756 27972
rect 14700 27918 14702 27970
rect 14702 27918 14754 27970
rect 14754 27918 14756 27970
rect 14700 27916 14756 27918
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 13916 27186 13972 27188
rect 13916 27134 13918 27186
rect 13918 27134 13970 27186
rect 13970 27134 13972 27186
rect 13916 27132 13972 27134
rect 13580 27020 13636 27076
rect 12796 25618 12852 25620
rect 12796 25566 12798 25618
rect 12798 25566 12850 25618
rect 12850 25566 12852 25618
rect 12796 25564 12852 25566
rect 12684 24556 12740 24612
rect 12348 24162 12404 24164
rect 12348 24110 12350 24162
rect 12350 24110 12402 24162
rect 12402 24110 12404 24162
rect 12348 24108 12404 24110
rect 12012 23826 12068 23828
rect 12012 23774 12014 23826
rect 12014 23774 12066 23826
rect 12066 23774 12068 23826
rect 12012 23772 12068 23774
rect 12460 23772 12516 23828
rect 14476 27692 14532 27748
rect 14252 27074 14308 27076
rect 14252 27022 14254 27074
rect 14254 27022 14306 27074
rect 14306 27022 14308 27074
rect 14252 27020 14308 27022
rect 13916 26290 13972 26292
rect 13916 26238 13918 26290
rect 13918 26238 13970 26290
rect 13970 26238 13972 26290
rect 13916 26236 13972 26238
rect 14252 25228 14308 25284
rect 13580 24668 13636 24724
rect 14588 27580 14644 27636
rect 15036 27132 15092 27188
rect 14700 26178 14756 26180
rect 14700 26126 14702 26178
rect 14702 26126 14754 26178
rect 14754 26126 14756 26178
rect 14700 26124 14756 26126
rect 15484 31388 15540 31444
rect 15708 31052 15764 31108
rect 15820 29596 15876 29652
rect 15820 29314 15876 29316
rect 15820 29262 15822 29314
rect 15822 29262 15874 29314
rect 15874 29262 15876 29314
rect 15820 29260 15876 29262
rect 15484 29148 15540 29204
rect 15484 27804 15540 27860
rect 17276 35868 17332 35924
rect 17388 35980 17444 36036
rect 17276 34690 17332 34692
rect 17276 34638 17278 34690
rect 17278 34638 17330 34690
rect 17330 34638 17332 34690
rect 17276 34636 17332 34638
rect 17836 36092 17892 36148
rect 17948 35980 18004 36036
rect 18284 39004 18340 39060
rect 18396 38668 18452 38724
rect 18172 38220 18228 38276
rect 17948 35756 18004 35812
rect 17724 35420 17780 35476
rect 17612 35308 17668 35364
rect 20412 44380 20468 44436
rect 20188 44210 20244 44212
rect 20188 44158 20190 44210
rect 20190 44158 20242 44210
rect 20242 44158 20244 44210
rect 20188 44156 20244 44158
rect 19852 44098 19908 44100
rect 19852 44046 19854 44098
rect 19854 44046 19906 44098
rect 19906 44046 19908 44098
rect 19852 44044 19908 44046
rect 21980 44380 22036 44436
rect 21756 44322 21812 44324
rect 21756 44270 21758 44322
rect 21758 44270 21810 44322
rect 21810 44270 21812 44322
rect 21756 44268 21812 44270
rect 20412 44044 20468 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19292 43708 19348 43764
rect 19180 43372 19236 43428
rect 19180 42364 19236 42420
rect 18956 39788 19012 39844
rect 18732 39564 18788 39620
rect 18620 38780 18676 38836
rect 18508 37154 18564 37156
rect 18508 37102 18510 37154
rect 18510 37102 18562 37154
rect 18562 37102 18564 37154
rect 18508 37100 18564 37102
rect 19292 41692 19348 41748
rect 20076 42978 20132 42980
rect 20076 42926 20078 42978
rect 20078 42926 20130 42978
rect 20130 42926 20132 42978
rect 20076 42924 20132 42926
rect 20860 44098 20916 44100
rect 20860 44046 20862 44098
rect 20862 44046 20914 44098
rect 20914 44046 20916 44098
rect 20860 44044 20916 44046
rect 21868 44210 21924 44212
rect 21868 44158 21870 44210
rect 21870 44158 21922 44210
rect 21922 44158 21924 44210
rect 21868 44156 21924 44158
rect 22428 44268 22484 44324
rect 22092 44098 22148 44100
rect 22092 44046 22094 44098
rect 22094 44046 22146 44098
rect 22146 44046 22148 44098
rect 22092 44044 22148 44046
rect 21980 43820 22036 43876
rect 21084 43596 21140 43652
rect 22764 44322 22820 44324
rect 22764 44270 22766 44322
rect 22766 44270 22818 44322
rect 22818 44270 22820 44322
rect 22764 44268 22820 44270
rect 22428 43708 22484 43764
rect 21644 43426 21700 43428
rect 21644 43374 21646 43426
rect 21646 43374 21698 43426
rect 21698 43374 21700 43426
rect 21644 43372 21700 43374
rect 22652 43932 22708 43988
rect 23100 44098 23156 44100
rect 23100 44046 23102 44098
rect 23102 44046 23154 44098
rect 23154 44046 23156 44098
rect 23100 44044 23156 44046
rect 22540 43372 22596 43428
rect 21868 42924 21924 42980
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19292 40236 19348 40292
rect 19292 39116 19348 39172
rect 20412 41186 20468 41188
rect 20412 41134 20414 41186
rect 20414 41134 20466 41186
rect 20466 41134 20468 41186
rect 20412 41132 20468 41134
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20188 40460 20244 40516
rect 20076 39788 20132 39844
rect 20524 39618 20580 39620
rect 20524 39566 20526 39618
rect 20526 39566 20578 39618
rect 20578 39566 20580 39618
rect 20524 39564 20580 39566
rect 19404 38892 19460 38948
rect 19404 38220 19460 38276
rect 19068 38050 19124 38052
rect 19068 37998 19070 38050
rect 19070 37998 19122 38050
rect 19122 37998 19124 38050
rect 19068 37996 19124 37998
rect 19180 36876 19236 36932
rect 18284 36482 18340 36484
rect 18284 36430 18286 36482
rect 18286 36430 18338 36482
rect 18338 36430 18340 36482
rect 18284 36428 18340 36430
rect 18396 36370 18452 36372
rect 18396 36318 18398 36370
rect 18398 36318 18450 36370
rect 18450 36318 18452 36370
rect 18396 36316 18452 36318
rect 18396 35756 18452 35812
rect 18060 35196 18116 35252
rect 17836 35026 17892 35028
rect 17836 34974 17838 35026
rect 17838 34974 17890 35026
rect 17890 34974 17892 35026
rect 17836 34972 17892 34974
rect 19180 36370 19236 36372
rect 19180 36318 19182 36370
rect 19182 36318 19234 36370
rect 19234 36318 19236 36370
rect 19180 36316 19236 36318
rect 18508 34636 18564 34692
rect 19068 34636 19124 34692
rect 18956 34300 19012 34356
rect 18620 34188 18676 34244
rect 16940 33516 16996 33572
rect 16828 32732 16884 32788
rect 16716 32620 16772 32676
rect 16268 32396 16324 32452
rect 16604 32562 16660 32564
rect 16604 32510 16606 32562
rect 16606 32510 16658 32562
rect 16658 32510 16660 32562
rect 16604 32508 16660 32510
rect 16380 32060 16436 32116
rect 16940 32060 16996 32116
rect 17052 33628 17108 33684
rect 16268 31948 16324 32004
rect 17500 33628 17556 33684
rect 17500 33458 17556 33460
rect 17500 33406 17502 33458
rect 17502 33406 17554 33458
rect 17554 33406 17556 33458
rect 17500 33404 17556 33406
rect 17948 33404 18004 33460
rect 18172 33628 18228 33684
rect 17500 33068 17556 33124
rect 17388 32674 17444 32676
rect 17388 32622 17390 32674
rect 17390 32622 17442 32674
rect 17442 32622 17444 32674
rect 17388 32620 17444 32622
rect 17948 32396 18004 32452
rect 17276 31778 17332 31780
rect 17276 31726 17278 31778
rect 17278 31726 17330 31778
rect 17330 31726 17332 31778
rect 17276 31724 17332 31726
rect 16380 30156 16436 30212
rect 17836 31554 17892 31556
rect 17836 31502 17838 31554
rect 17838 31502 17890 31554
rect 17890 31502 17892 31554
rect 17836 31500 17892 31502
rect 17388 30492 17444 30548
rect 17612 30156 17668 30212
rect 16380 29708 16436 29764
rect 17948 29932 18004 29988
rect 17836 29708 17892 29764
rect 17724 29650 17780 29652
rect 17724 29598 17726 29650
rect 17726 29598 17778 29650
rect 17778 29598 17780 29650
rect 17724 29596 17780 29598
rect 18060 32060 18116 32116
rect 16940 28588 16996 28644
rect 17164 29260 17220 29316
rect 15932 27356 15988 27412
rect 16268 27580 16324 27636
rect 14700 24610 14756 24612
rect 14700 24558 14702 24610
rect 14702 24558 14754 24610
rect 14754 24558 14756 24610
rect 14700 24556 14756 24558
rect 14812 24220 14868 24276
rect 12908 23938 12964 23940
rect 12908 23886 12910 23938
rect 12910 23886 12962 23938
rect 12962 23886 12964 23938
rect 12908 23884 12964 23886
rect 13244 23884 13300 23940
rect 13020 23324 13076 23380
rect 13580 23660 13636 23716
rect 12908 22482 12964 22484
rect 12908 22430 12910 22482
rect 12910 22430 12962 22482
rect 12962 22430 12964 22482
rect 12908 22428 12964 22430
rect 12796 22092 12852 22148
rect 13244 21756 13300 21812
rect 13804 23938 13860 23940
rect 13804 23886 13806 23938
rect 13806 23886 13858 23938
rect 13858 23886 13860 23938
rect 13804 23884 13860 23886
rect 13692 23324 13748 23380
rect 14140 23548 14196 23604
rect 13692 22428 13748 22484
rect 14028 22204 14084 22260
rect 13804 22146 13860 22148
rect 13804 22094 13806 22146
rect 13806 22094 13858 22146
rect 13858 22094 13860 22146
rect 13804 22092 13860 22094
rect 14140 21868 14196 21924
rect 12908 20972 12964 21028
rect 12684 20802 12740 20804
rect 12684 20750 12686 20802
rect 12686 20750 12738 20802
rect 12738 20750 12740 20802
rect 12684 20748 12740 20750
rect 11788 20578 11844 20580
rect 11788 20526 11790 20578
rect 11790 20526 11842 20578
rect 11842 20526 11844 20578
rect 11788 20524 11844 20526
rect 12012 19292 12068 19348
rect 13020 19852 13076 19908
rect 12236 19180 12292 19236
rect 11900 18396 11956 18452
rect 12908 19068 12964 19124
rect 13020 18508 13076 18564
rect 12572 17612 12628 17668
rect 12796 16994 12852 16996
rect 12796 16942 12798 16994
rect 12798 16942 12850 16994
rect 12850 16942 12852 16994
rect 12796 16940 12852 16942
rect 12908 16770 12964 16772
rect 12908 16718 12910 16770
rect 12910 16718 12962 16770
rect 12962 16718 12964 16770
rect 12908 16716 12964 16718
rect 14924 23714 14980 23716
rect 14924 23662 14926 23714
rect 14926 23662 14978 23714
rect 14978 23662 14980 23714
rect 14924 23660 14980 23662
rect 14700 23266 14756 23268
rect 14700 23214 14702 23266
rect 14702 23214 14754 23266
rect 14754 23214 14756 23266
rect 14700 23212 14756 23214
rect 14812 21868 14868 21924
rect 14252 20972 14308 21028
rect 13356 20748 13412 20804
rect 14028 20802 14084 20804
rect 14028 20750 14030 20802
rect 14030 20750 14082 20802
rect 14082 20750 14084 20802
rect 14028 20748 14084 20750
rect 13580 19404 13636 19460
rect 13804 19346 13860 19348
rect 13804 19294 13806 19346
rect 13806 19294 13858 19346
rect 13858 19294 13860 19346
rect 13804 19292 13860 19294
rect 14140 19180 14196 19236
rect 15372 20748 15428 20804
rect 15260 20130 15316 20132
rect 15260 20078 15262 20130
rect 15262 20078 15314 20130
rect 15314 20078 15316 20130
rect 15260 20076 15316 20078
rect 14476 19068 14532 19124
rect 14140 18396 14196 18452
rect 13244 17106 13300 17108
rect 13244 17054 13246 17106
rect 13246 17054 13298 17106
rect 13298 17054 13300 17106
rect 13244 17052 13300 17054
rect 14476 18060 14532 18116
rect 14252 17666 14308 17668
rect 14252 17614 14254 17666
rect 14254 17614 14306 17666
rect 14306 17614 14308 17666
rect 14252 17612 14308 17614
rect 16940 28364 16996 28420
rect 16828 27468 16884 27524
rect 16828 26236 16884 26292
rect 16380 25564 16436 25620
rect 16492 25340 16548 25396
rect 16828 25228 16884 25284
rect 16380 24722 16436 24724
rect 16380 24670 16382 24722
rect 16382 24670 16434 24722
rect 16434 24670 16436 24722
rect 16380 24668 16436 24670
rect 15708 24556 15764 24612
rect 15708 23548 15764 23604
rect 16156 23772 16212 23828
rect 15932 21810 15988 21812
rect 15932 21758 15934 21810
rect 15934 21758 15986 21810
rect 15986 21758 15988 21810
rect 15932 21756 15988 21758
rect 15708 20972 15764 21028
rect 16828 23100 16884 23156
rect 16380 22988 16436 23044
rect 16380 22652 16436 22708
rect 16268 22258 16324 22260
rect 16268 22206 16270 22258
rect 16270 22206 16322 22258
rect 16322 22206 16324 22258
rect 16268 22204 16324 22206
rect 16716 21196 16772 21252
rect 15484 19068 15540 19124
rect 15372 18450 15428 18452
rect 15372 18398 15374 18450
rect 15374 18398 15426 18450
rect 15426 18398 15428 18450
rect 15372 18396 15428 18398
rect 15260 18060 15316 18116
rect 15036 17612 15092 17668
rect 16268 18508 16324 18564
rect 16492 20524 16548 20580
rect 16716 20300 16772 20356
rect 16716 19852 16772 19908
rect 15932 18338 15988 18340
rect 15932 18286 15934 18338
rect 15934 18286 15986 18338
rect 15986 18286 15988 18338
rect 15932 18284 15988 18286
rect 15932 17724 15988 17780
rect 16044 17052 16100 17108
rect 15596 16940 15652 16996
rect 14588 16716 14644 16772
rect 14364 16268 14420 16324
rect 15036 16604 15092 16660
rect 15596 16322 15652 16324
rect 15596 16270 15598 16322
rect 15598 16270 15650 16322
rect 15650 16270 15652 16322
rect 15596 16268 15652 16270
rect 15260 15986 15316 15988
rect 15260 15934 15262 15986
rect 15262 15934 15314 15986
rect 15314 15934 15316 15986
rect 15260 15932 15316 15934
rect 15932 16716 15988 16772
rect 16156 16604 16212 16660
rect 16492 16716 16548 16772
rect 16380 15986 16436 15988
rect 16380 15934 16382 15986
rect 16382 15934 16434 15986
rect 16434 15934 16436 15986
rect 16380 15932 16436 15934
rect 15036 15708 15092 15764
rect 13132 14812 13188 14868
rect 11788 14364 11844 14420
rect 12236 14530 12292 14532
rect 12236 14478 12238 14530
rect 12238 14478 12290 14530
rect 12290 14478 12292 14530
rect 12236 14476 12292 14478
rect 12460 14418 12516 14420
rect 12460 14366 12462 14418
rect 12462 14366 12514 14418
rect 12514 14366 12516 14418
rect 12460 14364 12516 14366
rect 12124 13916 12180 13972
rect 12572 14252 12628 14308
rect 12012 13580 12068 13636
rect 12236 12348 12292 12404
rect 11788 10556 11844 10612
rect 12684 10556 12740 10612
rect 12348 10444 12404 10500
rect 12012 9938 12068 9940
rect 12012 9886 12014 9938
rect 12014 9886 12066 9938
rect 12066 9886 12068 9938
rect 12012 9884 12068 9886
rect 11900 9826 11956 9828
rect 11900 9774 11902 9826
rect 11902 9774 11954 9826
rect 11954 9774 11956 9826
rect 11900 9772 11956 9774
rect 12236 9772 12292 9828
rect 11788 9212 11844 9268
rect 11340 9154 11396 9156
rect 11340 9102 11342 9154
rect 11342 9102 11394 9154
rect 11394 9102 11396 9154
rect 11340 9100 11396 9102
rect 9884 8876 9940 8932
rect 9884 8652 9940 8708
rect 10108 8428 10164 8484
rect 8204 6690 8260 6692
rect 8204 6638 8206 6690
rect 8206 6638 8258 6690
rect 8258 6638 8260 6690
rect 8204 6636 8260 6638
rect 8204 6412 8260 6468
rect 7868 5964 7924 6020
rect 8316 6188 8372 6244
rect 7308 5180 7364 5236
rect 8764 6300 8820 6356
rect 8540 5234 8596 5236
rect 8540 5182 8542 5234
rect 8542 5182 8594 5234
rect 8594 5182 8596 5234
rect 8540 5180 8596 5182
rect 7756 4956 7812 5012
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 8652 4562 8708 4564
rect 8652 4510 8654 4562
rect 8654 4510 8706 4562
rect 8706 4510 8708 4562
rect 8652 4508 8708 4510
rect 6300 4226 6356 4228
rect 6300 4174 6302 4226
rect 6302 4174 6354 4226
rect 6354 4174 6356 4226
rect 6300 4172 6356 4174
rect 7532 4226 7588 4228
rect 7532 4174 7534 4226
rect 7534 4174 7586 4226
rect 7586 4174 7588 4226
rect 7532 4172 7588 4174
rect 9100 6188 9156 6244
rect 9100 6018 9156 6020
rect 9100 5966 9102 6018
rect 9102 5966 9154 6018
rect 9154 5966 9156 6018
rect 9100 5964 9156 5966
rect 9100 5628 9156 5684
rect 9436 6524 9492 6580
rect 8764 4284 8820 4340
rect 9548 6300 9604 6356
rect 10668 8316 10724 8372
rect 11788 8876 11844 8932
rect 12348 9714 12404 9716
rect 12348 9662 12350 9714
rect 12350 9662 12402 9714
rect 12402 9662 12404 9714
rect 12348 9660 12404 9662
rect 12684 9042 12740 9044
rect 12684 8990 12686 9042
rect 12686 8990 12738 9042
rect 12738 8990 12740 9042
rect 12684 8988 12740 8990
rect 11676 8316 11732 8372
rect 11452 8258 11508 8260
rect 11452 8206 11454 8258
rect 11454 8206 11506 8258
rect 11506 8206 11508 8258
rect 11452 8204 11508 8206
rect 11004 7420 11060 7476
rect 10780 6748 10836 6804
rect 9660 5740 9716 5796
rect 9548 5234 9604 5236
rect 9548 5182 9550 5234
rect 9550 5182 9602 5234
rect 9602 5182 9604 5234
rect 9548 5180 9604 5182
rect 12124 8204 12180 8260
rect 11676 7308 11732 7364
rect 12684 7980 12740 8036
rect 12236 6914 12292 6916
rect 12236 6862 12238 6914
rect 12238 6862 12290 6914
rect 12290 6862 12292 6914
rect 12236 6860 12292 6862
rect 12572 6802 12628 6804
rect 12572 6750 12574 6802
rect 12574 6750 12626 6802
rect 12626 6750 12628 6802
rect 12572 6748 12628 6750
rect 12012 6636 12068 6692
rect 11004 6412 11060 6468
rect 8988 4898 9044 4900
rect 8988 4846 8990 4898
rect 8990 4846 9042 4898
rect 9042 4846 9044 4898
rect 8988 4844 9044 4846
rect 10108 5122 10164 5124
rect 10108 5070 10110 5122
rect 10110 5070 10162 5122
rect 10162 5070 10164 5122
rect 10108 5068 10164 5070
rect 9660 4450 9716 4452
rect 9660 4398 9662 4450
rect 9662 4398 9714 4450
rect 9714 4398 9716 4450
rect 9660 4396 9716 4398
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 9772 4284 9828 4340
rect 8764 3778 8820 3780
rect 8764 3726 8766 3778
rect 8766 3726 8818 3778
rect 8818 3726 8820 3778
rect 8764 3724 8820 3726
rect 10556 4844 10612 4900
rect 8652 3442 8708 3444
rect 8652 3390 8654 3442
rect 8654 3390 8706 3442
rect 8706 3390 8708 3442
rect 8652 3388 8708 3390
rect 10444 3442 10500 3444
rect 10444 3390 10446 3442
rect 10446 3390 10498 3442
rect 10498 3390 10500 3442
rect 10444 3388 10500 3390
rect 12124 6466 12180 6468
rect 12124 6414 12126 6466
rect 12126 6414 12178 6466
rect 12178 6414 12180 6466
rect 12124 6412 12180 6414
rect 13020 14642 13076 14644
rect 13020 14590 13022 14642
rect 13022 14590 13074 14642
rect 13074 14590 13076 14642
rect 13020 14588 13076 14590
rect 13692 14530 13748 14532
rect 13692 14478 13694 14530
rect 13694 14478 13746 14530
rect 13746 14478 13748 14530
rect 13692 14476 13748 14478
rect 14140 15036 14196 15092
rect 14140 14588 14196 14644
rect 14924 15260 14980 15316
rect 13580 14418 13636 14420
rect 13580 14366 13582 14418
rect 13582 14366 13634 14418
rect 13634 14366 13636 14418
rect 13580 14364 13636 14366
rect 13468 14306 13524 14308
rect 13468 14254 13470 14306
rect 13470 14254 13522 14306
rect 13522 14254 13524 14306
rect 13468 14252 13524 14254
rect 14028 14028 14084 14084
rect 13132 13858 13188 13860
rect 13132 13806 13134 13858
rect 13134 13806 13186 13858
rect 13186 13806 13188 13858
rect 13132 13804 13188 13806
rect 15260 15314 15316 15316
rect 15260 15262 15262 15314
rect 15262 15262 15314 15314
rect 15314 15262 15316 15314
rect 15260 15260 15316 15262
rect 16268 15148 16324 15204
rect 16828 16770 16884 16772
rect 16828 16718 16830 16770
rect 16830 16718 16882 16770
rect 16882 16718 16884 16770
rect 16828 16716 16884 16718
rect 17948 28700 18004 28756
rect 17836 27970 17892 27972
rect 17836 27918 17838 27970
rect 17838 27918 17890 27970
rect 17890 27918 17892 27970
rect 17836 27916 17892 27918
rect 17500 27746 17556 27748
rect 17500 27694 17502 27746
rect 17502 27694 17554 27746
rect 17554 27694 17556 27746
rect 17500 27692 17556 27694
rect 17388 27634 17444 27636
rect 17388 27582 17390 27634
rect 17390 27582 17442 27634
rect 17442 27582 17444 27634
rect 17388 27580 17444 27582
rect 18396 32562 18452 32564
rect 18396 32510 18398 32562
rect 18398 32510 18450 32562
rect 18450 32510 18452 32562
rect 18396 32508 18452 32510
rect 18620 33404 18676 33460
rect 19068 32508 19124 32564
rect 18172 31276 18228 31332
rect 18172 30268 18228 30324
rect 20188 39340 20244 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20076 38780 20132 38836
rect 20300 39004 20356 39060
rect 20412 38668 20468 38724
rect 19628 37996 19684 38052
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19516 36370 19572 36372
rect 19516 36318 19518 36370
rect 19518 36318 19570 36370
rect 19570 36318 19572 36370
rect 19516 36316 19572 36318
rect 19404 35644 19460 35700
rect 19516 34412 19572 34468
rect 19404 33516 19460 33572
rect 20300 38220 20356 38276
rect 20300 37212 20356 37268
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19964 34802 20020 34804
rect 19964 34750 19966 34802
rect 19966 34750 20018 34802
rect 20018 34750 20020 34802
rect 19964 34748 20020 34750
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19964 34018 20020 34020
rect 19964 33966 19966 34018
rect 19966 33966 20018 34018
rect 20018 33966 20020 34018
rect 19964 33964 20020 33966
rect 19628 33458 19684 33460
rect 19628 33406 19630 33458
rect 19630 33406 19682 33458
rect 19682 33406 19684 33458
rect 19628 33404 19684 33406
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19740 32732 19796 32788
rect 20412 36258 20468 36260
rect 20412 36206 20414 36258
rect 20414 36206 20466 36258
rect 20466 36206 20468 36258
rect 20412 36204 20468 36206
rect 20412 35196 20468 35252
rect 21420 41020 21476 41076
rect 20860 40962 20916 40964
rect 20860 40910 20862 40962
rect 20862 40910 20914 40962
rect 20914 40910 20916 40962
rect 20860 40908 20916 40910
rect 21308 39506 21364 39508
rect 21308 39454 21310 39506
rect 21310 39454 21362 39506
rect 21362 39454 21364 39506
rect 21308 39452 21364 39454
rect 21644 40572 21700 40628
rect 21980 42700 22036 42756
rect 22876 40908 22932 40964
rect 23212 43708 23268 43764
rect 22988 40796 23044 40852
rect 23212 42700 23268 42756
rect 22876 40684 22932 40740
rect 21532 39004 21588 39060
rect 20860 38834 20916 38836
rect 20860 38782 20862 38834
rect 20862 38782 20914 38834
rect 20914 38782 20916 38834
rect 20860 38780 20916 38782
rect 21308 38834 21364 38836
rect 21308 38782 21310 38834
rect 21310 38782 21362 38834
rect 21362 38782 21364 38834
rect 21308 38780 21364 38782
rect 20748 38220 20804 38276
rect 20636 37212 20692 37268
rect 21756 38274 21812 38276
rect 21756 38222 21758 38274
rect 21758 38222 21810 38274
rect 21810 38222 21812 38274
rect 21756 38220 21812 38222
rect 21308 38050 21364 38052
rect 21308 37998 21310 38050
rect 21310 37998 21362 38050
rect 21362 37998 21364 38050
rect 21308 37996 21364 37998
rect 22204 37996 22260 38052
rect 20524 34972 20580 35028
rect 20636 34914 20692 34916
rect 20636 34862 20638 34914
rect 20638 34862 20690 34914
rect 20690 34862 20692 34914
rect 20636 34860 20692 34862
rect 20860 34524 20916 34580
rect 20860 34242 20916 34244
rect 20860 34190 20862 34242
rect 20862 34190 20914 34242
rect 20914 34190 20916 34242
rect 20860 34188 20916 34190
rect 20412 33234 20468 33236
rect 20412 33182 20414 33234
rect 20414 33182 20466 33234
rect 20466 33182 20468 33234
rect 20412 33180 20468 33182
rect 19516 32508 19572 32564
rect 18620 31388 18676 31444
rect 18508 30716 18564 30772
rect 19404 31388 19460 31444
rect 19292 31052 19348 31108
rect 19068 30492 19124 30548
rect 19404 30716 19460 30772
rect 18508 29708 18564 29764
rect 18396 28364 18452 28420
rect 18956 29260 19012 29316
rect 18732 29036 18788 29092
rect 18284 27132 18340 27188
rect 18396 27020 18452 27076
rect 18732 27746 18788 27748
rect 18732 27694 18734 27746
rect 18734 27694 18786 27746
rect 18786 27694 18788 27746
rect 18732 27692 18788 27694
rect 19068 28364 19124 28420
rect 18956 27074 19012 27076
rect 18956 27022 18958 27074
rect 18958 27022 19010 27074
rect 19010 27022 19012 27074
rect 18956 27020 19012 27022
rect 19068 26908 19124 26964
rect 17612 26572 17668 26628
rect 17500 25788 17556 25844
rect 17724 24722 17780 24724
rect 17724 24670 17726 24722
rect 17726 24670 17778 24722
rect 17778 24670 17780 24722
rect 17724 24668 17780 24670
rect 18284 26290 18340 26292
rect 18284 26238 18286 26290
rect 18286 26238 18338 26290
rect 18338 26238 18340 26290
rect 18284 26236 18340 26238
rect 18060 25506 18116 25508
rect 18060 25454 18062 25506
rect 18062 25454 18114 25506
rect 18114 25454 18116 25506
rect 18060 25452 18116 25454
rect 18732 25788 18788 25844
rect 18956 25676 19012 25732
rect 18620 25282 18676 25284
rect 18620 25230 18622 25282
rect 18622 25230 18674 25282
rect 18674 25230 18676 25282
rect 18620 25228 18676 25230
rect 19516 30268 19572 30324
rect 19292 30210 19348 30212
rect 19292 30158 19294 30210
rect 19294 30158 19346 30210
rect 19346 30158 19348 30210
rect 19292 30156 19348 30158
rect 20188 32284 20244 32340
rect 19852 31890 19908 31892
rect 19852 31838 19854 31890
rect 19854 31838 19906 31890
rect 19906 31838 19908 31890
rect 19852 31836 19908 31838
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20748 32508 20804 32564
rect 20412 31836 20468 31892
rect 20300 30994 20356 30996
rect 20300 30942 20302 30994
rect 20302 30942 20354 30994
rect 20354 30942 20356 30994
rect 20300 30940 20356 30942
rect 20412 31500 20468 31556
rect 20524 30268 20580 30324
rect 19628 30156 19684 30212
rect 20412 30210 20468 30212
rect 20412 30158 20414 30210
rect 20414 30158 20466 30210
rect 20466 30158 20468 30210
rect 20412 30156 20468 30158
rect 19404 28364 19460 28420
rect 19292 26684 19348 26740
rect 19292 26236 19348 26292
rect 19628 29986 19684 29988
rect 19628 29934 19630 29986
rect 19630 29934 19682 29986
rect 19682 29934 19684 29986
rect 19628 29932 19684 29934
rect 20076 29986 20132 29988
rect 20076 29934 20078 29986
rect 20078 29934 20130 29986
rect 20130 29934 20132 29986
rect 20076 29932 20132 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20860 32732 20916 32788
rect 20636 29484 20692 29540
rect 20300 29148 20356 29204
rect 20188 28754 20244 28756
rect 20188 28702 20190 28754
rect 20190 28702 20242 28754
rect 20242 28702 20244 28754
rect 20188 28700 20244 28702
rect 19628 28642 19684 28644
rect 19628 28590 19630 28642
rect 19630 28590 19682 28642
rect 19682 28590 19684 28642
rect 19628 28588 19684 28590
rect 20076 28418 20132 28420
rect 20076 28366 20078 28418
rect 20078 28366 20130 28418
rect 20130 28366 20132 28418
rect 20076 28364 20132 28366
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 28252 20244 28308
rect 19516 27970 19572 27972
rect 19516 27918 19518 27970
rect 19518 27918 19570 27970
rect 19570 27918 19572 27970
rect 19516 27916 19572 27918
rect 21308 36258 21364 36260
rect 21308 36206 21310 36258
rect 21310 36206 21362 36258
rect 21362 36206 21364 36258
rect 21308 36204 21364 36206
rect 21420 34748 21476 34804
rect 21532 34690 21588 34692
rect 21532 34638 21534 34690
rect 21534 34638 21586 34690
rect 21586 34638 21588 34690
rect 21532 34636 21588 34638
rect 21756 35196 21812 35252
rect 21420 33852 21476 33908
rect 21868 34914 21924 34916
rect 21868 34862 21870 34914
rect 21870 34862 21922 34914
rect 21922 34862 21924 34914
rect 21868 34860 21924 34862
rect 21420 32732 21476 32788
rect 21868 34636 21924 34692
rect 21420 31836 21476 31892
rect 21308 31778 21364 31780
rect 21308 31726 21310 31778
rect 21310 31726 21362 31778
rect 21362 31726 21364 31778
rect 21308 31724 21364 31726
rect 21084 31106 21140 31108
rect 21084 31054 21086 31106
rect 21086 31054 21138 31106
rect 21138 31054 21140 31106
rect 21084 31052 21140 31054
rect 21420 30716 21476 30772
rect 21980 34130 22036 34132
rect 21980 34078 21982 34130
rect 21982 34078 22034 34130
rect 22034 34078 22036 34130
rect 21980 34076 22036 34078
rect 22316 33964 22372 34020
rect 21980 33570 22036 33572
rect 21980 33518 21982 33570
rect 21982 33518 22034 33570
rect 22034 33518 22036 33570
rect 21980 33516 22036 33518
rect 21980 32956 22036 33012
rect 21532 30156 21588 30212
rect 21756 30994 21812 30996
rect 21756 30942 21758 30994
rect 21758 30942 21810 30994
rect 21810 30942 21812 30994
rect 21756 30940 21812 30942
rect 21308 29820 21364 29876
rect 20860 28812 20916 28868
rect 22876 39004 22932 39060
rect 23436 42924 23492 42980
rect 23548 43596 23604 43652
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 30604 44322 30660 44324
rect 30604 44270 30606 44322
rect 30606 44270 30658 44322
rect 30658 44270 30660 44322
rect 30604 44268 30660 44270
rect 27804 43708 27860 43764
rect 28476 43820 28532 43876
rect 24220 42476 24276 42532
rect 23436 41074 23492 41076
rect 23436 41022 23438 41074
rect 23438 41022 23490 41074
rect 23490 41022 23492 41074
rect 23436 41020 23492 41022
rect 23212 40514 23268 40516
rect 23212 40462 23214 40514
rect 23214 40462 23266 40514
rect 23266 40462 23268 40514
rect 23212 40460 23268 40462
rect 23100 39058 23156 39060
rect 23100 39006 23102 39058
rect 23102 39006 23154 39058
rect 23154 39006 23156 39058
rect 23100 39004 23156 39006
rect 23212 39452 23268 39508
rect 23548 40626 23604 40628
rect 23548 40574 23550 40626
rect 23550 40574 23602 40626
rect 23602 40574 23604 40626
rect 23548 40572 23604 40574
rect 23324 38946 23380 38948
rect 23324 38894 23326 38946
rect 23326 38894 23378 38946
rect 23378 38894 23380 38946
rect 23324 38892 23380 38894
rect 22540 38220 22596 38276
rect 23548 40236 23604 40292
rect 22540 38050 22596 38052
rect 22540 37998 22542 38050
rect 22542 37998 22594 38050
rect 22594 37998 22596 38050
rect 22540 37996 22596 37998
rect 22540 35756 22596 35812
rect 22876 36258 22932 36260
rect 22876 36206 22878 36258
rect 22878 36206 22930 36258
rect 22930 36206 22932 36258
rect 22876 36204 22932 36206
rect 23212 36876 23268 36932
rect 22988 35196 23044 35252
rect 23212 35868 23268 35924
rect 22652 34354 22708 34356
rect 22652 34302 22654 34354
rect 22654 34302 22706 34354
rect 22706 34302 22708 34354
rect 22652 34300 22708 34302
rect 23212 34524 23268 34580
rect 24220 41186 24276 41188
rect 24220 41134 24222 41186
rect 24222 41134 24274 41186
rect 24274 41134 24276 41186
rect 24220 41132 24276 41134
rect 24444 41916 24500 41972
rect 25004 43484 25060 43540
rect 24668 42588 24724 42644
rect 24780 42476 24836 42532
rect 25676 43538 25732 43540
rect 25676 43486 25678 43538
rect 25678 43486 25730 43538
rect 25730 43486 25732 43538
rect 25676 43484 25732 43486
rect 26460 43426 26516 43428
rect 26460 43374 26462 43426
rect 26462 43374 26514 43426
rect 26514 43374 26516 43426
rect 26460 43372 26516 43374
rect 25788 43148 25844 43204
rect 26684 42924 26740 42980
rect 26348 42754 26404 42756
rect 26348 42702 26350 42754
rect 26350 42702 26402 42754
rect 26402 42702 26404 42754
rect 26348 42700 26404 42702
rect 26124 42642 26180 42644
rect 26124 42590 26126 42642
rect 26126 42590 26178 42642
rect 26178 42590 26180 42642
rect 26124 42588 26180 42590
rect 28700 43484 28756 43540
rect 28476 42588 28532 42644
rect 26572 42364 26628 42420
rect 25340 41356 25396 41412
rect 27132 41356 27188 41412
rect 24556 41132 24612 41188
rect 24332 40684 24388 40740
rect 23660 40124 23716 40180
rect 23660 39004 23716 39060
rect 23548 36876 23604 36932
rect 24332 40124 24388 40180
rect 24108 39004 24164 39060
rect 25340 41186 25396 41188
rect 25340 41134 25342 41186
rect 25342 41134 25394 41186
rect 25394 41134 25396 41186
rect 25340 41132 25396 41134
rect 26012 40572 26068 40628
rect 27692 40908 27748 40964
rect 27356 40402 27412 40404
rect 27356 40350 27358 40402
rect 27358 40350 27410 40402
rect 27410 40350 27412 40402
rect 27356 40348 27412 40350
rect 25116 39116 25172 39172
rect 26572 39228 26628 39284
rect 26348 39004 26404 39060
rect 24444 38834 24500 38836
rect 24444 38782 24446 38834
rect 24446 38782 24498 38834
rect 24498 38782 24500 38834
rect 24444 38780 24500 38782
rect 25116 38780 25172 38836
rect 24332 38668 24388 38724
rect 23884 38220 23940 38276
rect 24108 37378 24164 37380
rect 24108 37326 24110 37378
rect 24110 37326 24162 37378
rect 24162 37326 24164 37378
rect 24108 37324 24164 37326
rect 25228 38722 25284 38724
rect 25228 38670 25230 38722
rect 25230 38670 25282 38722
rect 25282 38670 25284 38722
rect 25228 38668 25284 38670
rect 26124 38722 26180 38724
rect 26124 38670 26126 38722
rect 26126 38670 26178 38722
rect 26178 38670 26180 38722
rect 26124 38668 26180 38670
rect 25452 37996 25508 38052
rect 24668 37266 24724 37268
rect 24668 37214 24670 37266
rect 24670 37214 24722 37266
rect 24722 37214 24724 37266
rect 24668 37212 24724 37214
rect 25452 36988 25508 37044
rect 23100 34188 23156 34244
rect 23772 35868 23828 35924
rect 23100 33906 23156 33908
rect 23100 33854 23102 33906
rect 23102 33854 23154 33906
rect 23154 33854 23156 33906
rect 23100 33852 23156 33854
rect 25228 35922 25284 35924
rect 25228 35870 25230 35922
rect 25230 35870 25282 35922
rect 25282 35870 25284 35922
rect 25228 35868 25284 35870
rect 23772 34300 23828 34356
rect 24108 34130 24164 34132
rect 24108 34078 24110 34130
rect 24110 34078 24162 34130
rect 24162 34078 24164 34130
rect 24108 34076 24164 34078
rect 23884 33906 23940 33908
rect 23884 33854 23886 33906
rect 23886 33854 23938 33906
rect 23938 33854 23940 33906
rect 23884 33852 23940 33854
rect 23212 33516 23268 33572
rect 23996 33740 24052 33796
rect 22764 33234 22820 33236
rect 22764 33182 22766 33234
rect 22766 33182 22818 33234
rect 22818 33182 22820 33234
rect 22764 33180 22820 33182
rect 23436 33180 23492 33236
rect 22428 32284 22484 32340
rect 22988 32562 23044 32564
rect 22988 32510 22990 32562
rect 22990 32510 23042 32562
rect 23042 32510 23044 32562
rect 22988 32508 23044 32510
rect 23324 32562 23380 32564
rect 23324 32510 23326 32562
rect 23326 32510 23378 32562
rect 23378 32510 23380 32562
rect 23324 32508 23380 32510
rect 23436 32284 23492 32340
rect 23212 31612 23268 31668
rect 22316 30268 22372 30324
rect 21756 29820 21812 29876
rect 21532 29260 21588 29316
rect 20300 28028 20356 28084
rect 20188 27916 20244 27972
rect 19740 26796 19796 26852
rect 20636 27580 20692 27636
rect 20748 28588 20804 28644
rect 20412 26908 20468 26964
rect 20076 26796 20132 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19404 25676 19460 25732
rect 20412 26124 20468 26180
rect 20188 25564 20244 25620
rect 20300 25506 20356 25508
rect 20300 25454 20302 25506
rect 20302 25454 20354 25506
rect 20354 25454 20356 25506
rect 20300 25452 20356 25454
rect 17724 22876 17780 22932
rect 18284 23154 18340 23156
rect 18284 23102 18286 23154
rect 18286 23102 18338 23154
rect 18338 23102 18340 23154
rect 18284 23100 18340 23102
rect 17164 22316 17220 22372
rect 17724 22316 17780 22372
rect 17388 20300 17444 20356
rect 17164 20188 17220 20244
rect 17052 20076 17108 20132
rect 17948 21756 18004 21812
rect 18396 21756 18452 21812
rect 19068 23100 19124 23156
rect 19180 22428 19236 22484
rect 18508 21308 18564 21364
rect 18172 20748 18228 20804
rect 18172 20188 18228 20244
rect 17836 20130 17892 20132
rect 17836 20078 17838 20130
rect 17838 20078 17890 20130
rect 17890 20078 17892 20130
rect 17836 20076 17892 20078
rect 17948 19906 18004 19908
rect 17948 19854 17950 19906
rect 17950 19854 18002 19906
rect 18002 19854 18004 19906
rect 17948 19852 18004 19854
rect 18508 20578 18564 20580
rect 18508 20526 18510 20578
rect 18510 20526 18562 20578
rect 18562 20526 18564 20578
rect 18508 20524 18564 20526
rect 18956 20524 19012 20580
rect 18620 20076 18676 20132
rect 18172 19346 18228 19348
rect 18172 19294 18174 19346
rect 18174 19294 18226 19346
rect 18226 19294 18228 19346
rect 18172 19292 18228 19294
rect 17388 18060 17444 18116
rect 17500 18508 17556 18564
rect 19180 20802 19236 20804
rect 19180 20750 19182 20802
rect 19182 20750 19234 20802
rect 19234 20750 19236 20802
rect 19180 20748 19236 20750
rect 19068 20188 19124 20244
rect 19292 20188 19348 20244
rect 18956 20076 19012 20132
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20524 25116 20580 25172
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20412 23714 20468 23716
rect 20412 23662 20414 23714
rect 20414 23662 20466 23714
rect 20466 23662 20468 23714
rect 20412 23660 20468 23662
rect 20524 23548 20580 23604
rect 19740 22540 19796 22596
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19852 20802 19908 20804
rect 19852 20750 19854 20802
rect 19854 20750 19906 20802
rect 19906 20750 19908 20802
rect 19852 20748 19908 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20300 22764 20356 22820
rect 21644 28812 21700 28868
rect 21532 28476 21588 28532
rect 22764 30210 22820 30212
rect 22764 30158 22766 30210
rect 22766 30158 22818 30210
rect 22818 30158 22820 30210
rect 22764 30156 22820 30158
rect 22428 29986 22484 29988
rect 22428 29934 22430 29986
rect 22430 29934 22482 29986
rect 22482 29934 22484 29986
rect 22428 29932 22484 29934
rect 22764 29932 22820 29988
rect 22428 29426 22484 29428
rect 22428 29374 22430 29426
rect 22430 29374 22482 29426
rect 22482 29374 22484 29426
rect 22428 29372 22484 29374
rect 22428 29148 22484 29204
rect 21980 28812 22036 28868
rect 21756 27916 21812 27972
rect 21308 26796 21364 26852
rect 20748 23772 20804 23828
rect 20636 23154 20692 23156
rect 20636 23102 20638 23154
rect 20638 23102 20690 23154
rect 20690 23102 20692 23154
rect 20636 23100 20692 23102
rect 20972 25452 21028 25508
rect 20524 22540 20580 22596
rect 20300 20412 20356 20468
rect 20188 20188 20244 20244
rect 20076 19404 20132 19460
rect 20524 20076 20580 20132
rect 20412 19292 20468 19348
rect 18844 18732 18900 18788
rect 20412 19122 20468 19124
rect 20412 19070 20414 19122
rect 20414 19070 20466 19122
rect 20466 19070 20468 19122
rect 20412 19068 20468 19070
rect 19516 18732 19572 18788
rect 19292 18396 19348 18452
rect 17500 16940 17556 16996
rect 18284 18060 18340 18116
rect 18396 16828 18452 16884
rect 15820 14812 15876 14868
rect 17724 16044 17780 16100
rect 17836 15932 17892 15988
rect 17612 15708 17668 15764
rect 17836 15596 17892 15652
rect 17948 16210 18004 16212
rect 17948 16158 17950 16210
rect 17950 16158 18002 16210
rect 18002 16158 18004 16210
rect 17948 16156 18004 16158
rect 14588 14028 14644 14084
rect 14700 13692 14756 13748
rect 13804 13580 13860 13636
rect 12908 13132 12964 13188
rect 13692 13132 13748 13188
rect 12908 12962 12964 12964
rect 12908 12910 12910 12962
rect 12910 12910 12962 12962
rect 12962 12910 12964 12962
rect 12908 12908 12964 12910
rect 14252 12962 14308 12964
rect 14252 12910 14254 12962
rect 14254 12910 14306 12962
rect 14306 12910 14308 12962
rect 14252 12908 14308 12910
rect 13804 12684 13860 12740
rect 12908 11282 12964 11284
rect 12908 11230 12910 11282
rect 12910 11230 12962 11282
rect 12962 11230 12964 11282
rect 12908 11228 12964 11230
rect 13356 11282 13412 11284
rect 13356 11230 13358 11282
rect 13358 11230 13410 11282
rect 13410 11230 13412 11282
rect 13356 11228 13412 11230
rect 13692 11282 13748 11284
rect 13692 11230 13694 11282
rect 13694 11230 13746 11282
rect 13746 11230 13748 11282
rect 13692 11228 13748 11230
rect 12908 10444 12964 10500
rect 13020 9884 13076 9940
rect 13020 8876 13076 8932
rect 16156 12348 16212 12404
rect 15820 11732 15876 11788
rect 15484 11564 15540 11620
rect 15820 11564 15876 11620
rect 15484 11340 15540 11396
rect 15260 11282 15316 11284
rect 15260 11230 15262 11282
rect 15262 11230 15314 11282
rect 15314 11230 15316 11282
rect 15260 11228 15316 11230
rect 15148 11170 15204 11172
rect 15148 11118 15150 11170
rect 15150 11118 15202 11170
rect 15202 11118 15204 11170
rect 15148 11116 15204 11118
rect 15596 11228 15652 11284
rect 16268 12290 16324 12292
rect 16268 12238 16270 12290
rect 16270 12238 16322 12290
rect 16322 12238 16324 12290
rect 16268 12236 16324 12238
rect 19404 18060 19460 18116
rect 19516 18508 19572 18564
rect 19180 16882 19236 16884
rect 19180 16830 19182 16882
rect 19182 16830 19234 16882
rect 19234 16830 19236 16882
rect 19180 16828 19236 16830
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20076 18620 20132 18676
rect 19964 18450 20020 18452
rect 19964 18398 19966 18450
rect 19966 18398 20018 18450
rect 20018 18398 20020 18450
rect 19964 18396 20020 18398
rect 20188 18562 20244 18564
rect 20188 18510 20190 18562
rect 20190 18510 20242 18562
rect 20242 18510 20244 18562
rect 20188 18508 20244 18510
rect 20412 18450 20468 18452
rect 20412 18398 20414 18450
rect 20414 18398 20466 18450
rect 20466 18398 20468 18450
rect 20412 18396 20468 18398
rect 19628 18172 19684 18228
rect 19852 17778 19908 17780
rect 19852 17726 19854 17778
rect 19854 17726 19906 17778
rect 19906 17726 19908 17778
rect 19852 17724 19908 17726
rect 20188 17388 20244 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20972 21644 21028 21700
rect 21084 25340 21140 25396
rect 21196 25564 21252 25620
rect 21420 26012 21476 26068
rect 22876 29484 22932 29540
rect 22876 29148 22932 29204
rect 22652 28588 22708 28644
rect 21868 26796 21924 26852
rect 21756 26290 21812 26292
rect 21756 26238 21758 26290
rect 21758 26238 21810 26290
rect 21810 26238 21812 26290
rect 21756 26236 21812 26238
rect 21532 24556 21588 24612
rect 21532 23938 21588 23940
rect 21532 23886 21534 23938
rect 21534 23886 21586 23938
rect 21586 23886 21588 23938
rect 21532 23884 21588 23886
rect 21868 23660 21924 23716
rect 21308 23212 21364 23268
rect 21308 22876 21364 22932
rect 21532 22764 21588 22820
rect 21308 21474 21364 21476
rect 21308 21422 21310 21474
rect 21310 21422 21362 21474
rect 21362 21422 21364 21474
rect 21308 21420 21364 21422
rect 21084 21196 21140 21252
rect 21756 22988 21812 23044
rect 22652 26796 22708 26852
rect 22204 26572 22260 26628
rect 22652 26348 22708 26404
rect 22428 26066 22484 26068
rect 22428 26014 22430 26066
rect 22430 26014 22482 26066
rect 22482 26014 22484 26066
rect 22428 26012 22484 26014
rect 22988 27916 23044 27972
rect 23324 30940 23380 30996
rect 23324 30716 23380 30772
rect 23324 29260 23380 29316
rect 23212 28812 23268 28868
rect 23324 28476 23380 28532
rect 23660 31612 23716 31668
rect 23660 31052 23716 31108
rect 26684 39058 26740 39060
rect 26684 39006 26686 39058
rect 26686 39006 26738 39058
rect 26738 39006 26740 39058
rect 26684 39004 26740 39006
rect 26908 39004 26964 39060
rect 27020 38834 27076 38836
rect 27020 38782 27022 38834
rect 27022 38782 27074 38834
rect 27074 38782 27076 38834
rect 27020 38780 27076 38782
rect 27356 39228 27412 39284
rect 27468 39116 27524 39172
rect 28140 42530 28196 42532
rect 28140 42478 28142 42530
rect 28142 42478 28194 42530
rect 28194 42478 28196 42530
rect 28140 42476 28196 42478
rect 29148 43708 29204 43764
rect 28924 42476 28980 42532
rect 29484 43596 29540 43652
rect 29596 43484 29652 43540
rect 29260 42866 29316 42868
rect 29260 42814 29262 42866
rect 29262 42814 29314 42866
rect 29314 42814 29316 42866
rect 29260 42812 29316 42814
rect 29820 42700 29876 42756
rect 28700 42364 28756 42420
rect 28028 41132 28084 41188
rect 28140 41298 28196 41300
rect 28140 41246 28142 41298
rect 28142 41246 28194 41298
rect 28194 41246 28196 41298
rect 28140 41244 28196 41246
rect 28476 40962 28532 40964
rect 28476 40910 28478 40962
rect 28478 40910 28530 40962
rect 28530 40910 28532 40962
rect 28476 40908 28532 40910
rect 28476 40684 28532 40740
rect 28588 40348 28644 40404
rect 27804 39004 27860 39060
rect 26796 38444 26852 38500
rect 26796 37938 26852 37940
rect 26796 37886 26798 37938
rect 26798 37886 26850 37938
rect 26850 37886 26852 37938
rect 26796 37884 26852 37886
rect 26348 36316 26404 36372
rect 25452 35532 25508 35588
rect 25676 35420 25732 35476
rect 25116 35308 25172 35364
rect 25340 34412 25396 34468
rect 24444 34242 24500 34244
rect 24444 34190 24446 34242
rect 24446 34190 24498 34242
rect 24498 34190 24500 34242
rect 24444 34188 24500 34190
rect 25228 34242 25284 34244
rect 25228 34190 25230 34242
rect 25230 34190 25282 34242
rect 25282 34190 25284 34242
rect 25228 34188 25284 34190
rect 25340 33906 25396 33908
rect 25340 33854 25342 33906
rect 25342 33854 25394 33906
rect 25394 33854 25396 33906
rect 25340 33852 25396 33854
rect 25564 33852 25620 33908
rect 24332 33628 24388 33684
rect 26460 35420 26516 35476
rect 25900 33906 25956 33908
rect 25900 33854 25902 33906
rect 25902 33854 25954 33906
rect 25954 33854 25956 33906
rect 25900 33852 25956 33854
rect 25676 33740 25732 33796
rect 26012 33404 26068 33460
rect 26124 33628 26180 33684
rect 24108 32508 24164 32564
rect 24556 32562 24612 32564
rect 24556 32510 24558 32562
rect 24558 32510 24610 32562
rect 24610 32510 24612 32562
rect 24556 32508 24612 32510
rect 24444 32396 24500 32452
rect 24108 31612 24164 31668
rect 24444 32060 24500 32116
rect 24332 29708 24388 29764
rect 23996 28924 24052 28980
rect 22988 26572 23044 26628
rect 23212 26460 23268 26516
rect 23660 27580 23716 27636
rect 22316 25116 22372 25172
rect 22204 23938 22260 23940
rect 22204 23886 22206 23938
rect 22206 23886 22258 23938
rect 22258 23886 22260 23938
rect 22204 23884 22260 23886
rect 22316 24610 22372 24612
rect 22316 24558 22318 24610
rect 22318 24558 22370 24610
rect 22370 24558 22372 24610
rect 22316 24556 22372 24558
rect 22092 23548 22148 23604
rect 21980 22428 22036 22484
rect 22652 25564 22708 25620
rect 22540 24892 22596 24948
rect 22652 25004 22708 25060
rect 23100 25228 23156 25284
rect 23324 25004 23380 25060
rect 23436 26460 23492 26516
rect 23548 26290 23604 26292
rect 23548 26238 23550 26290
rect 23550 26238 23602 26290
rect 23602 26238 23604 26290
rect 23548 26236 23604 26238
rect 23212 24444 23268 24500
rect 22540 23436 22596 23492
rect 22428 23324 22484 23380
rect 20860 20412 20916 20468
rect 21196 20636 21252 20692
rect 22652 22652 22708 22708
rect 21980 21756 22036 21812
rect 21756 20802 21812 20804
rect 21756 20750 21758 20802
rect 21758 20750 21810 20802
rect 21810 20750 21812 20802
rect 21756 20748 21812 20750
rect 22428 21756 22484 21812
rect 22092 20076 22148 20132
rect 20748 19404 20804 19460
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 20636 17724 20692 17780
rect 20524 17442 20580 17444
rect 20524 17390 20526 17442
rect 20526 17390 20578 17442
rect 20578 17390 20580 17442
rect 20524 17388 20580 17390
rect 20524 17106 20580 17108
rect 20524 17054 20526 17106
rect 20526 17054 20578 17106
rect 20578 17054 20580 17106
rect 20524 17052 20580 17054
rect 18732 16156 18788 16212
rect 18284 16044 18340 16100
rect 18172 15820 18228 15876
rect 18732 15708 18788 15764
rect 18956 16098 19012 16100
rect 18956 16046 18958 16098
rect 18958 16046 19010 16098
rect 19010 16046 19012 16098
rect 18956 16044 19012 16046
rect 18844 15260 18900 15316
rect 17500 15202 17556 15204
rect 17500 15150 17502 15202
rect 17502 15150 17554 15202
rect 17554 15150 17556 15202
rect 17500 15148 17556 15150
rect 18396 15148 18452 15204
rect 16604 12348 16660 12404
rect 15932 11340 15988 11396
rect 16044 11170 16100 11172
rect 16044 11118 16046 11170
rect 16046 11118 16098 11170
rect 16098 11118 16100 11170
rect 16044 11116 16100 11118
rect 15372 10556 15428 10612
rect 15820 10610 15876 10612
rect 15820 10558 15822 10610
rect 15822 10558 15874 10610
rect 15874 10558 15876 10610
rect 15820 10556 15876 10558
rect 13468 9772 13524 9828
rect 14140 9212 14196 9268
rect 13804 9100 13860 9156
rect 13692 9042 13748 9044
rect 13692 8990 13694 9042
rect 13694 8990 13746 9042
rect 13746 8990 13748 9042
rect 13692 8988 13748 8990
rect 13244 8876 13300 8932
rect 12908 8146 12964 8148
rect 12908 8094 12910 8146
rect 12910 8094 12962 8146
rect 12962 8094 12964 8146
rect 12908 8092 12964 8094
rect 13804 8034 13860 8036
rect 13804 7982 13806 8034
rect 13806 7982 13858 8034
rect 13858 7982 13860 8034
rect 13804 7980 13860 7982
rect 14140 8146 14196 8148
rect 14140 8094 14142 8146
rect 14142 8094 14194 8146
rect 14194 8094 14196 8146
rect 14140 8092 14196 8094
rect 12908 6972 12964 7028
rect 13132 6748 13188 6804
rect 14028 6748 14084 6804
rect 13244 6636 13300 6692
rect 12796 5964 12852 6020
rect 13020 6524 13076 6580
rect 12908 5852 12964 5908
rect 12572 5404 12628 5460
rect 11564 3388 11620 3444
rect 12124 4396 12180 4452
rect 13132 5068 13188 5124
rect 13916 6466 13972 6468
rect 13916 6414 13918 6466
rect 13918 6414 13970 6466
rect 13970 6414 13972 6466
rect 13916 6412 13972 6414
rect 13580 6076 13636 6132
rect 13916 4508 13972 4564
rect 13580 4450 13636 4452
rect 13580 4398 13582 4450
rect 13582 4398 13634 4450
rect 13634 4398 13636 4450
rect 13580 4396 13636 4398
rect 13356 4226 13412 4228
rect 13356 4174 13358 4226
rect 13358 4174 13410 4226
rect 13410 4174 13412 4226
rect 13356 4172 13412 4174
rect 14700 9266 14756 9268
rect 14700 9214 14702 9266
rect 14702 9214 14754 9266
rect 14754 9214 14756 9266
rect 14700 9212 14756 9214
rect 14476 8764 14532 8820
rect 14588 8876 14644 8932
rect 15148 9154 15204 9156
rect 15148 9102 15150 9154
rect 15150 9102 15202 9154
rect 15202 9102 15204 9154
rect 15148 9100 15204 9102
rect 14812 8370 14868 8372
rect 14812 8318 14814 8370
rect 14814 8318 14866 8370
rect 14866 8318 14868 8370
rect 14812 8316 14868 8318
rect 14364 6636 14420 6692
rect 15148 6972 15204 7028
rect 14252 6578 14308 6580
rect 14252 6526 14254 6578
rect 14254 6526 14306 6578
rect 14306 6526 14308 6578
rect 14252 6524 14308 6526
rect 14476 6466 14532 6468
rect 14476 6414 14478 6466
rect 14478 6414 14530 6466
rect 14530 6414 14532 6466
rect 14476 6412 14532 6414
rect 14812 6466 14868 6468
rect 14812 6414 14814 6466
rect 14814 6414 14866 6466
rect 14866 6414 14868 6466
rect 14812 6412 14868 6414
rect 15596 6802 15652 6804
rect 15596 6750 15598 6802
rect 15598 6750 15650 6802
rect 15650 6750 15652 6802
rect 15596 6748 15652 6750
rect 15260 6412 15316 6468
rect 15708 6578 15764 6580
rect 15708 6526 15710 6578
rect 15710 6526 15762 6578
rect 15762 6526 15764 6578
rect 15708 6524 15764 6526
rect 15372 6130 15428 6132
rect 15372 6078 15374 6130
rect 15374 6078 15426 6130
rect 15426 6078 15428 6130
rect 15372 6076 15428 6078
rect 15820 6466 15876 6468
rect 15820 6414 15822 6466
rect 15822 6414 15874 6466
rect 15874 6414 15876 6466
rect 15820 6412 15876 6414
rect 15484 6300 15540 6356
rect 15820 6018 15876 6020
rect 15820 5966 15822 6018
rect 15822 5966 15874 6018
rect 15874 5966 15876 6018
rect 15820 5964 15876 5966
rect 14700 5404 14756 5460
rect 14700 5180 14756 5236
rect 16604 10556 16660 10612
rect 16604 9548 16660 9604
rect 16156 8930 16212 8932
rect 16156 8878 16158 8930
rect 16158 8878 16210 8930
rect 16210 8878 16212 8930
rect 16156 8876 16212 8878
rect 16492 8876 16548 8932
rect 16380 8316 16436 8372
rect 16380 7980 16436 8036
rect 16044 6748 16100 6804
rect 17052 12348 17108 12404
rect 18396 13020 18452 13076
rect 18172 12796 18228 12852
rect 17836 12402 17892 12404
rect 17836 12350 17838 12402
rect 17838 12350 17890 12402
rect 17890 12350 17892 12402
rect 17836 12348 17892 12350
rect 18732 12684 18788 12740
rect 18396 11788 18452 11844
rect 18396 11452 18452 11508
rect 19180 15708 19236 15764
rect 19964 16770 20020 16772
rect 19964 16718 19966 16770
rect 19966 16718 20018 16770
rect 20018 16718 20020 16770
rect 19964 16716 20020 16718
rect 19404 16210 19460 16212
rect 19404 16158 19406 16210
rect 19406 16158 19458 16210
rect 19458 16158 19460 16210
rect 19404 16156 19460 16158
rect 20412 16940 20468 16996
rect 20300 16604 20356 16660
rect 20300 15986 20356 15988
rect 20300 15934 20302 15986
rect 20302 15934 20354 15986
rect 20354 15934 20356 15986
rect 20300 15932 20356 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20524 15484 20580 15540
rect 19516 15260 19572 15316
rect 20300 15202 20356 15204
rect 20300 15150 20302 15202
rect 20302 15150 20354 15202
rect 20354 15150 20356 15202
rect 20300 15148 20356 15150
rect 17388 11116 17444 11172
rect 20748 16770 20804 16772
rect 20748 16718 20750 16770
rect 20750 16718 20802 16770
rect 20802 16718 20804 16770
rect 20748 16716 20804 16718
rect 20972 19068 21028 19124
rect 21532 19404 21588 19460
rect 22652 21868 22708 21924
rect 22876 23884 22932 23940
rect 22988 23714 23044 23716
rect 22988 23662 22990 23714
rect 22990 23662 23042 23714
rect 23042 23662 23044 23714
rect 22988 23660 23044 23662
rect 22988 23324 23044 23380
rect 23100 23266 23156 23268
rect 23100 23214 23102 23266
rect 23102 23214 23154 23266
rect 23154 23214 23156 23266
rect 23100 23212 23156 23214
rect 23100 22764 23156 22820
rect 23548 24332 23604 24388
rect 22876 21756 22932 21812
rect 23212 21810 23268 21812
rect 23212 21758 23214 21810
rect 23214 21758 23266 21810
rect 23266 21758 23268 21810
rect 23212 21756 23268 21758
rect 22988 21698 23044 21700
rect 22988 21646 22990 21698
rect 22990 21646 23042 21698
rect 23042 21646 23044 21698
rect 22988 21644 23044 21646
rect 22876 21586 22932 21588
rect 22876 21534 22878 21586
rect 22878 21534 22930 21586
rect 22930 21534 22932 21586
rect 22876 21532 22932 21534
rect 22764 20578 22820 20580
rect 22764 20526 22766 20578
rect 22766 20526 22818 20578
rect 22818 20526 22820 20578
rect 22764 20524 22820 20526
rect 23100 21474 23156 21476
rect 23100 21422 23102 21474
rect 23102 21422 23154 21474
rect 23154 21422 23156 21474
rect 23100 21420 23156 21422
rect 22988 20188 23044 20244
rect 23436 23548 23492 23604
rect 21420 19010 21476 19012
rect 21420 18958 21422 19010
rect 21422 18958 21474 19010
rect 21474 18958 21476 19010
rect 21420 18956 21476 18958
rect 21980 18956 22036 19012
rect 21756 18450 21812 18452
rect 21756 18398 21758 18450
rect 21758 18398 21810 18450
rect 21810 18398 21812 18450
rect 21756 18396 21812 18398
rect 21644 18338 21700 18340
rect 21644 18286 21646 18338
rect 21646 18286 21698 18338
rect 21698 18286 21700 18338
rect 21644 18284 21700 18286
rect 21532 18060 21588 18116
rect 20860 15426 20916 15428
rect 20860 15374 20862 15426
rect 20862 15374 20914 15426
rect 20914 15374 20916 15426
rect 20860 15372 20916 15374
rect 20076 14700 20132 14756
rect 20076 14418 20132 14420
rect 20076 14366 20078 14418
rect 20078 14366 20130 14418
rect 20130 14366 20132 14418
rect 20076 14364 20132 14366
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19180 13692 19236 13748
rect 19180 13074 19236 13076
rect 19180 13022 19182 13074
rect 19182 13022 19234 13074
rect 19234 13022 19236 13074
rect 19180 13020 19236 13022
rect 19516 12850 19572 12852
rect 19516 12798 19518 12850
rect 19518 12798 19570 12850
rect 19570 12798 19572 12850
rect 19516 12796 19572 12798
rect 19852 12738 19908 12740
rect 19852 12686 19854 12738
rect 19854 12686 19906 12738
rect 19906 12686 19908 12738
rect 19852 12684 19908 12686
rect 19628 12572 19684 12628
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20188 12460 20244 12516
rect 19292 12290 19348 12292
rect 19292 12238 19294 12290
rect 19294 12238 19346 12290
rect 19346 12238 19348 12290
rect 19292 12236 19348 12238
rect 19180 12124 19236 12180
rect 20076 12178 20132 12180
rect 20076 12126 20078 12178
rect 20078 12126 20130 12178
rect 20130 12126 20132 12178
rect 20076 12124 20132 12126
rect 20300 11788 20356 11844
rect 20188 11506 20244 11508
rect 20188 11454 20190 11506
rect 20190 11454 20242 11506
rect 20242 11454 20244 11506
rect 20188 11452 20244 11454
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 22316 18396 22372 18452
rect 22428 18172 22484 18228
rect 22540 17948 22596 18004
rect 23660 23154 23716 23156
rect 23660 23102 23662 23154
rect 23662 23102 23714 23154
rect 23714 23102 23716 23154
rect 23660 23100 23716 23102
rect 23660 22876 23716 22932
rect 24108 25228 24164 25284
rect 23996 24946 24052 24948
rect 23996 24894 23998 24946
rect 23998 24894 24050 24946
rect 24050 24894 24052 24946
rect 23996 24892 24052 24894
rect 24556 31948 24612 32004
rect 25452 33068 25508 33124
rect 25228 32620 25284 32676
rect 24780 31836 24836 31892
rect 24668 31052 24724 31108
rect 24668 30156 24724 30212
rect 24556 29650 24612 29652
rect 24556 29598 24558 29650
rect 24558 29598 24610 29650
rect 24610 29598 24612 29650
rect 24556 29596 24612 29598
rect 25452 32060 25508 32116
rect 25340 30156 25396 30212
rect 24892 30098 24948 30100
rect 24892 30046 24894 30098
rect 24894 30046 24946 30098
rect 24946 30046 24948 30098
rect 24892 30044 24948 30046
rect 24444 29426 24500 29428
rect 24444 29374 24446 29426
rect 24446 29374 24498 29426
rect 24498 29374 24500 29426
rect 24444 29372 24500 29374
rect 24556 28476 24612 28532
rect 25564 31836 25620 31892
rect 25340 29820 25396 29876
rect 25228 29596 25284 29652
rect 25452 28866 25508 28868
rect 25452 28814 25454 28866
rect 25454 28814 25506 28866
rect 25506 28814 25508 28866
rect 25452 28812 25508 28814
rect 25676 29986 25732 29988
rect 25676 29934 25678 29986
rect 25678 29934 25730 29986
rect 25730 29934 25732 29986
rect 25676 29932 25732 29934
rect 25564 29148 25620 29204
rect 24892 28754 24948 28756
rect 24892 28702 24894 28754
rect 24894 28702 24946 28754
rect 24946 28702 24948 28754
rect 24892 28700 24948 28702
rect 24668 27356 24724 27412
rect 24556 27132 24612 27188
rect 25340 28754 25396 28756
rect 25340 28702 25342 28754
rect 25342 28702 25394 28754
rect 25394 28702 25396 28754
rect 25340 28700 25396 28702
rect 27580 38668 27636 38724
rect 27244 37884 27300 37940
rect 27132 35980 27188 36036
rect 27244 35756 27300 35812
rect 26572 32732 26628 32788
rect 26908 34636 26964 34692
rect 26348 32674 26404 32676
rect 26348 32622 26350 32674
rect 26350 32622 26402 32674
rect 26402 32622 26404 32674
rect 26348 32620 26404 32622
rect 26908 32508 26964 32564
rect 26572 31948 26628 32004
rect 27020 31724 27076 31780
rect 27468 35308 27524 35364
rect 27356 34636 27412 34692
rect 27692 38050 27748 38052
rect 27692 37998 27694 38050
rect 27694 37998 27746 38050
rect 27746 37998 27748 38050
rect 27692 37996 27748 37998
rect 27692 37548 27748 37604
rect 27916 38892 27972 38948
rect 28028 39116 28084 39172
rect 28700 40178 28756 40180
rect 28700 40126 28702 40178
rect 28702 40126 28754 40178
rect 28754 40126 28756 40178
rect 28700 40124 28756 40126
rect 28476 39004 28532 39060
rect 28588 38892 28644 38948
rect 28028 38668 28084 38724
rect 28700 38668 28756 38724
rect 28364 37996 28420 38052
rect 28924 40012 28980 40068
rect 28924 39452 28980 39508
rect 28812 38108 28868 38164
rect 28252 37938 28308 37940
rect 28252 37886 28254 37938
rect 28254 37886 28306 37938
rect 28306 37886 28308 37938
rect 28252 37884 28308 37886
rect 28140 37826 28196 37828
rect 28140 37774 28142 37826
rect 28142 37774 28194 37826
rect 28194 37774 28196 37826
rect 28140 37772 28196 37774
rect 28140 37548 28196 37604
rect 28252 36204 28308 36260
rect 28364 36092 28420 36148
rect 27804 34412 27860 34468
rect 27244 32956 27300 33012
rect 28588 34690 28644 34692
rect 28588 34638 28590 34690
rect 28590 34638 28642 34690
rect 28642 34638 28644 34690
rect 28588 34636 28644 34638
rect 28364 34018 28420 34020
rect 28364 33966 28366 34018
rect 28366 33966 28418 34018
rect 28418 33966 28420 34018
rect 28364 33964 28420 33966
rect 28700 33516 28756 33572
rect 28252 33458 28308 33460
rect 28252 33406 28254 33458
rect 28254 33406 28306 33458
rect 28306 33406 28308 33458
rect 28252 33404 28308 33406
rect 28140 33234 28196 33236
rect 28140 33182 28142 33234
rect 28142 33182 28194 33234
rect 28194 33182 28196 33234
rect 28140 33180 28196 33182
rect 28588 33346 28644 33348
rect 28588 33294 28590 33346
rect 28590 33294 28642 33346
rect 28642 33294 28644 33346
rect 28588 33292 28644 33294
rect 28364 33068 28420 33124
rect 27468 31948 27524 32004
rect 27692 32450 27748 32452
rect 27692 32398 27694 32450
rect 27694 32398 27746 32450
rect 27746 32398 27748 32450
rect 27692 32396 27748 32398
rect 27580 31836 27636 31892
rect 26124 30716 26180 30772
rect 25900 30044 25956 30100
rect 26348 30044 26404 30100
rect 25788 29036 25844 29092
rect 26012 29036 26068 29092
rect 25228 26908 25284 26964
rect 24556 25340 24612 25396
rect 24444 24498 24500 24500
rect 24444 24446 24446 24498
rect 24446 24446 24498 24498
rect 24498 24446 24500 24498
rect 24444 24444 24500 24446
rect 24220 23266 24276 23268
rect 24220 23214 24222 23266
rect 24222 23214 24274 23266
rect 24274 23214 24276 23266
rect 24220 23212 24276 23214
rect 23884 22540 23940 22596
rect 24332 22092 24388 22148
rect 24332 21810 24388 21812
rect 24332 21758 24334 21810
rect 24334 21758 24386 21810
rect 24386 21758 24388 21810
rect 24332 21756 24388 21758
rect 24108 21698 24164 21700
rect 24108 21646 24110 21698
rect 24110 21646 24162 21698
rect 24162 21646 24164 21698
rect 24108 21644 24164 21646
rect 23996 21586 24052 21588
rect 23996 21534 23998 21586
rect 23998 21534 24050 21586
rect 24050 21534 24052 21586
rect 23996 21532 24052 21534
rect 23772 21420 23828 21476
rect 23100 18956 23156 19012
rect 21868 15874 21924 15876
rect 21868 15822 21870 15874
rect 21870 15822 21922 15874
rect 21922 15822 21924 15874
rect 21868 15820 21924 15822
rect 22876 18284 22932 18340
rect 22988 18060 23044 18116
rect 24220 20636 24276 20692
rect 24332 20188 24388 20244
rect 23436 20076 23492 20132
rect 23324 19964 23380 20020
rect 23324 18450 23380 18452
rect 23324 18398 23326 18450
rect 23326 18398 23378 18450
rect 23378 18398 23380 18450
rect 23324 18396 23380 18398
rect 23772 20018 23828 20020
rect 23772 19966 23774 20018
rect 23774 19966 23826 20018
rect 23826 19966 23828 20018
rect 23772 19964 23828 19966
rect 24556 23324 24612 23380
rect 25788 28530 25844 28532
rect 25788 28478 25790 28530
rect 25790 28478 25842 28530
rect 25842 28478 25844 28530
rect 25788 28476 25844 28478
rect 26684 31106 26740 31108
rect 26684 31054 26686 31106
rect 26686 31054 26738 31106
rect 26738 31054 26740 31106
rect 26684 31052 26740 31054
rect 26460 29708 26516 29764
rect 26684 30716 26740 30772
rect 26796 30322 26852 30324
rect 26796 30270 26798 30322
rect 26798 30270 26850 30322
rect 26850 30270 26852 30322
rect 26796 30268 26852 30270
rect 26908 29986 26964 29988
rect 26908 29934 26910 29986
rect 26910 29934 26962 29986
rect 26962 29934 26964 29986
rect 26908 29932 26964 29934
rect 26572 29036 26628 29092
rect 26236 28700 26292 28756
rect 26236 28418 26292 28420
rect 26236 28366 26238 28418
rect 26238 28366 26290 28418
rect 26290 28366 26292 28418
rect 26236 28364 26292 28366
rect 26124 27916 26180 27972
rect 26572 28812 26628 28868
rect 26796 28812 26852 28868
rect 26572 28364 26628 28420
rect 25452 26796 25508 26852
rect 26124 26850 26180 26852
rect 26124 26798 26126 26850
rect 26126 26798 26178 26850
rect 26178 26798 26180 26850
rect 26124 26796 26180 26798
rect 26012 26348 26068 26404
rect 26236 26402 26292 26404
rect 26236 26350 26238 26402
rect 26238 26350 26290 26402
rect 26290 26350 26292 26402
rect 26236 26348 26292 26350
rect 25564 25676 25620 25732
rect 25452 25394 25508 25396
rect 25452 25342 25454 25394
rect 25454 25342 25506 25394
rect 25506 25342 25508 25394
rect 25452 25340 25508 25342
rect 25340 25282 25396 25284
rect 25340 25230 25342 25282
rect 25342 25230 25394 25282
rect 25394 25230 25396 25282
rect 25340 25228 25396 25230
rect 26124 25228 26180 25284
rect 25676 24108 25732 24164
rect 25340 23826 25396 23828
rect 25340 23774 25342 23826
rect 25342 23774 25394 23826
rect 25394 23774 25396 23826
rect 25340 23772 25396 23774
rect 25228 23100 25284 23156
rect 25564 23154 25620 23156
rect 25564 23102 25566 23154
rect 25566 23102 25618 23154
rect 25618 23102 25620 23154
rect 25564 23100 25620 23102
rect 25900 23378 25956 23380
rect 25900 23326 25902 23378
rect 25902 23326 25954 23378
rect 25954 23326 25956 23378
rect 25900 23324 25956 23326
rect 26236 23436 26292 23492
rect 26124 23378 26180 23380
rect 26124 23326 26126 23378
rect 26126 23326 26178 23378
rect 26178 23326 26180 23378
rect 26124 23324 26180 23326
rect 26012 23266 26068 23268
rect 26012 23214 26014 23266
rect 26014 23214 26066 23266
rect 26066 23214 26068 23266
rect 26012 23212 26068 23214
rect 25788 23100 25844 23156
rect 26460 27074 26516 27076
rect 26460 27022 26462 27074
rect 26462 27022 26514 27074
rect 26514 27022 26516 27074
rect 26460 27020 26516 27022
rect 26460 26684 26516 26740
rect 25788 22652 25844 22708
rect 25452 22146 25508 22148
rect 25452 22094 25454 22146
rect 25454 22094 25506 22146
rect 25506 22094 25508 22146
rect 25452 22092 25508 22094
rect 26796 25394 26852 25396
rect 26796 25342 26798 25394
rect 26798 25342 26850 25394
rect 26850 25342 26852 25394
rect 26796 25340 26852 25342
rect 26572 24108 26628 24164
rect 26796 24780 26852 24836
rect 26796 23660 26852 23716
rect 26684 23436 26740 23492
rect 26572 23042 26628 23044
rect 26572 22990 26574 23042
rect 26574 22990 26626 23042
rect 26626 22990 26628 23042
rect 26572 22988 26628 22990
rect 27244 30268 27300 30324
rect 28140 32508 28196 32564
rect 28028 32002 28084 32004
rect 28028 31950 28030 32002
rect 28030 31950 28082 32002
rect 28082 31950 28084 32002
rect 28028 31948 28084 31950
rect 27916 31106 27972 31108
rect 27916 31054 27918 31106
rect 27918 31054 27970 31106
rect 27970 31054 27972 31106
rect 27916 31052 27972 31054
rect 28364 32172 28420 32228
rect 28364 31388 28420 31444
rect 29148 39340 29204 39396
rect 29484 40572 29540 40628
rect 29372 40514 29428 40516
rect 29372 40462 29374 40514
rect 29374 40462 29426 40514
rect 29426 40462 29428 40514
rect 29372 40460 29428 40462
rect 29484 40012 29540 40068
rect 29708 40908 29764 40964
rect 30268 43596 30324 43652
rect 30156 43260 30212 43316
rect 30044 42754 30100 42756
rect 30044 42702 30046 42754
rect 30046 42702 30098 42754
rect 30098 42702 30100 42754
rect 30044 42700 30100 42702
rect 30492 43260 30548 43316
rect 31052 43708 31108 43764
rect 31836 43708 31892 43764
rect 31388 43426 31444 43428
rect 31388 43374 31390 43426
rect 31390 43374 31442 43426
rect 31442 43374 31444 43426
rect 31388 43372 31444 43374
rect 31276 43260 31332 43316
rect 31052 43148 31108 43204
rect 29932 41916 29988 41972
rect 30156 42476 30212 42532
rect 30268 42252 30324 42308
rect 30044 41356 30100 41412
rect 30268 41298 30324 41300
rect 30268 41246 30270 41298
rect 30270 41246 30322 41298
rect 30322 41246 30324 41298
rect 30268 41244 30324 41246
rect 30716 42754 30772 42756
rect 30716 42702 30718 42754
rect 30718 42702 30770 42754
rect 30770 42702 30772 42754
rect 30716 42700 30772 42702
rect 30716 41356 30772 41412
rect 39228 44434 39284 44436
rect 39228 44382 39230 44434
rect 39230 44382 39282 44434
rect 39282 44382 39284 44434
rect 39228 44380 39284 44382
rect 32620 43650 32676 43652
rect 32620 43598 32622 43650
rect 32622 43598 32674 43650
rect 32674 43598 32676 43650
rect 32620 43596 32676 43598
rect 32844 43372 32900 43428
rect 32284 42812 32340 42868
rect 31164 41970 31220 41972
rect 31164 41918 31166 41970
rect 31166 41918 31218 41970
rect 31218 41918 31220 41970
rect 31164 41916 31220 41918
rect 31500 42530 31556 42532
rect 31500 42478 31502 42530
rect 31502 42478 31554 42530
rect 31554 42478 31556 42530
rect 31500 42476 31556 42478
rect 31948 42530 32004 42532
rect 31948 42478 31950 42530
rect 31950 42478 32002 42530
rect 32002 42478 32004 42530
rect 31948 42476 32004 42478
rect 31388 41356 31444 41412
rect 31276 40962 31332 40964
rect 31276 40910 31278 40962
rect 31278 40910 31330 40962
rect 31330 40910 31332 40962
rect 31276 40908 31332 40910
rect 31164 40796 31220 40852
rect 30492 40684 30548 40740
rect 30716 40684 30772 40740
rect 30492 40514 30548 40516
rect 30492 40462 30494 40514
rect 30494 40462 30546 40514
rect 30546 40462 30548 40514
rect 30492 40460 30548 40462
rect 30716 40514 30772 40516
rect 30716 40462 30718 40514
rect 30718 40462 30770 40514
rect 30770 40462 30772 40514
rect 30716 40460 30772 40462
rect 30268 39900 30324 39956
rect 29708 39730 29764 39732
rect 29708 39678 29710 39730
rect 29710 39678 29762 39730
rect 29762 39678 29764 39730
rect 29708 39676 29764 39678
rect 29820 39618 29876 39620
rect 29820 39566 29822 39618
rect 29822 39566 29874 39618
rect 29874 39566 29876 39618
rect 29820 39564 29876 39566
rect 29148 39116 29204 39172
rect 29372 38946 29428 38948
rect 29372 38894 29374 38946
rect 29374 38894 29426 38946
rect 29426 38894 29428 38946
rect 29372 38892 29428 38894
rect 29260 38834 29316 38836
rect 29260 38782 29262 38834
rect 29262 38782 29314 38834
rect 29314 38782 29316 38834
rect 29260 38780 29316 38782
rect 29148 38556 29204 38612
rect 29708 39340 29764 39396
rect 29596 38892 29652 38948
rect 29372 38050 29428 38052
rect 29372 37998 29374 38050
rect 29374 37998 29426 38050
rect 29426 37998 29428 38050
rect 29372 37996 29428 37998
rect 29148 37938 29204 37940
rect 29148 37886 29150 37938
rect 29150 37886 29202 37938
rect 29202 37886 29204 37938
rect 29148 37884 29204 37886
rect 29372 36428 29428 36484
rect 29260 35868 29316 35924
rect 29596 36370 29652 36372
rect 29596 36318 29598 36370
rect 29598 36318 29650 36370
rect 29650 36318 29652 36370
rect 29596 36316 29652 36318
rect 29148 35420 29204 35476
rect 29820 39116 29876 39172
rect 32172 41356 32228 41412
rect 33516 44210 33572 44212
rect 33516 44158 33518 44210
rect 33518 44158 33570 44210
rect 33570 44158 33572 44210
rect 33516 44156 33572 44158
rect 33404 43932 33460 43988
rect 32956 42812 33012 42868
rect 32396 42252 32452 42308
rect 32508 42588 32564 42644
rect 31948 41074 32004 41076
rect 31948 41022 31950 41074
rect 31950 41022 32002 41074
rect 32002 41022 32004 41074
rect 31948 41020 32004 41022
rect 31724 40460 31780 40516
rect 31388 40290 31444 40292
rect 31388 40238 31390 40290
rect 31390 40238 31442 40290
rect 31442 40238 31444 40290
rect 31388 40236 31444 40238
rect 30828 39900 30884 39956
rect 31276 40012 31332 40068
rect 30380 39564 30436 39620
rect 30492 39676 30548 39732
rect 30268 38892 30324 38948
rect 30716 39340 30772 39396
rect 30828 39228 30884 39284
rect 29932 38556 29988 38612
rect 30156 38108 30212 38164
rect 30492 38050 30548 38052
rect 30492 37998 30494 38050
rect 30494 37998 30546 38050
rect 30546 37998 30548 38050
rect 30492 37996 30548 37998
rect 30604 38444 30660 38500
rect 30268 37826 30324 37828
rect 30268 37774 30270 37826
rect 30270 37774 30322 37826
rect 30322 37774 30324 37826
rect 30268 37772 30324 37774
rect 31164 39004 31220 39060
rect 31948 40572 32004 40628
rect 31948 40236 32004 40292
rect 31724 40012 31780 40068
rect 31724 39676 31780 39732
rect 31612 39618 31668 39620
rect 31612 39566 31614 39618
rect 31614 39566 31666 39618
rect 31666 39566 31668 39618
rect 31612 39564 31668 39566
rect 32284 40572 32340 40628
rect 32396 40402 32452 40404
rect 32396 40350 32398 40402
rect 32398 40350 32450 40402
rect 32450 40350 32452 40402
rect 32396 40348 32452 40350
rect 33404 42700 33460 42756
rect 33068 42476 33124 42532
rect 33180 42252 33236 42308
rect 33404 42364 33460 42420
rect 33068 41692 33124 41748
rect 33180 41804 33236 41860
rect 32732 41356 32788 41412
rect 33292 41410 33348 41412
rect 33292 41358 33294 41410
rect 33294 41358 33346 41410
rect 33346 41358 33348 41410
rect 33292 41356 33348 41358
rect 34860 44156 34916 44212
rect 34188 44098 34244 44100
rect 34188 44046 34190 44098
rect 34190 44046 34242 44098
rect 34242 44046 34244 44098
rect 34188 44044 34244 44046
rect 33964 43932 34020 43988
rect 35196 43426 35252 43428
rect 35196 43374 35198 43426
rect 35198 43374 35250 43426
rect 35250 43374 35252 43426
rect 35196 43372 35252 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34860 42924 34916 42980
rect 34188 42700 34244 42756
rect 33852 42364 33908 42420
rect 33852 41132 33908 41188
rect 32284 39788 32340 39844
rect 31948 39394 32004 39396
rect 31948 39342 31950 39394
rect 31950 39342 32002 39394
rect 32002 39342 32004 39394
rect 31948 39340 32004 39342
rect 31052 38332 31108 38388
rect 30716 38220 30772 38276
rect 30940 37436 30996 37492
rect 29820 36092 29876 36148
rect 29932 36316 29988 36372
rect 30268 36370 30324 36372
rect 30268 36318 30270 36370
rect 30270 36318 30322 36370
rect 30322 36318 30324 36370
rect 30268 36316 30324 36318
rect 30156 36258 30212 36260
rect 30156 36206 30158 36258
rect 30158 36206 30210 36258
rect 30210 36206 30212 36258
rect 30156 36204 30212 36206
rect 30044 35868 30100 35924
rect 29932 35644 29988 35700
rect 29148 34412 29204 34468
rect 32172 39116 32228 39172
rect 31724 38946 31780 38948
rect 31724 38894 31726 38946
rect 31726 38894 31778 38946
rect 31778 38894 31780 38946
rect 31724 38892 31780 38894
rect 31724 38668 31780 38724
rect 31948 38108 32004 38164
rect 31836 38050 31892 38052
rect 31836 37998 31838 38050
rect 31838 37998 31890 38050
rect 31890 37998 31892 38050
rect 31836 37996 31892 37998
rect 32508 39676 32564 39732
rect 32508 38274 32564 38276
rect 32508 38222 32510 38274
rect 32510 38222 32562 38274
rect 32562 38222 32564 38274
rect 32508 38220 32564 38222
rect 32396 37772 32452 37828
rect 31948 37212 32004 37268
rect 30268 35308 30324 35364
rect 31836 36876 31892 36932
rect 32172 36876 32228 36932
rect 30940 36316 30996 36372
rect 31388 35980 31444 36036
rect 31276 35922 31332 35924
rect 31276 35870 31278 35922
rect 31278 35870 31330 35922
rect 31330 35870 31332 35922
rect 31276 35868 31332 35870
rect 31164 35810 31220 35812
rect 31164 35758 31166 35810
rect 31166 35758 31218 35810
rect 31218 35758 31220 35810
rect 31164 35756 31220 35758
rect 30940 35698 30996 35700
rect 30940 35646 30942 35698
rect 30942 35646 30994 35698
rect 30994 35646 30996 35698
rect 30940 35644 30996 35646
rect 30716 35308 30772 35364
rect 29260 33964 29316 34020
rect 29148 33516 29204 33572
rect 30044 33458 30100 33460
rect 30044 33406 30046 33458
rect 30046 33406 30098 33458
rect 30098 33406 30100 33458
rect 30044 33404 30100 33406
rect 30492 33740 30548 33796
rect 30604 33628 30660 33684
rect 30156 33346 30212 33348
rect 30156 33294 30158 33346
rect 30158 33294 30210 33346
rect 30210 33294 30212 33346
rect 30156 33292 30212 33294
rect 29708 33234 29764 33236
rect 29708 33182 29710 33234
rect 29710 33182 29762 33234
rect 29762 33182 29764 33234
rect 29708 33180 29764 33182
rect 29932 33122 29988 33124
rect 29932 33070 29934 33122
rect 29934 33070 29986 33122
rect 29986 33070 29988 33122
rect 29932 33068 29988 33070
rect 30492 32844 30548 32900
rect 29596 32674 29652 32676
rect 29596 32622 29598 32674
rect 29598 32622 29650 32674
rect 29650 32622 29652 32674
rect 29596 32620 29652 32622
rect 28588 31666 28644 31668
rect 28588 31614 28590 31666
rect 28590 31614 28642 31666
rect 28642 31614 28644 31666
rect 28588 31612 28644 31614
rect 28476 31276 28532 31332
rect 29484 32396 29540 32452
rect 29036 31724 29092 31780
rect 28812 31052 28868 31108
rect 31164 33516 31220 33572
rect 31052 33292 31108 33348
rect 29708 31388 29764 31444
rect 30156 32338 30212 32340
rect 30156 32286 30158 32338
rect 30158 32286 30210 32338
rect 30210 32286 30212 32338
rect 30156 32284 30212 32286
rect 27804 30044 27860 30100
rect 27692 29986 27748 29988
rect 27692 29934 27694 29986
rect 27694 29934 27746 29986
rect 27746 29934 27748 29986
rect 27692 29932 27748 29934
rect 27580 29820 27636 29876
rect 27132 29372 27188 29428
rect 28140 28700 28196 28756
rect 27804 28642 27860 28644
rect 27804 28590 27806 28642
rect 27806 28590 27858 28642
rect 27858 28590 27860 28642
rect 27804 28588 27860 28590
rect 27244 28082 27300 28084
rect 27244 28030 27246 28082
rect 27246 28030 27298 28082
rect 27298 28030 27300 28082
rect 27244 28028 27300 28030
rect 27580 27298 27636 27300
rect 27580 27246 27582 27298
rect 27582 27246 27634 27298
rect 27634 27246 27636 27298
rect 27580 27244 27636 27246
rect 27692 27020 27748 27076
rect 27244 24892 27300 24948
rect 26908 23436 26964 23492
rect 26460 21756 26516 21812
rect 26124 21644 26180 21700
rect 25564 21586 25620 21588
rect 25564 21534 25566 21586
rect 25566 21534 25618 21586
rect 25618 21534 25620 21586
rect 25564 21532 25620 21534
rect 26908 21532 26964 21588
rect 25788 21420 25844 21476
rect 26236 21474 26292 21476
rect 26236 21422 26238 21474
rect 26238 21422 26290 21474
rect 26290 21422 26292 21474
rect 26236 21420 26292 21422
rect 26572 21308 26628 21364
rect 26348 21196 26404 21252
rect 25340 20076 25396 20132
rect 23324 17554 23380 17556
rect 23324 17502 23326 17554
rect 23326 17502 23378 17554
rect 23378 17502 23380 17554
rect 23324 17500 23380 17502
rect 22540 15538 22596 15540
rect 22540 15486 22542 15538
rect 22542 15486 22594 15538
rect 22594 15486 22596 15538
rect 22540 15484 22596 15486
rect 20524 10668 20580 10724
rect 18396 10610 18452 10612
rect 18396 10558 18398 10610
rect 18398 10558 18450 10610
rect 18450 10558 18452 10610
rect 18396 10556 18452 10558
rect 18172 9602 18228 9604
rect 18172 9550 18174 9602
rect 18174 9550 18226 9602
rect 18226 9550 18228 9602
rect 18172 9548 18228 9550
rect 16716 9100 16772 9156
rect 16604 7868 16660 7924
rect 16828 8092 16884 8148
rect 18172 8930 18228 8932
rect 18172 8878 18174 8930
rect 18174 8878 18226 8930
rect 18226 8878 18228 8930
rect 18172 8876 18228 8878
rect 17388 7980 17444 8036
rect 17948 8204 18004 8260
rect 16828 7586 16884 7588
rect 16828 7534 16830 7586
rect 16830 7534 16882 7586
rect 16882 7534 16884 7586
rect 16828 7532 16884 7534
rect 17388 7474 17444 7476
rect 17388 7422 17390 7474
rect 17390 7422 17442 7474
rect 17442 7422 17444 7474
rect 17388 7420 17444 7422
rect 16716 6412 16772 6468
rect 16380 6300 16436 6356
rect 16604 5906 16660 5908
rect 16604 5854 16606 5906
rect 16606 5854 16658 5906
rect 16658 5854 16660 5906
rect 16604 5852 16660 5854
rect 16492 5794 16548 5796
rect 16492 5742 16494 5794
rect 16494 5742 16546 5794
rect 16546 5742 16548 5794
rect 16492 5740 16548 5742
rect 16156 5404 16212 5460
rect 16940 6412 16996 6468
rect 17724 6188 17780 6244
rect 16940 5964 16996 6020
rect 16828 5516 16884 5572
rect 14588 3724 14644 3780
rect 13692 3388 13748 3444
rect 17052 5516 17108 5572
rect 16044 3500 16100 3556
rect 17276 5516 17332 5572
rect 17164 5292 17220 5348
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19740 8258 19796 8260
rect 19740 8206 19742 8258
rect 19742 8206 19794 8258
rect 19794 8206 19796 8258
rect 19740 8204 19796 8206
rect 20188 8034 20244 8036
rect 20188 7982 20190 8034
rect 20190 7982 20242 8034
rect 20242 7982 20244 8034
rect 20188 7980 20244 7982
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 18396 7644 18452 7700
rect 19852 7644 19908 7700
rect 19628 7420 19684 7476
rect 18284 7196 18340 7252
rect 18060 6130 18116 6132
rect 18060 6078 18062 6130
rect 18062 6078 18114 6130
rect 18114 6078 18116 6130
rect 18060 6076 18116 6078
rect 18396 5906 18452 5908
rect 18396 5854 18398 5906
rect 18398 5854 18450 5906
rect 18450 5854 18452 5906
rect 18396 5852 18452 5854
rect 19068 7196 19124 7252
rect 18620 6188 18676 6244
rect 18620 5404 18676 5460
rect 18508 5292 18564 5348
rect 18060 5068 18116 5124
rect 18956 5516 19012 5572
rect 18844 5292 18900 5348
rect 20748 8316 20804 8372
rect 21084 12460 21140 12516
rect 21196 11788 21252 11844
rect 21644 13804 21700 13860
rect 21308 9884 21364 9940
rect 22092 14364 22148 14420
rect 22204 14306 22260 14308
rect 22204 14254 22206 14306
rect 22206 14254 22258 14306
rect 22258 14254 22260 14306
rect 22204 14252 22260 14254
rect 22092 13468 22148 13524
rect 22540 14306 22596 14308
rect 22540 14254 22542 14306
rect 22542 14254 22594 14306
rect 22594 14254 22596 14306
rect 22540 14252 22596 14254
rect 22540 13468 22596 13524
rect 22428 12460 22484 12516
rect 21868 11788 21924 11844
rect 21420 9212 21476 9268
rect 20860 8204 20916 8260
rect 21420 8204 21476 8260
rect 20748 8092 20804 8148
rect 20412 7532 20468 7588
rect 20972 8092 21028 8148
rect 19964 6466 20020 6468
rect 19964 6414 19966 6466
rect 19966 6414 20018 6466
rect 20018 6414 20020 6466
rect 19964 6412 20020 6414
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19628 6076 19684 6132
rect 19852 5122 19908 5124
rect 19852 5070 19854 5122
rect 19854 5070 19906 5122
rect 19906 5070 19908 5122
rect 19852 5068 19908 5070
rect 20748 7474 20804 7476
rect 20748 7422 20750 7474
rect 20750 7422 20802 7474
rect 20802 7422 20804 7474
rect 20748 7420 20804 7422
rect 21756 11340 21812 11396
rect 21644 10610 21700 10612
rect 21644 10558 21646 10610
rect 21646 10558 21698 10610
rect 21698 10558 21700 10610
rect 21644 10556 21700 10558
rect 21532 7868 21588 7924
rect 23100 16044 23156 16100
rect 24332 18450 24388 18452
rect 24332 18398 24334 18450
rect 24334 18398 24386 18450
rect 24386 18398 24388 18450
rect 24332 18396 24388 18398
rect 24556 19852 24612 19908
rect 24220 18172 24276 18228
rect 23884 16098 23940 16100
rect 23884 16046 23886 16098
rect 23886 16046 23938 16098
rect 23938 16046 23940 16098
rect 23884 16044 23940 16046
rect 24108 15260 24164 15316
rect 23436 15036 23492 15092
rect 23772 15148 23828 15204
rect 25340 19346 25396 19348
rect 25340 19294 25342 19346
rect 25342 19294 25394 19346
rect 25394 19294 25396 19346
rect 25340 19292 25396 19294
rect 26012 20076 26068 20132
rect 24668 17724 24724 17780
rect 24668 17106 24724 17108
rect 24668 17054 24670 17106
rect 24670 17054 24722 17106
rect 24722 17054 24724 17106
rect 24668 17052 24724 17054
rect 27580 23548 27636 23604
rect 27468 23436 27524 23492
rect 27580 23378 27636 23380
rect 27580 23326 27582 23378
rect 27582 23326 27634 23378
rect 27634 23326 27636 23378
rect 27580 23324 27636 23326
rect 27244 23154 27300 23156
rect 27244 23102 27246 23154
rect 27246 23102 27298 23154
rect 27298 23102 27300 23154
rect 27244 23100 27300 23102
rect 28140 28140 28196 28196
rect 28476 28754 28532 28756
rect 28476 28702 28478 28754
rect 28478 28702 28530 28754
rect 28530 28702 28532 28754
rect 28476 28700 28532 28702
rect 28476 28140 28532 28196
rect 28364 28028 28420 28084
rect 28700 27468 28756 27524
rect 28364 27074 28420 27076
rect 28364 27022 28366 27074
rect 28366 27022 28418 27074
rect 28418 27022 28420 27074
rect 28364 27020 28420 27022
rect 28476 27244 28532 27300
rect 28364 24892 28420 24948
rect 28140 23378 28196 23380
rect 28140 23326 28142 23378
rect 28142 23326 28194 23378
rect 28194 23326 28196 23378
rect 28140 23324 28196 23326
rect 28700 23436 28756 23492
rect 29260 30268 29316 30324
rect 29148 29148 29204 29204
rect 29596 30098 29652 30100
rect 29596 30046 29598 30098
rect 29598 30046 29650 30098
rect 29650 30046 29652 30098
rect 29596 30044 29652 30046
rect 29260 28588 29316 28644
rect 29484 29820 29540 29876
rect 29596 28700 29652 28756
rect 29932 29932 29988 29988
rect 29484 28588 29540 28644
rect 29148 28364 29204 28420
rect 28924 27916 28980 27972
rect 29148 27692 29204 27748
rect 29260 28028 29316 28084
rect 29932 28364 29988 28420
rect 29260 27244 29316 27300
rect 29484 27692 29540 27748
rect 28924 25564 28980 25620
rect 29148 25282 29204 25284
rect 29148 25230 29150 25282
rect 29150 25230 29202 25282
rect 29202 25230 29204 25282
rect 29148 25228 29204 25230
rect 30940 32284 30996 32340
rect 31164 33234 31220 33236
rect 31164 33182 31166 33234
rect 31166 33182 31218 33234
rect 31218 33182 31220 33234
rect 31164 33180 31220 33182
rect 31500 33628 31556 33684
rect 31612 33292 31668 33348
rect 32060 36092 32116 36148
rect 34188 40962 34244 40964
rect 34188 40910 34190 40962
rect 34190 40910 34242 40962
rect 34242 40910 34244 40962
rect 34188 40908 34244 40910
rect 34636 42700 34692 42756
rect 34412 42642 34468 42644
rect 34412 42590 34414 42642
rect 34414 42590 34466 42642
rect 34466 42590 34468 42642
rect 34412 42588 34468 42590
rect 33180 40626 33236 40628
rect 33180 40574 33182 40626
rect 33182 40574 33234 40626
rect 33234 40574 33236 40626
rect 33180 40572 33236 40574
rect 33180 40348 33236 40404
rect 32956 39730 33012 39732
rect 32956 39678 32958 39730
rect 32958 39678 33010 39730
rect 33010 39678 33012 39730
rect 32956 39676 33012 39678
rect 32732 39452 32788 39508
rect 33068 39618 33124 39620
rect 33068 39566 33070 39618
rect 33070 39566 33122 39618
rect 33122 39566 33124 39618
rect 33068 39564 33124 39566
rect 33180 39506 33236 39508
rect 33180 39454 33182 39506
rect 33182 39454 33234 39506
rect 33234 39454 33236 39506
rect 33180 39452 33236 39454
rect 32732 38108 32788 38164
rect 32620 37436 32676 37492
rect 32396 37154 32452 37156
rect 32396 37102 32398 37154
rect 32398 37102 32450 37154
rect 32450 37102 32452 37154
rect 32396 37100 32452 37102
rect 32508 36540 32564 36596
rect 32172 35532 32228 35588
rect 31836 34130 31892 34132
rect 31836 34078 31838 34130
rect 31838 34078 31890 34130
rect 31890 34078 31892 34130
rect 31836 34076 31892 34078
rect 32060 35196 32116 35252
rect 32060 33852 32116 33908
rect 32620 35980 32676 36036
rect 32396 35196 32452 35252
rect 32508 35420 32564 35476
rect 32284 34188 32340 34244
rect 31948 33516 32004 33572
rect 31276 32786 31332 32788
rect 31276 32734 31278 32786
rect 31278 32734 31330 32786
rect 31330 32734 31332 32786
rect 31276 32732 31332 32734
rect 32396 34076 32452 34132
rect 32396 32732 32452 32788
rect 31164 32620 31220 32676
rect 31052 32508 31108 32564
rect 30380 31836 30436 31892
rect 30156 30828 30212 30884
rect 30716 30828 30772 30884
rect 30828 31388 30884 31444
rect 30380 30268 30436 30324
rect 31388 30156 31444 30212
rect 30268 30098 30324 30100
rect 30268 30046 30270 30098
rect 30270 30046 30322 30098
rect 30322 30046 30324 30098
rect 30268 30044 30324 30046
rect 30156 29820 30212 29876
rect 30156 29484 30212 29540
rect 31276 29986 31332 29988
rect 31276 29934 31278 29986
rect 31278 29934 31330 29986
rect 31330 29934 31332 29986
rect 31276 29932 31332 29934
rect 31052 29820 31108 29876
rect 30716 29596 30772 29652
rect 30492 29484 30548 29540
rect 30380 27298 30436 27300
rect 30380 27246 30382 27298
rect 30382 27246 30434 27298
rect 30434 27246 30436 27298
rect 30380 27244 30436 27246
rect 31276 29596 31332 29652
rect 31836 32620 31892 32676
rect 31612 32508 31668 32564
rect 32172 32396 32228 32452
rect 32284 32508 32340 32564
rect 32956 36988 33012 37044
rect 33292 37548 33348 37604
rect 33068 36428 33124 36484
rect 33180 37100 33236 37156
rect 33292 35980 33348 36036
rect 33516 39676 33572 39732
rect 33628 39506 33684 39508
rect 33628 39454 33630 39506
rect 33630 39454 33682 39506
rect 33682 39454 33684 39506
rect 33628 39452 33684 39454
rect 33628 39058 33684 39060
rect 33628 39006 33630 39058
rect 33630 39006 33682 39058
rect 33682 39006 33684 39058
rect 33628 39004 33684 39006
rect 33516 37826 33572 37828
rect 33516 37774 33518 37826
rect 33518 37774 33570 37826
rect 33570 37774 33572 37826
rect 33516 37772 33572 37774
rect 34748 42476 34804 42532
rect 35868 44044 35924 44100
rect 35644 43372 35700 43428
rect 37100 44210 37156 44212
rect 37100 44158 37102 44210
rect 37102 44158 37154 44210
rect 37154 44158 37156 44210
rect 37100 44156 37156 44158
rect 39228 43932 39284 43988
rect 36428 43820 36484 43876
rect 37324 43820 37380 43876
rect 36316 43036 36372 43092
rect 35532 42252 35588 42308
rect 35196 41858 35252 41860
rect 35196 41806 35198 41858
rect 35198 41806 35250 41858
rect 35250 41806 35252 41858
rect 35196 41804 35252 41806
rect 34972 41692 35028 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35644 42028 35700 42084
rect 34300 40402 34356 40404
rect 34300 40350 34302 40402
rect 34302 40350 34354 40402
rect 34354 40350 34356 40402
rect 34300 40348 34356 40350
rect 33964 39900 34020 39956
rect 33852 39228 33908 39284
rect 34188 39116 34244 39172
rect 33852 38834 33908 38836
rect 33852 38782 33854 38834
rect 33854 38782 33906 38834
rect 33906 38782 33908 38834
rect 33852 38780 33908 38782
rect 34412 38834 34468 38836
rect 34412 38782 34414 38834
rect 34414 38782 34466 38834
rect 34466 38782 34468 38834
rect 34412 38780 34468 38782
rect 34636 38834 34692 38836
rect 34636 38782 34638 38834
rect 34638 38782 34690 38834
rect 34690 38782 34692 38834
rect 34636 38780 34692 38782
rect 34300 38668 34356 38724
rect 34636 38444 34692 38500
rect 33964 37938 34020 37940
rect 33964 37886 33966 37938
rect 33966 37886 34018 37938
rect 34018 37886 34020 37938
rect 33964 37884 34020 37886
rect 33852 37548 33908 37604
rect 33628 36594 33684 36596
rect 33628 36542 33630 36594
rect 33630 36542 33682 36594
rect 33682 36542 33684 36594
rect 33628 36540 33684 36542
rect 33516 36092 33572 36148
rect 33068 35308 33124 35364
rect 33516 34242 33572 34244
rect 33516 34190 33518 34242
rect 33518 34190 33570 34242
rect 33570 34190 33572 34242
rect 33516 34188 33572 34190
rect 32844 34076 32900 34132
rect 33628 34130 33684 34132
rect 33628 34078 33630 34130
rect 33630 34078 33682 34130
rect 33682 34078 33684 34130
rect 33628 34076 33684 34078
rect 33180 33516 33236 33572
rect 32620 32396 32676 32452
rect 31724 32060 31780 32116
rect 31724 30882 31780 30884
rect 31724 30830 31726 30882
rect 31726 30830 31778 30882
rect 31778 30830 31780 30882
rect 31724 30828 31780 30830
rect 33852 36540 33908 36596
rect 34076 35532 34132 35588
rect 34524 36988 34580 37044
rect 34188 35420 34244 35476
rect 34076 34242 34132 34244
rect 34076 34190 34078 34242
rect 34078 34190 34130 34242
rect 34130 34190 34132 34242
rect 34076 34188 34132 34190
rect 34188 33964 34244 34020
rect 34412 33628 34468 33684
rect 34300 33516 34356 33572
rect 34188 33404 34244 33460
rect 33404 32844 33460 32900
rect 33404 31948 33460 32004
rect 31612 29484 31668 29540
rect 30828 28812 30884 28868
rect 30940 28588 30996 28644
rect 30268 26796 30324 26852
rect 30268 26402 30324 26404
rect 30268 26350 30270 26402
rect 30270 26350 30322 26402
rect 30322 26350 30324 26402
rect 30268 26348 30324 26350
rect 29484 24162 29540 24164
rect 29484 24110 29486 24162
rect 29486 24110 29538 24162
rect 29538 24110 29540 24162
rect 29484 24108 29540 24110
rect 29708 24108 29764 24164
rect 30828 26348 30884 26404
rect 31164 26012 31220 26068
rect 30716 25618 30772 25620
rect 30716 25566 30718 25618
rect 30718 25566 30770 25618
rect 30770 25566 30772 25618
rect 30716 25564 30772 25566
rect 28812 23324 28868 23380
rect 28588 23212 28644 23268
rect 28476 23100 28532 23156
rect 28364 22876 28420 22932
rect 27244 21756 27300 21812
rect 27244 20690 27300 20692
rect 27244 20638 27246 20690
rect 27246 20638 27298 20690
rect 27298 20638 27300 20690
rect 27244 20636 27300 20638
rect 26348 19292 26404 19348
rect 26012 18172 26068 18228
rect 26796 20018 26852 20020
rect 26796 19966 26798 20018
rect 26798 19966 26850 20018
rect 26850 19966 26852 20018
rect 26796 19964 26852 19966
rect 26684 18508 26740 18564
rect 25452 17052 25508 17108
rect 26348 17052 26404 17108
rect 24332 16828 24388 16884
rect 25452 16882 25508 16884
rect 25452 16830 25454 16882
rect 25454 16830 25506 16882
rect 25506 16830 25508 16882
rect 25452 16828 25508 16830
rect 28252 20524 28308 20580
rect 28252 20188 28308 20244
rect 27356 20130 27412 20132
rect 27356 20078 27358 20130
rect 27358 20078 27410 20130
rect 27410 20078 27412 20130
rect 27356 20076 27412 20078
rect 27580 20018 27636 20020
rect 27580 19966 27582 20018
rect 27582 19966 27634 20018
rect 27634 19966 27636 20018
rect 27580 19964 27636 19966
rect 27692 19906 27748 19908
rect 27692 19854 27694 19906
rect 27694 19854 27746 19906
rect 27746 19854 27748 19906
rect 27692 19852 27748 19854
rect 27020 19740 27076 19796
rect 28252 18508 28308 18564
rect 27916 18284 27972 18340
rect 26908 17052 26964 17108
rect 27692 17106 27748 17108
rect 27692 17054 27694 17106
rect 27694 17054 27746 17106
rect 27746 17054 27748 17106
rect 27692 17052 27748 17054
rect 26124 16156 26180 16212
rect 26796 16210 26852 16212
rect 26796 16158 26798 16210
rect 26798 16158 26850 16210
rect 26850 16158 26852 16210
rect 26796 16156 26852 16158
rect 25340 15314 25396 15316
rect 25340 15262 25342 15314
rect 25342 15262 25394 15314
rect 25394 15262 25396 15314
rect 25340 15260 25396 15262
rect 25228 15202 25284 15204
rect 25228 15150 25230 15202
rect 25230 15150 25282 15202
rect 25282 15150 25284 15202
rect 25228 15148 25284 15150
rect 23548 13916 23604 13972
rect 24332 14252 24388 14308
rect 22988 13746 23044 13748
rect 22988 13694 22990 13746
rect 22990 13694 23042 13746
rect 23042 13694 23044 13746
rect 22988 13692 23044 13694
rect 23660 13858 23716 13860
rect 23660 13806 23662 13858
rect 23662 13806 23714 13858
rect 23714 13806 23716 13858
rect 23660 13804 23716 13806
rect 22876 12236 22932 12292
rect 22876 11788 22932 11844
rect 22764 9548 22820 9604
rect 22204 9324 22260 9380
rect 21980 8316 22036 8372
rect 21756 8146 21812 8148
rect 21756 8094 21758 8146
rect 21758 8094 21810 8146
rect 21810 8094 21812 8146
rect 21756 8092 21812 8094
rect 22316 7868 22372 7924
rect 21420 7084 21476 7140
rect 22204 7586 22260 7588
rect 22204 7534 22206 7586
rect 22206 7534 22258 7586
rect 22258 7534 22260 7586
rect 22204 7532 22260 7534
rect 21644 7362 21700 7364
rect 21644 7310 21646 7362
rect 21646 7310 21698 7362
rect 21698 7310 21700 7362
rect 21644 7308 21700 7310
rect 20972 6748 21028 6804
rect 20524 6076 20580 6132
rect 20748 6466 20804 6468
rect 20748 6414 20750 6466
rect 20750 6414 20802 6466
rect 20802 6414 20804 6466
rect 20748 6412 20804 6414
rect 20748 5628 20804 5684
rect 20636 5516 20692 5572
rect 20860 5292 20916 5348
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 18732 4396 18788 4452
rect 18732 4226 18788 4228
rect 18732 4174 18734 4226
rect 18734 4174 18786 4226
rect 18786 4174 18788 4226
rect 18732 4172 18788 4174
rect 17612 3554 17668 3556
rect 17612 3502 17614 3554
rect 17614 3502 17666 3554
rect 17666 3502 17668 3554
rect 17612 3500 17668 3502
rect 20076 3612 20132 3668
rect 21644 6636 21700 6692
rect 21532 6578 21588 6580
rect 21532 6526 21534 6578
rect 21534 6526 21586 6578
rect 21586 6526 21588 6578
rect 21532 6524 21588 6526
rect 21308 6076 21364 6132
rect 21308 5068 21364 5124
rect 21532 4396 21588 4452
rect 21868 6412 21924 6468
rect 23996 12290 24052 12292
rect 23996 12238 23998 12290
rect 23998 12238 24050 12290
rect 24050 12238 24052 12290
rect 23996 12236 24052 12238
rect 24108 12348 24164 12404
rect 23884 12178 23940 12180
rect 23884 12126 23886 12178
rect 23886 12126 23938 12178
rect 23938 12126 23940 12178
rect 23884 12124 23940 12126
rect 23660 12012 23716 12068
rect 23548 11340 23604 11396
rect 24556 13746 24612 13748
rect 24556 13694 24558 13746
rect 24558 13694 24610 13746
rect 24610 13694 24612 13746
rect 24556 13692 24612 13694
rect 24444 13522 24500 13524
rect 24444 13470 24446 13522
rect 24446 13470 24498 13522
rect 24498 13470 24500 13522
rect 24444 13468 24500 13470
rect 24444 11900 24500 11956
rect 25228 13522 25284 13524
rect 25228 13470 25230 13522
rect 25230 13470 25282 13522
rect 25282 13470 25284 13522
rect 25228 13468 25284 13470
rect 25564 15202 25620 15204
rect 25564 15150 25566 15202
rect 25566 15150 25618 15202
rect 25618 15150 25620 15202
rect 25564 15148 25620 15150
rect 26684 15314 26740 15316
rect 26684 15262 26686 15314
rect 26686 15262 26738 15314
rect 26738 15262 26740 15314
rect 26684 15260 26740 15262
rect 26796 15148 26852 15204
rect 26236 15036 26292 15092
rect 26908 14700 26964 14756
rect 27580 16940 27636 16996
rect 26348 14028 26404 14084
rect 26460 13692 26516 13748
rect 26572 14028 26628 14084
rect 26796 13858 26852 13860
rect 26796 13806 26798 13858
rect 26798 13806 26850 13858
rect 26850 13806 26852 13858
rect 26796 13804 26852 13806
rect 27244 14700 27300 14756
rect 27356 15932 27412 15988
rect 28140 16994 28196 16996
rect 28140 16942 28142 16994
rect 28142 16942 28194 16994
rect 28194 16942 28196 16994
rect 28140 16940 28196 16942
rect 28588 21420 28644 21476
rect 28476 20578 28532 20580
rect 28476 20526 28478 20578
rect 28478 20526 28530 20578
rect 28530 20526 28532 20578
rect 28476 20524 28532 20526
rect 29036 21308 29092 21364
rect 28588 20188 28644 20244
rect 29148 20076 29204 20132
rect 28700 19740 28756 19796
rect 28588 17554 28644 17556
rect 28588 17502 28590 17554
rect 28590 17502 28642 17554
rect 28642 17502 28644 17554
rect 28588 17500 28644 17502
rect 28364 16492 28420 16548
rect 27692 16156 27748 16212
rect 28588 16210 28644 16212
rect 28588 16158 28590 16210
rect 28590 16158 28642 16210
rect 28642 16158 28644 16210
rect 28588 16156 28644 16158
rect 27468 15484 27524 15540
rect 27580 15596 27636 15652
rect 27804 15986 27860 15988
rect 27804 15934 27806 15986
rect 27806 15934 27858 15986
rect 27858 15934 27860 15986
rect 27804 15932 27860 15934
rect 27916 15426 27972 15428
rect 27916 15374 27918 15426
rect 27918 15374 27970 15426
rect 27970 15374 27972 15426
rect 27916 15372 27972 15374
rect 27356 15036 27412 15092
rect 27356 14588 27412 14644
rect 27132 14476 27188 14532
rect 28028 15314 28084 15316
rect 28028 15262 28030 15314
rect 28030 15262 28082 15314
rect 28082 15262 28084 15314
rect 28028 15260 28084 15262
rect 28476 15596 28532 15652
rect 28364 15260 28420 15316
rect 27692 15036 27748 15092
rect 28364 15036 28420 15092
rect 27692 14418 27748 14420
rect 27692 14366 27694 14418
rect 27694 14366 27746 14418
rect 27746 14366 27748 14418
rect 27692 14364 27748 14366
rect 28028 14028 28084 14084
rect 25788 13634 25844 13636
rect 25788 13582 25790 13634
rect 25790 13582 25842 13634
rect 25842 13582 25844 13634
rect 25788 13580 25844 13582
rect 26572 13580 26628 13636
rect 26460 13468 26516 13524
rect 25564 12348 25620 12404
rect 26460 12236 26516 12292
rect 25788 12178 25844 12180
rect 25788 12126 25790 12178
rect 25790 12126 25842 12178
rect 25842 12126 25844 12178
rect 25788 12124 25844 12126
rect 26124 12066 26180 12068
rect 26124 12014 26126 12066
rect 26126 12014 26178 12066
rect 26178 12014 26180 12066
rect 26124 12012 26180 12014
rect 28028 13858 28084 13860
rect 28028 13806 28030 13858
rect 28030 13806 28082 13858
rect 28082 13806 28084 13858
rect 28028 13804 28084 13806
rect 27692 13020 27748 13076
rect 27468 12684 27524 12740
rect 26908 12178 26964 12180
rect 26908 12126 26910 12178
rect 26910 12126 26962 12178
rect 26962 12126 26964 12178
rect 26908 12124 26964 12126
rect 26684 11900 26740 11956
rect 27244 12290 27300 12292
rect 27244 12238 27246 12290
rect 27246 12238 27298 12290
rect 27298 12238 27300 12290
rect 27244 12236 27300 12238
rect 27132 11900 27188 11956
rect 27244 11170 27300 11172
rect 27244 11118 27246 11170
rect 27246 11118 27298 11170
rect 27298 11118 27300 11170
rect 27244 11116 27300 11118
rect 27244 10892 27300 10948
rect 24220 9938 24276 9940
rect 24220 9886 24222 9938
rect 24222 9886 24274 9938
rect 24274 9886 24276 9938
rect 24220 9884 24276 9886
rect 23436 9602 23492 9604
rect 23436 9550 23438 9602
rect 23438 9550 23490 9602
rect 23490 9550 23492 9602
rect 23436 9548 23492 9550
rect 22876 8092 22932 8148
rect 23212 8034 23268 8036
rect 23212 7982 23214 8034
rect 23214 7982 23266 8034
rect 23266 7982 23268 8034
rect 23212 7980 23268 7982
rect 22876 7586 22932 7588
rect 22876 7534 22878 7586
rect 22878 7534 22930 7586
rect 22930 7534 22932 7586
rect 22876 7532 22932 7534
rect 22428 7420 22484 7476
rect 22652 7308 22708 7364
rect 23100 7196 23156 7252
rect 22764 5516 22820 5572
rect 23324 7196 23380 7252
rect 23436 6748 23492 6804
rect 24332 8988 24388 9044
rect 23660 8370 23716 8372
rect 23660 8318 23662 8370
rect 23662 8318 23714 8370
rect 23714 8318 23716 8370
rect 23660 8316 23716 8318
rect 23660 8092 23716 8148
rect 24108 8258 24164 8260
rect 24108 8206 24110 8258
rect 24110 8206 24162 8258
rect 24162 8206 24164 8258
rect 24108 8204 24164 8206
rect 25340 9996 25396 10052
rect 27132 9996 27188 10052
rect 25004 9884 25060 9940
rect 24780 9266 24836 9268
rect 24780 9214 24782 9266
rect 24782 9214 24834 9266
rect 24834 9214 24836 9266
rect 24780 9212 24836 9214
rect 24444 8764 24500 8820
rect 26572 9884 26628 9940
rect 25004 9100 25060 9156
rect 25228 9660 25284 9716
rect 26348 9714 26404 9716
rect 26348 9662 26350 9714
rect 26350 9662 26402 9714
rect 26402 9662 26404 9714
rect 26348 9660 26404 9662
rect 25228 9212 25284 9268
rect 27356 9212 27412 9268
rect 25564 9042 25620 9044
rect 25564 8990 25566 9042
rect 25566 8990 25618 9042
rect 25618 8990 25620 9042
rect 25564 8988 25620 8990
rect 25340 8146 25396 8148
rect 25340 8094 25342 8146
rect 25342 8094 25394 8146
rect 25394 8094 25396 8146
rect 25340 8092 25396 8094
rect 23548 6636 23604 6692
rect 23660 7084 23716 7140
rect 23212 5852 23268 5908
rect 22876 5180 22932 5236
rect 23660 5404 23716 5460
rect 21980 5068 22036 5124
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 23772 5068 23828 5124
rect 21868 3666 21924 3668
rect 21868 3614 21870 3666
rect 21870 3614 21922 3666
rect 21922 3614 21924 3666
rect 21868 3612 21924 3614
rect 24444 7868 24500 7924
rect 24332 7474 24388 7476
rect 24332 7422 24334 7474
rect 24334 7422 24386 7474
rect 24386 7422 24388 7474
rect 24332 7420 24388 7422
rect 24220 7362 24276 7364
rect 24220 7310 24222 7362
rect 24222 7310 24274 7362
rect 24274 7310 24276 7362
rect 24220 7308 24276 7310
rect 24780 6636 24836 6692
rect 24780 6076 24836 6132
rect 24220 5628 24276 5684
rect 24556 5404 24612 5460
rect 24220 5234 24276 5236
rect 24220 5182 24222 5234
rect 24222 5182 24274 5234
rect 24274 5182 24276 5234
rect 24220 5180 24276 5182
rect 25788 8092 25844 8148
rect 26012 9154 26068 9156
rect 26012 9102 26014 9154
rect 26014 9102 26066 9154
rect 26066 9102 26068 9154
rect 26012 9100 26068 9102
rect 26124 8092 26180 8148
rect 27580 12348 27636 12404
rect 27916 13244 27972 13300
rect 28028 12962 28084 12964
rect 28028 12910 28030 12962
rect 28030 12910 28082 12962
rect 28082 12910 28084 12962
rect 28028 12908 28084 12910
rect 28028 12178 28084 12180
rect 28028 12126 28030 12178
rect 28030 12126 28082 12178
rect 28082 12126 28084 12178
rect 28028 12124 28084 12126
rect 27692 10668 27748 10724
rect 28028 10668 28084 10724
rect 28700 15260 28756 15316
rect 29708 23154 29764 23156
rect 29708 23102 29710 23154
rect 29710 23102 29762 23154
rect 29762 23102 29764 23154
rect 29708 23100 29764 23102
rect 30044 22930 30100 22932
rect 30044 22878 30046 22930
rect 30046 22878 30098 22930
rect 30098 22878 30100 22930
rect 30044 22876 30100 22878
rect 29484 21586 29540 21588
rect 29484 21534 29486 21586
rect 29486 21534 29538 21586
rect 29538 21534 29540 21586
rect 29484 21532 29540 21534
rect 30380 22428 30436 22484
rect 30044 22370 30100 22372
rect 30044 22318 30046 22370
rect 30046 22318 30098 22370
rect 30098 22318 30100 22370
rect 30044 22316 30100 22318
rect 30044 21532 30100 21588
rect 29708 20802 29764 20804
rect 29708 20750 29710 20802
rect 29710 20750 29762 20802
rect 29762 20750 29764 20802
rect 29708 20748 29764 20750
rect 29596 20636 29652 20692
rect 29484 20412 29540 20468
rect 29372 20188 29428 20244
rect 29036 18844 29092 18900
rect 30828 23042 30884 23044
rect 30828 22990 30830 23042
rect 30830 22990 30882 23042
rect 30882 22990 30884 23042
rect 30828 22988 30884 22990
rect 30492 22316 30548 22372
rect 30380 21756 30436 21812
rect 31276 25788 31332 25844
rect 31164 25618 31220 25620
rect 31164 25566 31166 25618
rect 31166 25566 31218 25618
rect 31218 25566 31220 25618
rect 31164 25564 31220 25566
rect 31164 25394 31220 25396
rect 31164 25342 31166 25394
rect 31166 25342 31218 25394
rect 31218 25342 31220 25394
rect 31164 25340 31220 25342
rect 31164 24108 31220 24164
rect 31164 23154 31220 23156
rect 31164 23102 31166 23154
rect 31166 23102 31218 23154
rect 31218 23102 31220 23154
rect 31164 23100 31220 23102
rect 31612 28924 31668 28980
rect 31612 28140 31668 28196
rect 31500 25506 31556 25508
rect 31500 25454 31502 25506
rect 31502 25454 31554 25506
rect 31554 25454 31556 25506
rect 31500 25452 31556 25454
rect 32508 30828 32564 30884
rect 32172 29820 32228 29876
rect 32060 28754 32116 28756
rect 32060 28702 32062 28754
rect 32062 28702 32114 28754
rect 32114 28702 32116 28754
rect 32060 28700 32116 28702
rect 32284 29596 32340 29652
rect 32284 29426 32340 29428
rect 32284 29374 32286 29426
rect 32286 29374 32338 29426
rect 32338 29374 32340 29426
rect 32284 29372 32340 29374
rect 31836 25788 31892 25844
rect 32956 29820 33012 29876
rect 32620 29372 32676 29428
rect 32396 28530 32452 28532
rect 32396 28478 32398 28530
rect 32398 28478 32450 28530
rect 32450 28478 32452 28530
rect 32396 28476 32452 28478
rect 32508 28418 32564 28420
rect 32508 28366 32510 28418
rect 32510 28366 32562 28418
rect 32562 28366 32564 28418
rect 32508 28364 32564 28366
rect 32060 28140 32116 28196
rect 32284 28082 32340 28084
rect 32284 28030 32286 28082
rect 32286 28030 32338 28082
rect 32338 28030 32340 28082
rect 32284 28028 32340 28030
rect 32172 27746 32228 27748
rect 32172 27694 32174 27746
rect 32174 27694 32226 27746
rect 32226 27694 32228 27746
rect 32172 27692 32228 27694
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 34076 31948 34132 32004
rect 33404 30156 33460 30212
rect 33852 31276 33908 31332
rect 33404 29986 33460 29988
rect 33404 29934 33406 29986
rect 33406 29934 33458 29986
rect 33458 29934 33460 29986
rect 33404 29932 33460 29934
rect 33180 29650 33236 29652
rect 33180 29598 33182 29650
rect 33182 29598 33234 29650
rect 33234 29598 33236 29650
rect 33180 29596 33236 29598
rect 33404 29650 33460 29652
rect 33404 29598 33406 29650
rect 33406 29598 33458 29650
rect 33458 29598 33460 29650
rect 33404 29596 33460 29598
rect 33292 29426 33348 29428
rect 33292 29374 33294 29426
rect 33294 29374 33346 29426
rect 33346 29374 33348 29426
rect 33292 29372 33348 29374
rect 33180 28754 33236 28756
rect 33180 28702 33182 28754
rect 33182 28702 33234 28754
rect 33234 28702 33236 28754
rect 33180 28700 33236 28702
rect 33292 28252 33348 28308
rect 33404 28588 33460 28644
rect 33628 29372 33684 29428
rect 34300 33180 34356 33236
rect 34636 36258 34692 36260
rect 34636 36206 34638 36258
rect 34638 36206 34690 36258
rect 34690 36206 34692 36258
rect 34636 36204 34692 36206
rect 35196 40796 35252 40852
rect 35084 40572 35140 40628
rect 35532 40514 35588 40516
rect 35532 40462 35534 40514
rect 35534 40462 35586 40514
rect 35586 40462 35588 40514
rect 35532 40460 35588 40462
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36092 42754 36148 42756
rect 36092 42702 36094 42754
rect 36094 42702 36146 42754
rect 36146 42702 36148 42754
rect 36092 42700 36148 42702
rect 35980 41244 36036 41300
rect 35868 40124 35924 40180
rect 35756 39618 35812 39620
rect 35756 39566 35758 39618
rect 35758 39566 35810 39618
rect 35810 39566 35812 39618
rect 35756 39564 35812 39566
rect 35084 39340 35140 39396
rect 35868 39452 35924 39508
rect 34972 39116 35028 39172
rect 34972 38834 35028 38836
rect 34972 38782 34974 38834
rect 34974 38782 35026 38834
rect 35026 38782 35028 38834
rect 34972 38780 35028 38782
rect 36316 42364 36372 42420
rect 36204 42028 36260 42084
rect 36428 41804 36484 41860
rect 37100 43426 37156 43428
rect 37100 43374 37102 43426
rect 37102 43374 37154 43426
rect 37154 43374 37156 43426
rect 37100 43372 37156 43374
rect 36652 42364 36708 42420
rect 37100 41970 37156 41972
rect 37100 41918 37102 41970
rect 37102 41918 37154 41970
rect 37154 41918 37156 41970
rect 37100 41916 37156 41918
rect 36988 41858 37044 41860
rect 36988 41806 36990 41858
rect 36990 41806 37042 41858
rect 37042 41806 37044 41858
rect 36988 41804 37044 41806
rect 39116 43484 39172 43540
rect 37996 43372 38052 43428
rect 37548 42364 37604 42420
rect 36540 41244 36596 41300
rect 36316 40460 36372 40516
rect 36764 40460 36820 40516
rect 36204 40348 36260 40404
rect 36876 40290 36932 40292
rect 36876 40238 36878 40290
rect 36878 40238 36930 40290
rect 36930 40238 36932 40290
rect 36876 40236 36932 40238
rect 36092 39564 36148 39620
rect 35084 38668 35140 38724
rect 34972 38332 35028 38388
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35980 38050 36036 38052
rect 35980 37998 35982 38050
rect 35982 37998 36034 38050
rect 36034 37998 36036 38050
rect 35980 37996 36036 37998
rect 37212 41298 37268 41300
rect 37212 41246 37214 41298
rect 37214 41246 37266 41298
rect 37266 41246 37268 41298
rect 37212 41244 37268 41246
rect 38444 42978 38500 42980
rect 38444 42926 38446 42978
rect 38446 42926 38498 42978
rect 38498 42926 38500 42978
rect 38444 42924 38500 42926
rect 39900 43932 39956 43988
rect 40124 43820 40180 43876
rect 40460 44044 40516 44100
rect 39676 43426 39732 43428
rect 39676 43374 39678 43426
rect 39678 43374 39730 43426
rect 39730 43374 39732 43426
rect 39676 43372 39732 43374
rect 39452 43036 39508 43092
rect 39564 43260 39620 43316
rect 37884 42530 37940 42532
rect 37884 42478 37886 42530
rect 37886 42478 37938 42530
rect 37938 42478 37940 42530
rect 37884 42476 37940 42478
rect 38220 41132 38276 41188
rect 38556 41804 38612 41860
rect 37660 40348 37716 40404
rect 37884 40460 37940 40516
rect 38332 40348 38388 40404
rect 37772 40236 37828 40292
rect 38108 40290 38164 40292
rect 38108 40238 38110 40290
rect 38110 40238 38162 40290
rect 38162 40238 38164 40290
rect 38108 40236 38164 40238
rect 38332 40124 38388 40180
rect 38780 40460 38836 40516
rect 38892 40908 38948 40964
rect 38892 40402 38948 40404
rect 38892 40350 38894 40402
rect 38894 40350 38946 40402
rect 38946 40350 38948 40402
rect 38892 40348 38948 40350
rect 40012 41916 40068 41972
rect 40012 40684 40068 40740
rect 40124 42924 40180 42980
rect 40124 42588 40180 42644
rect 36428 37938 36484 37940
rect 36428 37886 36430 37938
rect 36430 37886 36482 37938
rect 36482 37886 36484 37938
rect 36428 37884 36484 37886
rect 36092 37772 36148 37828
rect 34972 36988 35028 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 34860 36540 34916 36596
rect 35644 36428 35700 36484
rect 35308 35980 35364 36036
rect 35420 35868 35476 35924
rect 34860 35084 34916 35140
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34860 34242 34916 34244
rect 34860 34190 34862 34242
rect 34862 34190 34914 34242
rect 34914 34190 34916 34242
rect 34860 34188 34916 34190
rect 34636 34076 34692 34132
rect 35644 34914 35700 34916
rect 35644 34862 35646 34914
rect 35646 34862 35698 34914
rect 35698 34862 35700 34914
rect 35644 34860 35700 34862
rect 35532 34748 35588 34804
rect 35644 34300 35700 34356
rect 35980 35420 36036 35476
rect 37212 39452 37268 39508
rect 39004 40178 39060 40180
rect 39004 40126 39006 40178
rect 39006 40126 39058 40178
rect 39058 40126 39060 40178
rect 39004 40124 39060 40126
rect 38780 39506 38836 39508
rect 38780 39454 38782 39506
rect 38782 39454 38834 39506
rect 38834 39454 38836 39506
rect 38780 39452 38836 39454
rect 39116 39452 39172 39508
rect 38220 38780 38276 38836
rect 37212 37826 37268 37828
rect 37212 37774 37214 37826
rect 37214 37774 37266 37826
rect 37266 37774 37268 37826
rect 37212 37772 37268 37774
rect 36876 37436 36932 37492
rect 37884 37772 37940 37828
rect 36876 37100 36932 37156
rect 36204 36876 36260 36932
rect 36652 35756 36708 35812
rect 39340 39228 39396 39284
rect 40348 41858 40404 41860
rect 40348 41806 40350 41858
rect 40350 41806 40402 41858
rect 40402 41806 40404 41858
rect 40348 41804 40404 41806
rect 41468 44156 41524 44212
rect 41356 43932 41412 43988
rect 40572 40684 40628 40740
rect 40236 40348 40292 40404
rect 40348 40236 40404 40292
rect 38332 38050 38388 38052
rect 38332 37998 38334 38050
rect 38334 37998 38386 38050
rect 38386 37998 38388 38050
rect 38332 37996 38388 37998
rect 38444 37436 38500 37492
rect 37212 36428 37268 36484
rect 37100 35980 37156 36036
rect 36988 35922 37044 35924
rect 36988 35870 36990 35922
rect 36990 35870 37042 35922
rect 37042 35870 37044 35922
rect 36988 35868 37044 35870
rect 36428 35196 36484 35252
rect 36316 35026 36372 35028
rect 36316 34974 36318 35026
rect 36318 34974 36370 35026
rect 36370 34974 36372 35026
rect 36316 34972 36372 34974
rect 36988 34802 37044 34804
rect 36988 34750 36990 34802
rect 36990 34750 37042 34802
rect 37042 34750 37044 34802
rect 36988 34748 37044 34750
rect 35868 34130 35924 34132
rect 35868 34078 35870 34130
rect 35870 34078 35922 34130
rect 35922 34078 35924 34130
rect 35868 34076 35924 34078
rect 34748 33740 34804 33796
rect 34524 32508 34580 32564
rect 34300 32396 34356 32452
rect 33964 30828 34020 30884
rect 34412 31836 34468 31892
rect 33852 28812 33908 28868
rect 33740 28700 33796 28756
rect 33516 28028 33572 28084
rect 32508 27186 32564 27188
rect 32508 27134 32510 27186
rect 32510 27134 32562 27186
rect 32562 27134 32564 27186
rect 32508 27132 32564 27134
rect 33068 27692 33124 27748
rect 32396 26348 32452 26404
rect 32172 26012 32228 26068
rect 32508 25506 32564 25508
rect 32508 25454 32510 25506
rect 32510 25454 32562 25506
rect 32562 25454 32564 25506
rect 32508 25452 32564 25454
rect 32732 25506 32788 25508
rect 32732 25454 32734 25506
rect 32734 25454 32786 25506
rect 32786 25454 32788 25506
rect 32732 25452 32788 25454
rect 31948 25340 32004 25396
rect 32284 25282 32340 25284
rect 32284 25230 32286 25282
rect 32286 25230 32338 25282
rect 32338 25230 32340 25282
rect 32284 25228 32340 25230
rect 31724 24556 31780 24612
rect 32508 24610 32564 24612
rect 32508 24558 32510 24610
rect 32510 24558 32562 24610
rect 32562 24558 32564 24610
rect 32508 24556 32564 24558
rect 31836 24444 31892 24500
rect 31388 22204 31444 22260
rect 30940 21980 30996 22036
rect 30156 20748 30212 20804
rect 30044 20578 30100 20580
rect 30044 20526 30046 20578
rect 30046 20526 30098 20578
rect 30098 20526 30100 20578
rect 30044 20524 30100 20526
rect 30604 21308 30660 21364
rect 30716 20690 30772 20692
rect 30716 20638 30718 20690
rect 30718 20638 30770 20690
rect 30770 20638 30772 20690
rect 30716 20636 30772 20638
rect 30268 20524 30324 20580
rect 30828 20578 30884 20580
rect 30828 20526 30830 20578
rect 30830 20526 30882 20578
rect 30882 20526 30884 20578
rect 30828 20524 30884 20526
rect 31388 21532 31444 21588
rect 31724 23212 31780 23268
rect 31724 23042 31780 23044
rect 31724 22990 31726 23042
rect 31726 22990 31778 23042
rect 31778 22990 31780 23042
rect 31724 22988 31780 22990
rect 32396 23154 32452 23156
rect 32396 23102 32398 23154
rect 32398 23102 32450 23154
rect 32450 23102 32452 23154
rect 32396 23100 32452 23102
rect 31836 22428 31892 22484
rect 31612 21868 31668 21924
rect 31948 21980 32004 22036
rect 31500 21756 31556 21812
rect 31724 20242 31780 20244
rect 31724 20190 31726 20242
rect 31726 20190 31778 20242
rect 31778 20190 31780 20242
rect 31724 20188 31780 20190
rect 31836 19964 31892 20020
rect 30380 19852 30436 19908
rect 29260 19010 29316 19012
rect 29260 18958 29262 19010
rect 29262 18958 29314 19010
rect 29314 18958 29316 19010
rect 29260 18956 29316 18958
rect 30044 18562 30100 18564
rect 30044 18510 30046 18562
rect 30046 18510 30098 18562
rect 30098 18510 30100 18562
rect 30044 18508 30100 18510
rect 29148 18396 29204 18452
rect 30156 18450 30212 18452
rect 30156 18398 30158 18450
rect 30158 18398 30210 18450
rect 30210 18398 30212 18450
rect 30156 18396 30212 18398
rect 29932 18338 29988 18340
rect 29932 18286 29934 18338
rect 29934 18286 29986 18338
rect 29986 18286 29988 18338
rect 29932 18284 29988 18286
rect 29484 17500 29540 17556
rect 29484 16156 29540 16212
rect 30716 18508 30772 18564
rect 30716 18338 30772 18340
rect 30716 18286 30718 18338
rect 30718 18286 30770 18338
rect 30770 18286 30772 18338
rect 30716 18284 30772 18286
rect 30828 18396 30884 18452
rect 31500 18450 31556 18452
rect 31500 18398 31502 18450
rect 31502 18398 31554 18450
rect 31554 18398 31556 18450
rect 31500 18396 31556 18398
rect 32060 21810 32116 21812
rect 32060 21758 32062 21810
rect 32062 21758 32114 21810
rect 32114 21758 32116 21810
rect 32060 21756 32116 21758
rect 32172 20860 32228 20916
rect 32396 20076 32452 20132
rect 32060 19292 32116 19348
rect 31388 17948 31444 18004
rect 31500 17612 31556 17668
rect 30268 16716 30324 16772
rect 31388 17052 31444 17108
rect 30492 16380 30548 16436
rect 30044 15986 30100 15988
rect 30044 15934 30046 15986
rect 30046 15934 30098 15986
rect 30098 15934 30100 15986
rect 30044 15932 30100 15934
rect 28588 14924 28644 14980
rect 28476 14530 28532 14532
rect 28476 14478 28478 14530
rect 28478 14478 28530 14530
rect 28530 14478 28532 14530
rect 28476 14476 28532 14478
rect 28700 14028 28756 14084
rect 28476 13132 28532 13188
rect 28588 12850 28644 12852
rect 28588 12798 28590 12850
rect 28590 12798 28642 12850
rect 28642 12798 28644 12850
rect 28588 12796 28644 12798
rect 28476 12066 28532 12068
rect 28476 12014 28478 12066
rect 28478 12014 28530 12066
rect 28530 12014 28532 12066
rect 28476 12012 28532 12014
rect 28588 11564 28644 11620
rect 28924 12908 28980 12964
rect 28700 11900 28756 11956
rect 28812 12796 28868 12852
rect 28812 11788 28868 11844
rect 28364 11116 28420 11172
rect 28364 10668 28420 10724
rect 27692 10220 27748 10276
rect 27468 8428 27524 8484
rect 27580 8988 27636 9044
rect 28476 10220 28532 10276
rect 28140 9602 28196 9604
rect 28140 9550 28142 9602
rect 28142 9550 28194 9602
rect 28194 9550 28196 9602
rect 28140 9548 28196 9550
rect 27916 9266 27972 9268
rect 27916 9214 27918 9266
rect 27918 9214 27970 9266
rect 27970 9214 27972 9266
rect 27916 9212 27972 9214
rect 29260 14924 29316 14980
rect 29820 14924 29876 14980
rect 29372 14700 29428 14756
rect 29708 14700 29764 14756
rect 31276 15260 31332 15316
rect 30380 14642 30436 14644
rect 30380 14590 30382 14642
rect 30382 14590 30434 14642
rect 30434 14590 30436 14642
rect 30380 14588 30436 14590
rect 30828 14642 30884 14644
rect 30828 14590 30830 14642
rect 30830 14590 30882 14642
rect 30882 14590 30884 14642
rect 30828 14588 30884 14590
rect 29484 14364 29540 14420
rect 29260 14306 29316 14308
rect 29260 14254 29262 14306
rect 29262 14254 29314 14306
rect 29314 14254 29316 14306
rect 29260 14252 29316 14254
rect 29148 13020 29204 13076
rect 29372 12850 29428 12852
rect 29372 12798 29374 12850
rect 29374 12798 29426 12850
rect 29426 12798 29428 12850
rect 29372 12796 29428 12798
rect 29260 12348 29316 12404
rect 29148 12290 29204 12292
rect 29148 12238 29150 12290
rect 29150 12238 29202 12290
rect 29202 12238 29204 12290
rect 29148 12236 29204 12238
rect 29260 12066 29316 12068
rect 29260 12014 29262 12066
rect 29262 12014 29314 12066
rect 29314 12014 29316 12066
rect 29260 12012 29316 12014
rect 29372 11788 29428 11844
rect 29036 11004 29092 11060
rect 29820 13468 29876 13524
rect 29708 13132 29764 13188
rect 29596 12460 29652 12516
rect 30380 14418 30436 14420
rect 30380 14366 30382 14418
rect 30382 14366 30434 14418
rect 30434 14366 30436 14418
rect 30380 14364 30436 14366
rect 30268 14028 30324 14084
rect 30268 13858 30324 13860
rect 30268 13806 30270 13858
rect 30270 13806 30322 13858
rect 30322 13806 30324 13858
rect 30268 13804 30324 13806
rect 30940 14364 30996 14420
rect 30492 12460 30548 12516
rect 30268 12402 30324 12404
rect 30268 12350 30270 12402
rect 30270 12350 30322 12402
rect 30322 12350 30324 12402
rect 30268 12348 30324 12350
rect 30156 12236 30212 12292
rect 30828 12124 30884 12180
rect 30604 11564 30660 11620
rect 29372 10556 29428 10612
rect 29260 9996 29316 10052
rect 28476 8930 28532 8932
rect 28476 8878 28478 8930
rect 28478 8878 28530 8930
rect 28530 8878 28532 8930
rect 28476 8876 28532 8878
rect 27692 8204 27748 8260
rect 27804 8316 27860 8372
rect 26012 7420 26068 7476
rect 25564 6748 25620 6804
rect 25228 5906 25284 5908
rect 25228 5854 25230 5906
rect 25230 5854 25282 5906
rect 25282 5854 25284 5906
rect 25228 5852 25284 5854
rect 25116 5122 25172 5124
rect 25116 5070 25118 5122
rect 25118 5070 25170 5122
rect 25170 5070 25172 5122
rect 25116 5068 25172 5070
rect 26796 7362 26852 7364
rect 26796 7310 26798 7362
rect 26798 7310 26850 7362
rect 26850 7310 26852 7362
rect 26796 7308 26852 7310
rect 26908 6748 26964 6804
rect 26348 6524 26404 6580
rect 26236 6130 26292 6132
rect 26236 6078 26238 6130
rect 26238 6078 26290 6130
rect 26290 6078 26292 6130
rect 26236 6076 26292 6078
rect 26012 5852 26068 5908
rect 25676 5516 25732 5572
rect 26572 5906 26628 5908
rect 26572 5854 26574 5906
rect 26574 5854 26626 5906
rect 26626 5854 26628 5906
rect 26572 5852 26628 5854
rect 26684 5516 26740 5572
rect 28364 8204 28420 8260
rect 28252 6748 28308 6804
rect 28476 8146 28532 8148
rect 28476 8094 28478 8146
rect 28478 8094 28530 8146
rect 28530 8094 28532 8146
rect 28476 8092 28532 8094
rect 28364 7308 28420 7364
rect 28140 6690 28196 6692
rect 28140 6638 28142 6690
rect 28142 6638 28194 6690
rect 28194 6638 28196 6690
rect 28140 6636 28196 6638
rect 28588 6578 28644 6580
rect 28588 6526 28590 6578
rect 28590 6526 28642 6578
rect 28642 6526 28644 6578
rect 28588 6524 28644 6526
rect 23996 4620 24052 4676
rect 25228 4620 25284 4676
rect 24444 4450 24500 4452
rect 24444 4398 24446 4450
rect 24446 4398 24498 4450
rect 24498 4398 24500 4450
rect 24444 4396 24500 4398
rect 26460 5234 26516 5236
rect 26460 5182 26462 5234
rect 26462 5182 26514 5234
rect 26514 5182 26516 5234
rect 26460 5180 26516 5182
rect 26236 5068 26292 5124
rect 27244 5068 27300 5124
rect 23996 3554 24052 3556
rect 23996 3502 23998 3554
rect 23998 3502 24050 3554
rect 24050 3502 24052 3554
rect 23996 3500 24052 3502
rect 26012 3388 26068 3444
rect 23100 3276 23156 3332
rect 25340 3330 25396 3332
rect 25340 3278 25342 3330
rect 25342 3278 25394 3330
rect 25394 3278 25396 3330
rect 25340 3276 25396 3278
rect 26908 4898 26964 4900
rect 26908 4846 26910 4898
rect 26910 4846 26962 4898
rect 26962 4846 26964 4898
rect 26908 4844 26964 4846
rect 27580 5852 27636 5908
rect 27468 5404 27524 5460
rect 27580 5292 27636 5348
rect 27804 5122 27860 5124
rect 27804 5070 27806 5122
rect 27806 5070 27858 5122
rect 27858 5070 27860 5122
rect 27804 5068 27860 5070
rect 27356 4620 27412 4676
rect 28588 4620 28644 4676
rect 30604 10444 30660 10500
rect 30156 9154 30212 9156
rect 30156 9102 30158 9154
rect 30158 9102 30210 9154
rect 30210 9102 30212 9154
rect 30156 9100 30212 9102
rect 31052 11900 31108 11956
rect 33292 27298 33348 27300
rect 33292 27246 33294 27298
rect 33294 27246 33346 27298
rect 33346 27246 33348 27298
rect 33292 27244 33348 27246
rect 32956 26348 33012 26404
rect 33852 27244 33908 27300
rect 34076 28700 34132 28756
rect 34860 31276 34916 31332
rect 34748 30828 34804 30884
rect 34076 27244 34132 27300
rect 34188 28252 34244 28308
rect 33180 25788 33236 25844
rect 32956 25228 33012 25284
rect 33628 25282 33684 25284
rect 33628 25230 33630 25282
rect 33630 25230 33682 25282
rect 33682 25230 33684 25282
rect 33628 25228 33684 25230
rect 32396 18396 32452 18452
rect 32956 23772 33012 23828
rect 32844 19346 32900 19348
rect 32844 19294 32846 19346
rect 32846 19294 32898 19346
rect 32898 19294 32900 19346
rect 32844 19292 32900 19294
rect 34860 29820 34916 29876
rect 35868 33852 35924 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 33516 35252 33572
rect 35084 33404 35140 33460
rect 35084 33068 35140 33124
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 36540 34242 36596 34244
rect 36540 34190 36542 34242
rect 36542 34190 36594 34242
rect 36594 34190 36596 34242
rect 36540 34188 36596 34190
rect 36204 33234 36260 33236
rect 36204 33182 36206 33234
rect 36206 33182 36258 33234
rect 36258 33182 36260 33234
rect 36204 33180 36260 33182
rect 37548 35138 37604 35140
rect 37548 35086 37550 35138
rect 37550 35086 37602 35138
rect 37602 35086 37604 35138
rect 37548 35084 37604 35086
rect 37212 34914 37268 34916
rect 37212 34862 37214 34914
rect 37214 34862 37266 34914
rect 37266 34862 37268 34914
rect 37212 34860 37268 34862
rect 37212 34300 37268 34356
rect 37324 34188 37380 34244
rect 37772 35196 37828 35252
rect 37660 34076 37716 34132
rect 37772 34972 37828 35028
rect 35980 32508 36036 32564
rect 35868 32172 35924 32228
rect 36092 32396 36148 32452
rect 35756 31836 35812 31892
rect 35532 31778 35588 31780
rect 35532 31726 35534 31778
rect 35534 31726 35586 31778
rect 35586 31726 35588 31778
rect 35532 31724 35588 31726
rect 35868 31164 35924 31220
rect 35084 30716 35140 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 29484 35028 29540
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35756 29596 35812 29652
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34860 27132 34916 27188
rect 35308 27020 35364 27076
rect 33740 23772 33796 23828
rect 33964 23884 34020 23940
rect 34188 25676 34244 25732
rect 34188 24610 34244 24612
rect 34188 24558 34190 24610
rect 34190 24558 34242 24610
rect 34242 24558 34244 24610
rect 34188 24556 34244 24558
rect 34636 23938 34692 23940
rect 34636 23886 34638 23938
rect 34638 23886 34690 23938
rect 34690 23886 34692 23938
rect 34636 23884 34692 23886
rect 34076 23436 34132 23492
rect 33628 23324 33684 23380
rect 34188 23324 34244 23380
rect 33740 23266 33796 23268
rect 33740 23214 33742 23266
rect 33742 23214 33794 23266
rect 33794 23214 33796 23266
rect 33740 23212 33796 23214
rect 34636 23154 34692 23156
rect 34636 23102 34638 23154
rect 34638 23102 34690 23154
rect 34690 23102 34692 23154
rect 34636 23100 34692 23102
rect 33852 22258 33908 22260
rect 33852 22206 33854 22258
rect 33854 22206 33906 22258
rect 33906 22206 33908 22258
rect 33852 22204 33908 22206
rect 34524 22204 34580 22260
rect 33068 20860 33124 20916
rect 33628 20860 33684 20916
rect 33068 20076 33124 20132
rect 33516 20018 33572 20020
rect 33516 19966 33518 20018
rect 33518 19966 33570 20018
rect 33570 19966 33572 20018
rect 33516 19964 33572 19966
rect 34188 20914 34244 20916
rect 34188 20862 34190 20914
rect 34190 20862 34242 20914
rect 34242 20862 34244 20914
rect 34188 20860 34244 20862
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 25282 35252 25284
rect 35196 25230 35198 25282
rect 35198 25230 35250 25282
rect 35250 25230 35252 25282
rect 35196 25228 35252 25230
rect 34972 24668 35028 24724
rect 36204 31276 36260 31332
rect 35980 30882 36036 30884
rect 35980 30830 35982 30882
rect 35982 30830 36034 30882
rect 36034 30830 36036 30882
rect 35980 30828 36036 30830
rect 35980 30156 36036 30212
rect 36092 30098 36148 30100
rect 36092 30046 36094 30098
rect 36094 30046 36146 30098
rect 36146 30046 36148 30098
rect 36092 30044 36148 30046
rect 36092 29538 36148 29540
rect 36092 29486 36094 29538
rect 36094 29486 36146 29538
rect 36146 29486 36148 29538
rect 36092 29484 36148 29486
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 36988 31948 37044 32004
rect 37100 31890 37156 31892
rect 37100 31838 37102 31890
rect 37102 31838 37154 31890
rect 37154 31838 37156 31890
rect 37100 31836 37156 31838
rect 38892 37884 38948 37940
rect 38892 37490 38948 37492
rect 38892 37438 38894 37490
rect 38894 37438 38946 37490
rect 38946 37438 38948 37490
rect 38892 37436 38948 37438
rect 39340 38834 39396 38836
rect 39340 38782 39342 38834
rect 39342 38782 39394 38834
rect 39394 38782 39396 38834
rect 39340 38780 39396 38782
rect 40236 38780 40292 38836
rect 39116 37436 39172 37492
rect 39340 37548 39396 37604
rect 39564 37772 39620 37828
rect 40684 40460 40740 40516
rect 39676 37436 39732 37492
rect 39228 37100 39284 37156
rect 39452 36482 39508 36484
rect 39452 36430 39454 36482
rect 39454 36430 39506 36482
rect 39506 36430 39508 36482
rect 39452 36428 39508 36430
rect 39564 36988 39620 37044
rect 38780 36204 38836 36260
rect 38668 35756 38724 35812
rect 38444 35084 38500 35140
rect 38220 34188 38276 34244
rect 39004 35756 39060 35812
rect 39788 38220 39844 38276
rect 40236 37548 40292 37604
rect 39676 36876 39732 36932
rect 39676 35420 39732 35476
rect 41020 43372 41076 43428
rect 41244 43538 41300 43540
rect 41244 43486 41246 43538
rect 41246 43486 41298 43538
rect 41298 43486 41300 43538
rect 41244 43484 41300 43486
rect 41132 42700 41188 42756
rect 42924 45052 42980 45108
rect 42364 44044 42420 44100
rect 41692 43596 41748 43652
rect 42252 43820 42308 43876
rect 42140 43538 42196 43540
rect 42140 43486 42142 43538
rect 42142 43486 42194 43538
rect 42194 43486 42196 43538
rect 42140 43484 42196 43486
rect 41692 43314 41748 43316
rect 41692 43262 41694 43314
rect 41694 43262 41746 43314
rect 41746 43262 41748 43314
rect 41692 43260 41748 43262
rect 42476 43314 42532 43316
rect 42476 43262 42478 43314
rect 42478 43262 42530 43314
rect 42530 43262 42532 43314
rect 42476 43260 42532 43262
rect 41468 41244 41524 41300
rect 41692 42476 41748 42532
rect 41356 40572 41412 40628
rect 41020 40402 41076 40404
rect 41020 40350 41022 40402
rect 41022 40350 41074 40402
rect 41074 40350 41076 40402
rect 41020 40348 41076 40350
rect 41244 39506 41300 39508
rect 41244 39454 41246 39506
rect 41246 39454 41298 39506
rect 41298 39454 41300 39506
rect 41244 39452 41300 39454
rect 40796 38332 40852 38388
rect 40908 38220 40964 38276
rect 41356 37996 41412 38052
rect 41916 41916 41972 41972
rect 41020 37324 41076 37380
rect 40908 35980 40964 36036
rect 40236 34860 40292 34916
rect 39116 34300 39172 34356
rect 39340 34242 39396 34244
rect 39340 34190 39342 34242
rect 39342 34190 39394 34242
rect 39394 34190 39396 34242
rect 39340 34188 39396 34190
rect 41020 35308 41076 35364
rect 41244 35084 41300 35140
rect 41132 34914 41188 34916
rect 41132 34862 41134 34914
rect 41134 34862 41186 34914
rect 41186 34862 41188 34914
rect 41132 34860 41188 34862
rect 41468 37436 41524 37492
rect 41916 40124 41972 40180
rect 41916 39228 41972 39284
rect 42140 38892 42196 38948
rect 43036 44434 43092 44436
rect 43036 44382 43038 44434
rect 43038 44382 43090 44434
rect 43090 44382 43092 44434
rect 43036 44380 43092 44382
rect 45164 44380 45220 44436
rect 44156 44268 44212 44324
rect 43596 44210 43652 44212
rect 43596 44158 43598 44210
rect 43598 44158 43650 44210
rect 43650 44158 43652 44210
rect 43596 44156 43652 44158
rect 43708 43820 43764 43876
rect 43148 43708 43204 43764
rect 42924 42924 42980 42980
rect 42812 42866 42868 42868
rect 42812 42814 42814 42866
rect 42814 42814 42866 42866
rect 42866 42814 42868 42866
rect 42812 42812 42868 42814
rect 43148 43484 43204 43540
rect 43148 42364 43204 42420
rect 43484 42812 43540 42868
rect 43484 42252 43540 42308
rect 43932 43484 43988 43540
rect 44380 44098 44436 44100
rect 44380 44046 44382 44098
rect 44382 44046 44434 44098
rect 44434 44046 44436 44098
rect 44380 44044 44436 44046
rect 44268 43484 44324 43540
rect 44940 43708 44996 43764
rect 44492 43372 44548 43428
rect 43820 42476 43876 42532
rect 43820 42252 43876 42308
rect 43596 42028 43652 42084
rect 43708 42140 43764 42196
rect 43484 41804 43540 41860
rect 42588 40684 42644 40740
rect 42700 40348 42756 40404
rect 41356 34636 41412 34692
rect 41580 36092 41636 36148
rect 40460 34076 40516 34132
rect 38668 33740 38724 33796
rect 39788 33740 39844 33796
rect 40908 34130 40964 34132
rect 40908 34078 40910 34130
rect 40910 34078 40962 34130
rect 40962 34078 40964 34130
rect 40908 34076 40964 34078
rect 39788 33180 39844 33236
rect 38108 32620 38164 32676
rect 37996 32450 38052 32452
rect 37996 32398 37998 32450
rect 37998 32398 38050 32450
rect 38050 32398 38052 32450
rect 37996 32396 38052 32398
rect 37884 32284 37940 32340
rect 37324 31778 37380 31780
rect 37324 31726 37326 31778
rect 37326 31726 37378 31778
rect 37378 31726 37380 31778
rect 37324 31724 37380 31726
rect 37660 32060 37716 32116
rect 37548 31666 37604 31668
rect 37548 31614 37550 31666
rect 37550 31614 37602 31666
rect 37602 31614 37604 31666
rect 37548 31612 37604 31614
rect 37212 31388 37268 31444
rect 38892 32732 38948 32788
rect 39452 32620 39508 32676
rect 39004 32562 39060 32564
rect 39004 32510 39006 32562
rect 39006 32510 39058 32562
rect 39058 32510 39060 32562
rect 39004 32508 39060 32510
rect 39228 32450 39284 32452
rect 39228 32398 39230 32450
rect 39230 32398 39282 32450
rect 39282 32398 39284 32450
rect 39228 32396 39284 32398
rect 39340 31836 39396 31892
rect 40012 31666 40068 31668
rect 40012 31614 40014 31666
rect 40014 31614 40066 31666
rect 40066 31614 40068 31666
rect 40012 31612 40068 31614
rect 38332 31388 38388 31444
rect 37660 31276 37716 31332
rect 41468 32450 41524 32452
rect 41468 32398 41470 32450
rect 41470 32398 41522 32450
rect 41522 32398 41524 32450
rect 41468 32396 41524 32398
rect 41020 32060 41076 32116
rect 43932 41580 43988 41636
rect 43932 41356 43988 41412
rect 44268 42642 44324 42644
rect 44268 42590 44270 42642
rect 44270 42590 44322 42642
rect 44322 42590 44324 42642
rect 44268 42588 44324 42590
rect 44828 42642 44884 42644
rect 44828 42590 44830 42642
rect 44830 42590 44882 42642
rect 44882 42590 44884 42642
rect 44828 42588 44884 42590
rect 44156 42530 44212 42532
rect 44156 42478 44158 42530
rect 44158 42478 44210 42530
rect 44210 42478 44212 42530
rect 44156 42476 44212 42478
rect 43484 40684 43540 40740
rect 43148 39788 43204 39844
rect 43484 40460 43540 40516
rect 44156 40124 44212 40180
rect 43820 39676 43876 39732
rect 44268 39618 44324 39620
rect 44268 39566 44270 39618
rect 44270 39566 44322 39618
rect 44322 39566 44324 39618
rect 44268 39564 44324 39566
rect 43372 38444 43428 38500
rect 43484 38050 43540 38052
rect 43484 37998 43486 38050
rect 43486 37998 43538 38050
rect 43538 37998 43540 38050
rect 43484 37996 43540 37998
rect 43036 37772 43092 37828
rect 41916 36370 41972 36372
rect 41916 36318 41918 36370
rect 41918 36318 41970 36370
rect 41970 36318 41972 36370
rect 41916 36316 41972 36318
rect 41804 35868 41860 35924
rect 42028 35474 42084 35476
rect 42028 35422 42030 35474
rect 42030 35422 42082 35474
rect 42082 35422 42084 35474
rect 42028 35420 42084 35422
rect 42252 35868 42308 35924
rect 42476 36988 42532 37044
rect 42364 35308 42420 35364
rect 41692 34242 41748 34244
rect 41692 34190 41694 34242
rect 41694 34190 41746 34242
rect 41746 34190 41748 34242
rect 41692 34188 41748 34190
rect 41804 33292 41860 33348
rect 41916 32844 41972 32900
rect 41804 32732 41860 32788
rect 42140 34748 42196 34804
rect 42252 33292 42308 33348
rect 42028 32620 42084 32676
rect 40460 31836 40516 31892
rect 40236 31164 40292 31220
rect 36428 29986 36484 29988
rect 36428 29934 36430 29986
rect 36430 29934 36482 29986
rect 36482 29934 36484 29986
rect 36428 29932 36484 29934
rect 36092 27916 36148 27972
rect 36988 27916 37044 27972
rect 35980 27804 36036 27860
rect 36428 27132 36484 27188
rect 35980 26460 36036 26516
rect 36316 26178 36372 26180
rect 36316 26126 36318 26178
rect 36318 26126 36370 26178
rect 36370 26126 36372 26178
rect 36316 26124 36372 26126
rect 36316 25730 36372 25732
rect 36316 25678 36318 25730
rect 36318 25678 36370 25730
rect 36370 25678 36372 25730
rect 36316 25676 36372 25678
rect 36092 25340 36148 25396
rect 35868 24780 35924 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35868 24498 35924 24500
rect 35868 24446 35870 24498
rect 35870 24446 35922 24498
rect 35922 24446 35924 24498
rect 35868 24444 35924 24446
rect 35868 24220 35924 24276
rect 36204 24220 36260 24276
rect 36316 24780 36372 24836
rect 35196 23772 35252 23828
rect 34972 23212 35028 23268
rect 35868 23212 35924 23268
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35756 23154 35812 23156
rect 35756 23102 35758 23154
rect 35758 23102 35810 23154
rect 35810 23102 35812 23154
rect 35756 23100 35812 23102
rect 36204 23938 36260 23940
rect 36204 23886 36206 23938
rect 36206 23886 36258 23938
rect 36258 23886 36260 23938
rect 36204 23884 36260 23886
rect 39564 30940 39620 30996
rect 38332 30716 38388 30772
rect 37548 30210 37604 30212
rect 37548 30158 37550 30210
rect 37550 30158 37602 30210
rect 37602 30158 37604 30210
rect 37548 30156 37604 30158
rect 37212 29820 37268 29876
rect 38444 28812 38500 28868
rect 38444 28588 38500 28644
rect 37436 28364 37492 28420
rect 37324 27858 37380 27860
rect 37324 27806 37326 27858
rect 37326 27806 37378 27858
rect 37378 27806 37380 27858
rect 37324 27804 37380 27806
rect 37324 27132 37380 27188
rect 37548 27804 37604 27860
rect 37996 27244 38052 27300
rect 37884 27186 37940 27188
rect 37884 27134 37886 27186
rect 37886 27134 37938 27186
rect 37938 27134 37940 27186
rect 37884 27132 37940 27134
rect 37884 26460 37940 26516
rect 36764 26178 36820 26180
rect 36764 26126 36766 26178
rect 36766 26126 36818 26178
rect 36818 26126 36820 26178
rect 36764 26124 36820 26126
rect 39116 28642 39172 28644
rect 39116 28590 39118 28642
rect 39118 28590 39170 28642
rect 39170 28590 39172 28642
rect 39116 28588 39172 28590
rect 40124 30770 40180 30772
rect 40124 30718 40126 30770
rect 40126 30718 40178 30770
rect 40178 30718 40180 30770
rect 40124 30716 40180 30718
rect 39788 30156 39844 30212
rect 39676 29932 39732 29988
rect 39788 29708 39844 29764
rect 40348 30156 40404 30212
rect 39788 28924 39844 28980
rect 39900 28812 39956 28868
rect 39900 28642 39956 28644
rect 39900 28590 39902 28642
rect 39902 28590 39954 28642
rect 39954 28590 39956 28642
rect 39900 28588 39956 28590
rect 39564 28364 39620 28420
rect 40124 28364 40180 28420
rect 38892 27970 38948 27972
rect 38892 27918 38894 27970
rect 38894 27918 38946 27970
rect 38946 27918 38948 27970
rect 38892 27916 38948 27918
rect 38780 27858 38836 27860
rect 38780 27806 38782 27858
rect 38782 27806 38834 27858
rect 38834 27806 38836 27858
rect 38780 27804 38836 27806
rect 38780 27244 38836 27300
rect 39228 27804 39284 27860
rect 37660 26178 37716 26180
rect 37660 26126 37662 26178
rect 37662 26126 37714 26178
rect 37714 26126 37716 26178
rect 37660 26124 37716 26126
rect 37324 25452 37380 25508
rect 37548 25452 37604 25508
rect 36652 25228 36708 25284
rect 37436 25340 37492 25396
rect 37100 25116 37156 25172
rect 36764 24834 36820 24836
rect 36764 24782 36766 24834
rect 36766 24782 36818 24834
rect 36818 24782 36820 24834
rect 36764 24780 36820 24782
rect 36204 23212 36260 23268
rect 36540 24220 36596 24276
rect 35644 22204 35700 22260
rect 35308 22092 35364 22148
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35308 21026 35364 21028
rect 35308 20974 35310 21026
rect 35310 20974 35362 21026
rect 35362 20974 35364 21026
rect 35308 20972 35364 20974
rect 33740 20188 33796 20244
rect 33292 19852 33348 19908
rect 34188 20130 34244 20132
rect 34188 20078 34190 20130
rect 34190 20078 34242 20130
rect 34242 20078 34244 20130
rect 34188 20076 34244 20078
rect 33740 19740 33796 19796
rect 33404 18620 33460 18676
rect 31724 17890 31780 17892
rect 31724 17838 31726 17890
rect 31726 17838 31778 17890
rect 31778 17838 31780 17890
rect 31724 17836 31780 17838
rect 31948 17948 32004 18004
rect 31836 17500 31892 17556
rect 31724 16994 31780 16996
rect 31724 16942 31726 16994
rect 31726 16942 31778 16994
rect 31778 16942 31780 16994
rect 31724 16940 31780 16942
rect 31724 16492 31780 16548
rect 31276 14476 31332 14532
rect 31948 16716 32004 16772
rect 32396 17666 32452 17668
rect 32396 17614 32398 17666
rect 32398 17614 32450 17666
rect 32450 17614 32452 17666
rect 32396 17612 32452 17614
rect 32060 16380 32116 16436
rect 32284 16882 32340 16884
rect 32284 16830 32286 16882
rect 32286 16830 32338 16882
rect 32338 16830 32340 16882
rect 32284 16828 32340 16830
rect 32060 16210 32116 16212
rect 32060 16158 32062 16210
rect 32062 16158 32114 16210
rect 32114 16158 32116 16210
rect 32060 16156 32116 16158
rect 32172 15148 32228 15204
rect 31500 13692 31556 13748
rect 31948 14476 32004 14532
rect 31388 13580 31444 13636
rect 31388 10892 31444 10948
rect 31276 10610 31332 10612
rect 31276 10558 31278 10610
rect 31278 10558 31330 10610
rect 31330 10558 31332 10610
rect 31276 10556 31332 10558
rect 31276 9996 31332 10052
rect 31500 9996 31556 10052
rect 30940 9548 30996 9604
rect 31164 9884 31220 9940
rect 31164 9212 31220 9268
rect 30492 8988 30548 9044
rect 29036 8258 29092 8260
rect 29036 8206 29038 8258
rect 29038 8206 29090 8258
rect 29090 8206 29092 8258
rect 29036 8204 29092 8206
rect 29260 8146 29316 8148
rect 29260 8094 29262 8146
rect 29262 8094 29314 8146
rect 29314 8094 29316 8146
rect 29260 8092 29316 8094
rect 29820 8764 29876 8820
rect 29484 7756 29540 7812
rect 29596 8316 29652 8372
rect 29260 6636 29316 6692
rect 29148 5346 29204 5348
rect 29148 5294 29150 5346
rect 29150 5294 29202 5346
rect 29202 5294 29204 5346
rect 29148 5292 29204 5294
rect 26684 3612 26740 3668
rect 27580 3666 27636 3668
rect 27580 3614 27582 3666
rect 27582 3614 27634 3666
rect 27634 3614 27636 3666
rect 27580 3612 27636 3614
rect 28140 3612 28196 3668
rect 28812 4284 28868 4340
rect 29484 4844 29540 4900
rect 29260 4226 29316 4228
rect 29260 4174 29262 4226
rect 29262 4174 29314 4226
rect 29314 4174 29316 4226
rect 29260 4172 29316 4174
rect 29932 8316 29988 8372
rect 30156 7868 30212 7924
rect 30268 6748 30324 6804
rect 30044 6524 30100 6580
rect 30940 6636 30996 6692
rect 30380 5346 30436 5348
rect 30380 5294 30382 5346
rect 30382 5294 30434 5346
rect 30434 5294 30436 5346
rect 30380 5292 30436 5294
rect 31388 9100 31444 9156
rect 31836 12850 31892 12852
rect 31836 12798 31838 12850
rect 31838 12798 31890 12850
rect 31890 12798 31892 12850
rect 31836 12796 31892 12798
rect 31724 12460 31780 12516
rect 31948 10892 32004 10948
rect 32620 16828 32676 16884
rect 32396 16492 32452 16548
rect 32172 13970 32228 13972
rect 32172 13918 32174 13970
rect 32174 13918 32226 13970
rect 32226 13918 32228 13970
rect 32172 13916 32228 13918
rect 32732 14530 32788 14532
rect 32732 14478 32734 14530
rect 32734 14478 32786 14530
rect 32786 14478 32788 14530
rect 32732 14476 32788 14478
rect 32508 13634 32564 13636
rect 32508 13582 32510 13634
rect 32510 13582 32562 13634
rect 32562 13582 32564 13634
rect 32508 13580 32564 13582
rect 33292 18396 33348 18452
rect 33964 18508 34020 18564
rect 33740 18172 33796 18228
rect 33628 17836 33684 17892
rect 33068 17052 33124 17108
rect 33404 16492 33460 16548
rect 33516 16882 33572 16884
rect 33516 16830 33518 16882
rect 33518 16830 33570 16882
rect 33570 16830 33572 16882
rect 33516 16828 33572 16830
rect 33180 16380 33236 16436
rect 33180 16098 33236 16100
rect 33180 16046 33182 16098
rect 33182 16046 33234 16098
rect 33234 16046 33236 16098
rect 33180 16044 33236 16046
rect 33180 14700 33236 14756
rect 33292 14364 33348 14420
rect 32844 13132 32900 13188
rect 33180 14140 33236 14196
rect 32620 12962 32676 12964
rect 32620 12910 32622 12962
rect 32622 12910 32674 12962
rect 32674 12910 32676 12962
rect 32620 12908 32676 12910
rect 32396 12572 32452 12628
rect 32172 12066 32228 12068
rect 32172 12014 32174 12066
rect 32174 12014 32226 12066
rect 32226 12014 32228 12066
rect 32172 12012 32228 12014
rect 32508 12124 32564 12180
rect 32508 11116 32564 11172
rect 32620 11788 32676 11844
rect 32508 10780 32564 10836
rect 32172 10498 32228 10500
rect 32172 10446 32174 10498
rect 32174 10446 32226 10498
rect 32226 10446 32228 10498
rect 32172 10444 32228 10446
rect 31724 8876 31780 8932
rect 31612 8764 31668 8820
rect 31836 7644 31892 7700
rect 32508 9938 32564 9940
rect 32508 9886 32510 9938
rect 32510 9886 32562 9938
rect 32562 9886 32564 9938
rect 32508 9884 32564 9886
rect 32284 8818 32340 8820
rect 32284 8766 32286 8818
rect 32286 8766 32338 8818
rect 32338 8766 32340 8818
rect 32284 8764 32340 8766
rect 33292 13692 33348 13748
rect 33180 12738 33236 12740
rect 33180 12686 33182 12738
rect 33182 12686 33234 12738
rect 33234 12686 33236 12738
rect 33180 12684 33236 12686
rect 33180 12348 33236 12404
rect 33180 12124 33236 12180
rect 34524 20018 34580 20020
rect 34524 19966 34526 20018
rect 34526 19966 34578 20018
rect 34578 19966 34580 20018
rect 34524 19964 34580 19966
rect 34412 19906 34468 19908
rect 34412 19854 34414 19906
rect 34414 19854 34466 19906
rect 34466 19854 34468 19906
rect 34412 19852 34468 19854
rect 34524 19740 34580 19796
rect 34412 18396 34468 18452
rect 34188 17612 34244 17668
rect 34300 17554 34356 17556
rect 34300 17502 34302 17554
rect 34302 17502 34354 17554
rect 34354 17502 34356 17554
rect 34300 17500 34356 17502
rect 34748 19180 34804 19236
rect 34860 18396 34916 18452
rect 34972 20524 35028 20580
rect 34076 17052 34132 17108
rect 34748 17442 34804 17444
rect 34748 17390 34750 17442
rect 34750 17390 34802 17442
rect 34802 17390 34804 17442
rect 34748 17388 34804 17390
rect 34300 16492 34356 16548
rect 34188 16156 34244 16212
rect 33628 15202 33684 15204
rect 33628 15150 33630 15202
rect 33630 15150 33682 15202
rect 33682 15150 33684 15202
rect 33628 15148 33684 15150
rect 33740 14140 33796 14196
rect 33852 14418 33908 14420
rect 33852 14366 33854 14418
rect 33854 14366 33906 14418
rect 33906 14366 33908 14418
rect 33852 14364 33908 14366
rect 33628 12962 33684 12964
rect 33628 12910 33630 12962
rect 33630 12910 33682 12962
rect 33682 12910 33684 12962
rect 33628 12908 33684 12910
rect 33404 12572 33460 12628
rect 33068 10892 33124 10948
rect 33068 10610 33124 10612
rect 33068 10558 33070 10610
rect 33070 10558 33122 10610
rect 33122 10558 33124 10610
rect 33068 10556 33124 10558
rect 32956 9938 33012 9940
rect 32956 9886 32958 9938
rect 32958 9886 33010 9938
rect 33010 9886 33012 9938
rect 32956 9884 33012 9886
rect 33292 9996 33348 10052
rect 32620 8316 32676 8372
rect 33068 8876 33124 8932
rect 33180 8204 33236 8260
rect 34636 16882 34692 16884
rect 34636 16830 34638 16882
rect 34638 16830 34690 16882
rect 34690 16830 34692 16882
rect 34636 16828 34692 16830
rect 34524 15036 34580 15092
rect 35644 19906 35700 19908
rect 35644 19854 35646 19906
rect 35646 19854 35698 19906
rect 35698 19854 35700 19906
rect 35644 19852 35700 19854
rect 35196 19794 35252 19796
rect 35196 19742 35198 19794
rect 35198 19742 35250 19794
rect 35250 19742 35252 19794
rect 35196 19740 35252 19742
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 18620 35140 18676
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35644 19628 35700 19684
rect 35756 18620 35812 18676
rect 35196 17442 35252 17444
rect 35196 17390 35198 17442
rect 35198 17390 35250 17442
rect 35250 17390 35252 17442
rect 35196 17388 35252 17390
rect 34748 15148 34804 15204
rect 34972 16940 35028 16996
rect 35644 17388 35700 17444
rect 35532 16716 35588 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35084 15932 35140 15988
rect 33964 12348 34020 12404
rect 33740 12178 33796 12180
rect 33740 12126 33742 12178
rect 33742 12126 33794 12178
rect 33794 12126 33796 12178
rect 33740 12124 33796 12126
rect 34300 12012 34356 12068
rect 33852 11116 33908 11172
rect 34412 11394 34468 11396
rect 34412 11342 34414 11394
rect 34414 11342 34466 11394
rect 34466 11342 34468 11394
rect 34412 11340 34468 11342
rect 34412 9884 34468 9940
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 13468 35028 13524
rect 35644 15372 35700 15428
rect 36092 20130 36148 20132
rect 36092 20078 36094 20130
rect 36094 20078 36146 20130
rect 36146 20078 36148 20130
rect 36092 20076 36148 20078
rect 36204 19404 36260 19460
rect 38108 24892 38164 24948
rect 38220 25564 38276 25620
rect 39564 26572 39620 26628
rect 38444 26514 38500 26516
rect 38444 26462 38446 26514
rect 38446 26462 38498 26514
rect 38498 26462 38500 26514
rect 38444 26460 38500 26462
rect 39788 27692 39844 27748
rect 40012 27074 40068 27076
rect 40012 27022 40014 27074
rect 40014 27022 40066 27074
rect 40066 27022 40068 27074
rect 40012 27020 40068 27022
rect 41580 31836 41636 31892
rect 41804 31724 41860 31780
rect 40348 28812 40404 28868
rect 40796 29596 40852 29652
rect 41020 28924 41076 28980
rect 41804 31218 41860 31220
rect 41804 31166 41806 31218
rect 41806 31166 41858 31218
rect 41858 31166 41860 31218
rect 41804 31164 41860 31166
rect 41580 30994 41636 30996
rect 41580 30942 41582 30994
rect 41582 30942 41634 30994
rect 41634 30942 41636 30994
rect 41580 30940 41636 30942
rect 40572 28418 40628 28420
rect 40572 28366 40574 28418
rect 40574 28366 40626 28418
rect 40626 28366 40628 28418
rect 40572 28364 40628 28366
rect 40796 27468 40852 27524
rect 40348 27132 40404 27188
rect 40572 26796 40628 26852
rect 40348 26684 40404 26740
rect 38556 25564 38612 25620
rect 38332 25282 38388 25284
rect 38332 25230 38334 25282
rect 38334 25230 38386 25282
rect 38386 25230 38388 25282
rect 38332 25228 38388 25230
rect 38780 25452 38836 25508
rect 38892 26124 38948 26180
rect 38108 24722 38164 24724
rect 38108 24670 38110 24722
rect 38110 24670 38162 24722
rect 38162 24670 38164 24722
rect 38108 24668 38164 24670
rect 37660 24108 37716 24164
rect 38332 24108 38388 24164
rect 36988 23826 37044 23828
rect 36988 23774 36990 23826
rect 36990 23774 37042 23826
rect 37042 23774 37044 23826
rect 36988 23772 37044 23774
rect 36540 21644 36596 21700
rect 36652 19964 36708 20020
rect 36092 17164 36148 17220
rect 35980 16940 36036 16996
rect 36092 16098 36148 16100
rect 36092 16046 36094 16098
rect 36094 16046 36146 16098
rect 36146 16046 36148 16098
rect 36092 16044 36148 16046
rect 35868 14700 35924 14756
rect 35868 14530 35924 14532
rect 35868 14478 35870 14530
rect 35870 14478 35922 14530
rect 35922 14478 35924 14530
rect 35868 14476 35924 14478
rect 35644 13580 35700 13636
rect 36204 14530 36260 14532
rect 36204 14478 36206 14530
rect 36206 14478 36258 14530
rect 36258 14478 36260 14530
rect 36204 14476 36260 14478
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 12348 35140 12404
rect 35196 12012 35252 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36092 13468 36148 13524
rect 35532 11228 35588 11284
rect 35532 11004 35588 11060
rect 34300 9324 34356 9380
rect 34748 9996 34804 10052
rect 33628 9266 33684 9268
rect 33628 9214 33630 9266
rect 33630 9214 33682 9266
rect 33682 9214 33684 9266
rect 33628 9212 33684 9214
rect 33292 7868 33348 7924
rect 33180 7698 33236 7700
rect 33180 7646 33182 7698
rect 33182 7646 33234 7698
rect 33234 7646 33236 7698
rect 33180 7644 33236 7646
rect 32508 7586 32564 7588
rect 32508 7534 32510 7586
rect 32510 7534 32562 7586
rect 32562 7534 32564 7586
rect 32508 7532 32564 7534
rect 32284 7474 32340 7476
rect 32284 7422 32286 7474
rect 32286 7422 32338 7474
rect 32338 7422 32340 7474
rect 32284 7420 32340 7422
rect 31948 6690 32004 6692
rect 31948 6638 31950 6690
rect 31950 6638 32002 6690
rect 32002 6638 32004 6690
rect 31948 6636 32004 6638
rect 31836 5852 31892 5908
rect 32172 6188 32228 6244
rect 31948 5740 32004 5796
rect 31276 5292 31332 5348
rect 31612 5516 31668 5572
rect 30940 5122 30996 5124
rect 30940 5070 30942 5122
rect 30942 5070 30994 5122
rect 30994 5070 30996 5122
rect 30940 5068 30996 5070
rect 29820 4508 29876 4564
rect 31388 3724 31444 3780
rect 30940 3612 30996 3668
rect 31724 5010 31780 5012
rect 31724 4958 31726 5010
rect 31726 4958 31778 5010
rect 31778 4958 31780 5010
rect 31724 4956 31780 4958
rect 31836 4562 31892 4564
rect 31836 4510 31838 4562
rect 31838 4510 31890 4562
rect 31890 4510 31892 4562
rect 31836 4508 31892 4510
rect 31612 4172 31668 4228
rect 33852 9042 33908 9044
rect 33852 8990 33854 9042
rect 33854 8990 33906 9042
rect 33906 8990 33908 9042
rect 33852 8988 33908 8990
rect 33404 8316 33460 8372
rect 34300 8428 34356 8484
rect 33516 8092 33572 8148
rect 33404 7196 33460 7252
rect 33516 7420 33572 7476
rect 34524 9212 34580 9268
rect 34076 8258 34132 8260
rect 34076 8206 34078 8258
rect 34078 8206 34130 8258
rect 34130 8206 34132 8258
rect 34076 8204 34132 8206
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35756 10780 35812 10836
rect 35868 12124 35924 12180
rect 35980 12012 36036 12068
rect 36204 11900 36260 11956
rect 35644 10108 35700 10164
rect 35756 10556 35812 10612
rect 35532 9436 35588 9492
rect 35980 11676 36036 11732
rect 35980 11282 36036 11284
rect 35980 11230 35982 11282
rect 35982 11230 36034 11282
rect 36034 11230 36036 11282
rect 35980 11228 36036 11230
rect 36652 18620 36708 18676
rect 36540 16828 36596 16884
rect 36652 17164 36708 17220
rect 37436 23212 37492 23268
rect 37884 23660 37940 23716
rect 37324 22258 37380 22260
rect 37324 22206 37326 22258
rect 37326 22206 37378 22258
rect 37378 22206 37380 22258
rect 37324 22204 37380 22206
rect 36988 22146 37044 22148
rect 36988 22094 36990 22146
rect 36990 22094 37042 22146
rect 37042 22094 37044 22146
rect 36988 22092 37044 22094
rect 37772 22988 37828 23044
rect 38108 23714 38164 23716
rect 38108 23662 38110 23714
rect 38110 23662 38162 23714
rect 38162 23662 38164 23714
rect 38108 23660 38164 23662
rect 38444 23660 38500 23716
rect 38332 23324 38388 23380
rect 38780 25228 38836 25284
rect 39004 25228 39060 25284
rect 38780 24556 38836 24612
rect 39004 24610 39060 24612
rect 39004 24558 39006 24610
rect 39006 24558 39058 24610
rect 39058 24558 39060 24610
rect 39004 24556 39060 24558
rect 39452 24722 39508 24724
rect 39452 24670 39454 24722
rect 39454 24670 39506 24722
rect 39506 24670 39508 24722
rect 39452 24668 39508 24670
rect 39676 25228 39732 25284
rect 38556 23154 38612 23156
rect 38556 23102 38558 23154
rect 38558 23102 38610 23154
rect 38610 23102 38612 23154
rect 38556 23100 38612 23102
rect 37996 22876 38052 22932
rect 39116 23266 39172 23268
rect 39116 23214 39118 23266
rect 39118 23214 39170 23266
rect 39170 23214 39172 23266
rect 39116 23212 39172 23214
rect 36988 20972 37044 21028
rect 38444 21980 38500 22036
rect 37884 21196 37940 21252
rect 37100 19906 37156 19908
rect 37100 19854 37102 19906
rect 37102 19854 37154 19906
rect 37154 19854 37156 19906
rect 37100 19852 37156 19854
rect 38892 22146 38948 22148
rect 38892 22094 38894 22146
rect 38894 22094 38946 22146
rect 38946 22094 38948 22146
rect 38892 22092 38948 22094
rect 39228 23154 39284 23156
rect 39228 23102 39230 23154
rect 39230 23102 39282 23154
rect 39282 23102 39284 23154
rect 39228 23100 39284 23102
rect 39900 25004 39956 25060
rect 40236 26178 40292 26180
rect 40236 26126 40238 26178
rect 40238 26126 40290 26178
rect 40290 26126 40292 26178
rect 40236 26124 40292 26126
rect 40236 25564 40292 25620
rect 40124 24780 40180 24836
rect 40796 25618 40852 25620
rect 40796 25566 40798 25618
rect 40798 25566 40850 25618
rect 40850 25566 40852 25618
rect 40796 25564 40852 25566
rect 41244 27804 41300 27860
rect 41020 27692 41076 27748
rect 41020 27074 41076 27076
rect 41020 27022 41022 27074
rect 41022 27022 41074 27074
rect 41074 27022 41076 27074
rect 41020 27020 41076 27022
rect 41244 27074 41300 27076
rect 41244 27022 41246 27074
rect 41246 27022 41298 27074
rect 41298 27022 41300 27074
rect 41244 27020 41300 27022
rect 43260 37436 43316 37492
rect 43372 37154 43428 37156
rect 43372 37102 43374 37154
rect 43374 37102 43426 37154
rect 43426 37102 43428 37154
rect 43372 37100 43428 37102
rect 43036 35868 43092 35924
rect 43484 36988 43540 37044
rect 44156 37938 44212 37940
rect 44156 37886 44158 37938
rect 44158 37886 44210 37938
rect 44210 37886 44212 37938
rect 44156 37884 44212 37886
rect 44380 37826 44436 37828
rect 44380 37774 44382 37826
rect 44382 37774 44434 37826
rect 44434 37774 44436 37826
rect 44380 37772 44436 37774
rect 44044 37548 44100 37604
rect 43932 37100 43988 37156
rect 43708 36764 43764 36820
rect 43148 35138 43204 35140
rect 43148 35086 43150 35138
rect 43150 35086 43202 35138
rect 43202 35086 43204 35138
rect 43148 35084 43204 35086
rect 44940 42364 44996 42420
rect 44604 42252 44660 42308
rect 44604 42028 44660 42084
rect 44716 41970 44772 41972
rect 44716 41918 44718 41970
rect 44718 41918 44770 41970
rect 44770 41918 44772 41970
rect 44716 41916 44772 41918
rect 44828 41186 44884 41188
rect 44828 41134 44830 41186
rect 44830 41134 44882 41186
rect 44882 41134 44884 41186
rect 44828 41132 44884 41134
rect 44716 41020 44772 41076
rect 44604 40572 44660 40628
rect 45612 44098 45668 44100
rect 45612 44046 45614 44098
rect 45614 44046 45666 44098
rect 45666 44046 45668 44098
rect 45612 44044 45668 44046
rect 45948 43596 46004 43652
rect 45276 42812 45332 42868
rect 45164 42140 45220 42196
rect 45500 42140 45556 42196
rect 45388 41580 45444 41636
rect 45164 41410 45220 41412
rect 45164 41358 45166 41410
rect 45166 41358 45218 41410
rect 45218 41358 45220 41410
rect 45164 41356 45220 41358
rect 44940 40684 44996 40740
rect 45164 40402 45220 40404
rect 45164 40350 45166 40402
rect 45166 40350 45218 40402
rect 45218 40350 45220 40402
rect 45164 40348 45220 40350
rect 45836 41298 45892 41300
rect 45836 41246 45838 41298
rect 45838 41246 45890 41298
rect 45890 41246 45892 41298
rect 45836 41244 45892 41246
rect 46060 42476 46116 42532
rect 45948 41132 46004 41188
rect 46284 42252 46340 42308
rect 45612 41020 45668 41076
rect 45052 39564 45108 39620
rect 45164 39394 45220 39396
rect 45164 39342 45166 39394
rect 45166 39342 45218 39394
rect 45218 39342 45220 39394
rect 45164 39340 45220 39342
rect 45164 38834 45220 38836
rect 45164 38782 45166 38834
rect 45166 38782 45218 38834
rect 45218 38782 45220 38834
rect 45164 38780 45220 38782
rect 44716 38444 44772 38500
rect 44940 38162 44996 38164
rect 44940 38110 44942 38162
rect 44942 38110 44994 38162
rect 44994 38110 44996 38162
rect 44940 38108 44996 38110
rect 45052 38050 45108 38052
rect 45052 37998 45054 38050
rect 45054 37998 45106 38050
rect 45106 37998 45108 38050
rect 45052 37996 45108 37998
rect 45612 40626 45668 40628
rect 45612 40574 45614 40626
rect 45614 40574 45666 40626
rect 45666 40574 45668 40626
rect 45612 40572 45668 40574
rect 45948 40962 46004 40964
rect 45948 40910 45950 40962
rect 45950 40910 46002 40962
rect 46002 40910 46004 40962
rect 45948 40908 46004 40910
rect 45836 40684 45892 40740
rect 45724 40348 45780 40404
rect 45948 39340 46004 39396
rect 45612 39004 45668 39060
rect 44940 36764 44996 36820
rect 44828 36370 44884 36372
rect 44828 36318 44830 36370
rect 44830 36318 44882 36370
rect 44882 36318 44884 36370
rect 44828 36316 44884 36318
rect 44940 36258 44996 36260
rect 44940 36206 44942 36258
rect 44942 36206 44994 36258
rect 44994 36206 44996 36258
rect 44940 36204 44996 36206
rect 43708 35084 43764 35140
rect 43820 34972 43876 35028
rect 43372 34636 43428 34692
rect 43708 34300 43764 34356
rect 43484 34188 43540 34244
rect 45948 38332 46004 38388
rect 46172 39394 46228 39396
rect 46172 39342 46174 39394
rect 46174 39342 46226 39394
rect 46226 39342 46228 39394
rect 46172 39340 46228 39342
rect 45276 36204 45332 36260
rect 44828 34802 44884 34804
rect 44828 34750 44830 34802
rect 44830 34750 44882 34802
rect 44882 34750 44884 34802
rect 44828 34748 44884 34750
rect 45052 34636 45108 34692
rect 44828 34354 44884 34356
rect 44828 34302 44830 34354
rect 44830 34302 44882 34354
rect 44882 34302 44884 34354
rect 44828 34300 44884 34302
rect 43932 33740 43988 33796
rect 42476 33516 42532 33572
rect 42812 33346 42868 33348
rect 42812 33294 42814 33346
rect 42814 33294 42866 33346
rect 42866 33294 42868 33346
rect 42812 33292 42868 33294
rect 42476 32844 42532 32900
rect 44156 32732 44212 32788
rect 42476 32284 42532 32340
rect 42812 32172 42868 32228
rect 42588 31500 42644 31556
rect 42364 31106 42420 31108
rect 42364 31054 42366 31106
rect 42366 31054 42418 31106
rect 42418 31054 42420 31106
rect 42364 31052 42420 31054
rect 42252 30156 42308 30212
rect 42588 30044 42644 30100
rect 41916 28924 41972 28980
rect 42476 28924 42532 28980
rect 41692 28700 41748 28756
rect 42364 28812 42420 28868
rect 42252 28588 42308 28644
rect 42140 27858 42196 27860
rect 42140 27806 42142 27858
rect 42142 27806 42194 27858
rect 42194 27806 42196 27858
rect 42140 27804 42196 27806
rect 41916 27580 41972 27636
rect 41804 27132 41860 27188
rect 41468 26684 41524 26740
rect 41580 26796 41636 26852
rect 41132 25564 41188 25620
rect 41468 26124 41524 26180
rect 40124 24556 40180 24612
rect 40684 25282 40740 25284
rect 40684 25230 40686 25282
rect 40686 25230 40738 25282
rect 40738 25230 40740 25282
rect 40684 25228 40740 25230
rect 40460 24668 40516 24724
rect 40124 23938 40180 23940
rect 40124 23886 40126 23938
rect 40126 23886 40178 23938
rect 40178 23886 40180 23938
rect 40124 23884 40180 23886
rect 40460 23772 40516 23828
rect 39228 22482 39284 22484
rect 39228 22430 39230 22482
rect 39230 22430 39282 22482
rect 39282 22430 39284 22482
rect 39228 22428 39284 22430
rect 38108 21698 38164 21700
rect 38108 21646 38110 21698
rect 38110 21646 38162 21698
rect 38162 21646 38164 21698
rect 38108 21644 38164 21646
rect 38108 20748 38164 20804
rect 37996 20690 38052 20692
rect 37996 20638 37998 20690
rect 37998 20638 38050 20690
rect 38050 20638 38052 20690
rect 37996 20636 38052 20638
rect 38556 21084 38612 21140
rect 39676 21810 39732 21812
rect 39676 21758 39678 21810
rect 39678 21758 39730 21810
rect 39730 21758 39732 21810
rect 39676 21756 39732 21758
rect 39676 21532 39732 21588
rect 39340 21196 39396 21252
rect 39564 21420 39620 21476
rect 41692 26572 41748 26628
rect 42140 26572 42196 26628
rect 41804 26460 41860 26516
rect 42028 25506 42084 25508
rect 42028 25454 42030 25506
rect 42030 25454 42082 25506
rect 42082 25454 42084 25506
rect 42028 25452 42084 25454
rect 41468 25228 41524 25284
rect 40908 25116 40964 25172
rect 41468 25004 41524 25060
rect 41132 24892 41188 24948
rect 41020 24834 41076 24836
rect 41020 24782 41022 24834
rect 41022 24782 41074 24834
rect 41074 24782 41076 24834
rect 41020 24780 41076 24782
rect 40908 24556 40964 24612
rect 41580 24722 41636 24724
rect 41580 24670 41582 24722
rect 41582 24670 41634 24722
rect 41634 24670 41636 24722
rect 41580 24668 41636 24670
rect 41692 24444 41748 24500
rect 43484 32284 43540 32340
rect 42812 29596 42868 29652
rect 42924 31836 42980 31892
rect 43036 31778 43092 31780
rect 43036 31726 43038 31778
rect 43038 31726 43090 31778
rect 43090 31726 43092 31778
rect 43036 31724 43092 31726
rect 43036 30492 43092 30548
rect 43820 31890 43876 31892
rect 43820 31838 43822 31890
rect 43822 31838 43874 31890
rect 43874 31838 43876 31890
rect 43820 31836 43876 31838
rect 43932 31500 43988 31556
rect 44940 33180 44996 33236
rect 44492 32508 44548 32564
rect 44940 31890 44996 31892
rect 44940 31838 44942 31890
rect 44942 31838 44994 31890
rect 44994 31838 44996 31890
rect 44940 31836 44996 31838
rect 45388 35980 45444 36036
rect 46284 35644 46340 35700
rect 45836 35308 45892 35364
rect 45836 35084 45892 35140
rect 45500 34188 45556 34244
rect 45724 33740 45780 33796
rect 45836 34188 45892 34244
rect 45164 33404 45220 33460
rect 44268 30492 44324 30548
rect 44380 31052 44436 31108
rect 44156 30098 44212 30100
rect 44156 30046 44158 30098
rect 44158 30046 44210 30098
rect 44210 30046 44212 30098
rect 44156 30044 44212 30046
rect 43484 28812 43540 28868
rect 43484 28642 43540 28644
rect 43484 28590 43486 28642
rect 43486 28590 43538 28642
rect 43538 28590 43540 28642
rect 43484 28588 43540 28590
rect 43372 28476 43428 28532
rect 42924 27468 42980 27524
rect 42700 26572 42756 26628
rect 43260 27746 43316 27748
rect 43260 27694 43262 27746
rect 43262 27694 43314 27746
rect 43314 27694 43316 27746
rect 43260 27692 43316 27694
rect 43036 25676 43092 25732
rect 43148 26796 43204 26852
rect 42700 25564 42756 25620
rect 43260 26572 43316 26628
rect 43260 25506 43316 25508
rect 43260 25454 43262 25506
rect 43262 25454 43314 25506
rect 43314 25454 43316 25506
rect 43260 25452 43316 25454
rect 42364 24780 42420 24836
rect 42252 24722 42308 24724
rect 42252 24670 42254 24722
rect 42254 24670 42306 24722
rect 42306 24670 42308 24722
rect 42252 24668 42308 24670
rect 41132 23884 41188 23940
rect 41020 23660 41076 23716
rect 41468 23772 41524 23828
rect 40236 23436 40292 23492
rect 40348 23378 40404 23380
rect 40348 23326 40350 23378
rect 40350 23326 40402 23378
rect 40402 23326 40404 23378
rect 40348 23324 40404 23326
rect 40236 21810 40292 21812
rect 40236 21758 40238 21810
rect 40238 21758 40290 21810
rect 40290 21758 40292 21810
rect 40236 21756 40292 21758
rect 40348 21474 40404 21476
rect 40348 21422 40350 21474
rect 40350 21422 40402 21474
rect 40402 21422 40404 21474
rect 40348 21420 40404 21422
rect 41356 23378 41412 23380
rect 41356 23326 41358 23378
rect 41358 23326 41410 23378
rect 41410 23326 41412 23378
rect 41356 23324 41412 23326
rect 41804 23714 41860 23716
rect 41804 23662 41806 23714
rect 41806 23662 41858 23714
rect 41858 23662 41860 23714
rect 41804 23660 41860 23662
rect 41580 23324 41636 23380
rect 42812 25004 42868 25060
rect 42476 24668 42532 24724
rect 42364 23938 42420 23940
rect 42364 23886 42366 23938
rect 42366 23886 42418 23938
rect 42418 23886 42420 23938
rect 42364 23884 42420 23886
rect 42924 24610 42980 24612
rect 42924 24558 42926 24610
rect 42926 24558 42978 24610
rect 42978 24558 42980 24610
rect 42924 24556 42980 24558
rect 43148 24892 43204 24948
rect 43260 25004 43316 25060
rect 42140 23772 42196 23828
rect 43148 24668 43204 24724
rect 42924 23884 42980 23940
rect 42588 23714 42644 23716
rect 42588 23662 42590 23714
rect 42590 23662 42642 23714
rect 42642 23662 42644 23714
rect 42588 23660 42644 23662
rect 42028 23100 42084 23156
rect 42252 23324 42308 23380
rect 42700 23436 42756 23492
rect 44156 28476 44212 28532
rect 43932 27244 43988 27300
rect 44044 27074 44100 27076
rect 44044 27022 44046 27074
rect 44046 27022 44098 27074
rect 44098 27022 44100 27074
rect 44044 27020 44100 27022
rect 44940 30210 44996 30212
rect 44940 30158 44942 30210
rect 44942 30158 44994 30210
rect 44994 30158 44996 30210
rect 44940 30156 44996 30158
rect 44940 28754 44996 28756
rect 44940 28702 44942 28754
rect 44942 28702 44994 28754
rect 44994 28702 44996 28754
rect 44940 28700 44996 28702
rect 44828 28642 44884 28644
rect 44828 28590 44830 28642
rect 44830 28590 44882 28642
rect 44882 28590 44884 28642
rect 44828 28588 44884 28590
rect 45388 31890 45444 31892
rect 45388 31838 45390 31890
rect 45390 31838 45442 31890
rect 45442 31838 45444 31890
rect 45388 31836 45444 31838
rect 45724 31724 45780 31780
rect 45388 30210 45444 30212
rect 45388 30158 45390 30210
rect 45390 30158 45442 30210
rect 45442 30158 45444 30210
rect 45388 30156 45444 30158
rect 45388 29596 45444 29652
rect 44828 27804 44884 27860
rect 44716 27298 44772 27300
rect 44716 27246 44718 27298
rect 44718 27246 44770 27298
rect 44770 27246 44772 27298
rect 44716 27244 44772 27246
rect 44380 27020 44436 27076
rect 44268 25228 44324 25284
rect 44156 24108 44212 24164
rect 43260 23772 43316 23828
rect 42252 22316 42308 22372
rect 42364 22876 42420 22932
rect 41804 22258 41860 22260
rect 41804 22206 41806 22258
rect 41806 22206 41858 22258
rect 41858 22206 41860 22258
rect 41804 22204 41860 22206
rect 40908 21532 40964 21588
rect 40460 21084 40516 21140
rect 39676 20860 39732 20916
rect 40348 20914 40404 20916
rect 40348 20862 40350 20914
rect 40350 20862 40402 20914
rect 40402 20862 40404 20914
rect 40348 20860 40404 20862
rect 38780 20690 38836 20692
rect 38780 20638 38782 20690
rect 38782 20638 38834 20690
rect 38834 20638 38836 20690
rect 38780 20636 38836 20638
rect 38556 20076 38612 20132
rect 38220 19964 38276 20020
rect 37772 19404 37828 19460
rect 37548 19180 37604 19236
rect 37212 18620 37268 18676
rect 37100 17388 37156 17444
rect 37212 17500 37268 17556
rect 36988 16716 37044 16772
rect 37212 17052 37268 17108
rect 37436 16828 37492 16884
rect 37996 18396 38052 18452
rect 37884 17836 37940 17892
rect 38780 20018 38836 20020
rect 38780 19966 38782 20018
rect 38782 19966 38834 20018
rect 38834 19966 38836 20018
rect 38780 19964 38836 19966
rect 39116 20130 39172 20132
rect 39116 20078 39118 20130
rect 39118 20078 39170 20130
rect 39170 20078 39172 20130
rect 39116 20076 39172 20078
rect 39340 20076 39396 20132
rect 38780 19292 38836 19348
rect 39116 19292 39172 19348
rect 39004 19234 39060 19236
rect 39004 19182 39006 19234
rect 39006 19182 39058 19234
rect 39058 19182 39060 19234
rect 39004 19180 39060 19182
rect 38332 18844 38388 18900
rect 38668 18620 38724 18676
rect 38444 18396 38500 18452
rect 38332 17106 38388 17108
rect 38332 17054 38334 17106
rect 38334 17054 38386 17106
rect 38386 17054 38388 17106
rect 38332 17052 38388 17054
rect 39676 19346 39732 19348
rect 39676 19294 39678 19346
rect 39678 19294 39730 19346
rect 39730 19294 39732 19346
rect 39676 19292 39732 19294
rect 39564 19180 39620 19236
rect 39228 18620 39284 18676
rect 39340 18844 39396 18900
rect 38780 18172 38836 18228
rect 38668 17164 38724 17220
rect 38220 16940 38276 16996
rect 39788 18674 39844 18676
rect 39788 18622 39790 18674
rect 39790 18622 39842 18674
rect 39842 18622 39844 18674
rect 39788 18620 39844 18622
rect 39452 18172 39508 18228
rect 39900 16994 39956 16996
rect 39900 16942 39902 16994
rect 39902 16942 39954 16994
rect 39954 16942 39956 16994
rect 39900 16940 39956 16942
rect 38556 16882 38612 16884
rect 38556 16830 38558 16882
rect 38558 16830 38610 16882
rect 38610 16830 38612 16882
rect 38556 16828 38612 16830
rect 40012 16882 40068 16884
rect 40012 16830 40014 16882
rect 40014 16830 40066 16882
rect 40066 16830 40068 16882
rect 40012 16828 40068 16830
rect 38892 16268 38948 16324
rect 38668 15372 38724 15428
rect 36764 14700 36820 14756
rect 36428 13074 36484 13076
rect 36428 13022 36430 13074
rect 36430 13022 36482 13074
rect 36482 13022 36484 13074
rect 36428 13020 36484 13022
rect 36652 12290 36708 12292
rect 36652 12238 36654 12290
rect 36654 12238 36706 12290
rect 36706 12238 36708 12290
rect 36652 12236 36708 12238
rect 36428 12178 36484 12180
rect 36428 12126 36430 12178
rect 36430 12126 36482 12178
rect 36482 12126 36484 12178
rect 36428 12124 36484 12126
rect 36652 12012 36708 12068
rect 36540 10892 36596 10948
rect 36428 10834 36484 10836
rect 36428 10782 36430 10834
rect 36430 10782 36482 10834
rect 36482 10782 36484 10834
rect 36428 10780 36484 10782
rect 36316 10668 36372 10724
rect 37212 14364 37268 14420
rect 36988 14306 37044 14308
rect 36988 14254 36990 14306
rect 36990 14254 37042 14306
rect 37042 14254 37044 14306
rect 36988 14252 37044 14254
rect 36876 11900 36932 11956
rect 37324 11788 37380 11844
rect 37212 11676 37268 11732
rect 37548 14476 37604 14532
rect 37996 13468 38052 13524
rect 37884 13020 37940 13076
rect 37436 11564 37492 11620
rect 37548 12236 37604 12292
rect 39788 15538 39844 15540
rect 39788 15486 39790 15538
rect 39790 15486 39842 15538
rect 39842 15486 39844 15538
rect 39788 15484 39844 15486
rect 41580 21362 41636 21364
rect 41580 21310 41582 21362
rect 41582 21310 41634 21362
rect 41634 21310 41636 21362
rect 41580 21308 41636 21310
rect 40908 20748 40964 20804
rect 41356 20914 41412 20916
rect 41356 20862 41358 20914
rect 41358 20862 41410 20914
rect 41410 20862 41412 20914
rect 41356 20860 41412 20862
rect 42252 22146 42308 22148
rect 42252 22094 42254 22146
rect 42254 22094 42306 22146
rect 42306 22094 42308 22146
rect 42252 22092 42308 22094
rect 42924 22930 42980 22932
rect 42924 22878 42926 22930
rect 42926 22878 42978 22930
rect 42978 22878 42980 22930
rect 42924 22876 42980 22878
rect 42700 22370 42756 22372
rect 42700 22318 42702 22370
rect 42702 22318 42754 22370
rect 42754 22318 42756 22370
rect 42700 22316 42756 22318
rect 43372 23884 43428 23940
rect 43148 22482 43204 22484
rect 43148 22430 43150 22482
rect 43150 22430 43202 22482
rect 43202 22430 43204 22482
rect 43148 22428 43204 22430
rect 42700 21362 42756 21364
rect 42700 21310 42702 21362
rect 42702 21310 42754 21362
rect 42754 21310 42756 21362
rect 42700 21308 42756 21310
rect 42140 20860 42196 20916
rect 42476 21084 42532 21140
rect 41804 20636 41860 20692
rect 40796 19404 40852 19460
rect 40236 18844 40292 18900
rect 40908 19292 40964 19348
rect 41356 19346 41412 19348
rect 41356 19294 41358 19346
rect 41358 19294 41410 19346
rect 41410 19294 41412 19346
rect 41356 19292 41412 19294
rect 40460 18620 40516 18676
rect 40236 16716 40292 16772
rect 40796 17724 40852 17780
rect 40348 16492 40404 16548
rect 40348 16268 40404 16324
rect 41804 19292 41860 19348
rect 41356 17612 41412 17668
rect 41132 17052 41188 17108
rect 41580 17164 41636 17220
rect 42252 17052 42308 17108
rect 41468 16770 41524 16772
rect 41468 16718 41470 16770
rect 41470 16718 41522 16770
rect 41522 16718 41524 16770
rect 41468 16716 41524 16718
rect 41468 16492 41524 16548
rect 44044 23714 44100 23716
rect 44044 23662 44046 23714
rect 44046 23662 44098 23714
rect 44098 23662 44100 23714
rect 44044 23660 44100 23662
rect 44828 25730 44884 25732
rect 44828 25678 44830 25730
rect 44830 25678 44882 25730
rect 44882 25678 44884 25730
rect 44828 25676 44884 25678
rect 45052 27132 45108 27188
rect 45276 26460 45332 26516
rect 46172 35026 46228 35028
rect 46172 34974 46174 35026
rect 46174 34974 46226 35026
rect 46226 34974 46228 35026
rect 46172 34972 46228 34974
rect 46508 38780 46564 38836
rect 46060 34300 46116 34356
rect 46172 33458 46228 33460
rect 46172 33406 46174 33458
rect 46174 33406 46226 33458
rect 46226 33406 46228 33458
rect 46172 33404 46228 33406
rect 46844 40124 46900 40180
rect 46844 39340 46900 39396
rect 46620 35644 46676 35700
rect 45948 31554 46004 31556
rect 45948 31502 45950 31554
rect 45950 31502 46002 31554
rect 46002 31502 46004 31554
rect 45948 31500 46004 31502
rect 46172 30940 46228 30996
rect 45836 30492 45892 30548
rect 45836 28364 45892 28420
rect 46060 28476 46116 28532
rect 45612 27074 45668 27076
rect 45612 27022 45614 27074
rect 45614 27022 45666 27074
rect 45666 27022 45668 27074
rect 45612 27020 45668 27022
rect 46396 31500 46452 31556
rect 46060 26796 46116 26852
rect 46284 26684 46340 26740
rect 45948 26236 46004 26292
rect 45612 25618 45668 25620
rect 45612 25566 45614 25618
rect 45614 25566 45666 25618
rect 45666 25566 45668 25618
rect 45612 25564 45668 25566
rect 44940 25116 44996 25172
rect 44828 24556 44884 24612
rect 44380 23548 44436 23604
rect 44156 23324 44212 23380
rect 43820 22876 43876 22932
rect 43708 22482 43764 22484
rect 43708 22430 43710 22482
rect 43710 22430 43762 22482
rect 43762 22430 43764 22482
rect 43708 22428 43764 22430
rect 44156 21644 44212 21700
rect 44268 21532 44324 21588
rect 44044 20972 44100 21028
rect 44156 21420 44212 21476
rect 43596 20748 43652 20804
rect 43484 20690 43540 20692
rect 43484 20638 43486 20690
rect 43486 20638 43538 20690
rect 43538 20638 43540 20690
rect 43484 20636 43540 20638
rect 43372 19852 43428 19908
rect 42588 18620 42644 18676
rect 42700 18396 42756 18452
rect 42700 17164 42756 17220
rect 44156 20412 44212 20468
rect 43484 19122 43540 19124
rect 43484 19070 43486 19122
rect 43486 19070 43538 19122
rect 43538 19070 43540 19122
rect 43484 19068 43540 19070
rect 45052 23548 45108 23604
rect 46060 25506 46116 25508
rect 46060 25454 46062 25506
rect 46062 25454 46114 25506
rect 46114 25454 46116 25506
rect 46060 25452 46116 25454
rect 46060 25228 46116 25284
rect 46060 24162 46116 24164
rect 46060 24110 46062 24162
rect 46062 24110 46114 24162
rect 46114 24110 46116 24162
rect 46060 24108 46116 24110
rect 46508 28364 46564 28420
rect 46060 23154 46116 23156
rect 46060 23102 46062 23154
rect 46062 23102 46114 23154
rect 46114 23102 46116 23154
rect 46060 23100 46116 23102
rect 46172 22258 46228 22260
rect 46172 22206 46174 22258
rect 46174 22206 46226 22258
rect 46226 22206 46228 22258
rect 46172 22204 46228 22206
rect 45276 22092 45332 22148
rect 44940 21420 44996 21476
rect 45052 21868 45108 21924
rect 44940 21026 44996 21028
rect 44940 20974 44942 21026
rect 44942 20974 44994 21026
rect 44994 20974 44996 21026
rect 44940 20972 44996 20974
rect 44828 20690 44884 20692
rect 44828 20638 44830 20690
rect 44830 20638 44882 20690
rect 44882 20638 44884 20690
rect 44828 20636 44884 20638
rect 43820 18396 43876 18452
rect 44380 18172 44436 18228
rect 43484 17276 43540 17332
rect 43036 17052 43092 17108
rect 43372 17164 43428 17220
rect 42588 16770 42644 16772
rect 42588 16718 42590 16770
rect 42590 16718 42642 16770
rect 42642 16718 42644 16770
rect 42588 16716 42644 16718
rect 41804 16044 41860 16100
rect 43596 16380 43652 16436
rect 42924 15932 42980 15988
rect 43596 16044 43652 16100
rect 40236 14476 40292 14532
rect 39564 14364 39620 14420
rect 42812 15372 42868 15428
rect 41132 15148 41188 15204
rect 42700 15260 42756 15316
rect 40460 14418 40516 14420
rect 40460 14366 40462 14418
rect 40462 14366 40514 14418
rect 40514 14366 40516 14418
rect 40460 14364 40516 14366
rect 42700 14364 42756 14420
rect 41692 14252 41748 14308
rect 40236 13916 40292 13972
rect 41132 13580 41188 13636
rect 40012 13356 40068 13412
rect 37660 11788 37716 11844
rect 37660 11564 37716 11620
rect 37660 11340 37716 11396
rect 36988 10892 37044 10948
rect 37100 11228 37156 11284
rect 36540 10556 36596 10612
rect 33964 8092 34020 8148
rect 34076 7756 34132 7812
rect 33964 7586 34020 7588
rect 33964 7534 33966 7586
rect 33966 7534 34018 7586
rect 34018 7534 34020 7586
rect 33964 7532 34020 7534
rect 35756 9100 35812 9156
rect 35084 8764 35140 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34300 7644 34356 7700
rect 35084 8204 35140 8260
rect 35532 8428 35588 8484
rect 35084 7868 35140 7924
rect 35084 7644 35140 7700
rect 34524 7308 34580 7364
rect 34412 7196 34468 7252
rect 33964 6860 34020 6916
rect 33628 6636 33684 6692
rect 33852 6748 33908 6804
rect 33740 6188 33796 6244
rect 33180 5906 33236 5908
rect 33180 5854 33182 5906
rect 33182 5854 33234 5906
rect 33234 5854 33236 5906
rect 33180 5852 33236 5854
rect 32732 5516 32788 5572
rect 32284 4956 32340 5012
rect 33068 5068 33124 5124
rect 33516 4956 33572 5012
rect 34300 5852 34356 5908
rect 34300 5292 34356 5348
rect 34636 5794 34692 5796
rect 34636 5742 34638 5794
rect 34638 5742 34690 5794
rect 34690 5742 34692 5794
rect 34636 5740 34692 5742
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35308 5852 35364 5908
rect 36092 8428 36148 8484
rect 37884 11228 37940 11284
rect 37212 10892 37268 10948
rect 37324 11004 37380 11060
rect 37100 9602 37156 9604
rect 37100 9550 37102 9602
rect 37102 9550 37154 9602
rect 37154 9550 37156 9602
rect 37100 9548 37156 9550
rect 37100 8988 37156 9044
rect 37212 8258 37268 8260
rect 37212 8206 37214 8258
rect 37214 8206 37266 8258
rect 37266 8206 37268 8258
rect 37212 8204 37268 8206
rect 36092 6748 36148 6804
rect 36204 6690 36260 6692
rect 36204 6638 36206 6690
rect 36206 6638 36258 6690
rect 36258 6638 36260 6690
rect 36204 6636 36260 6638
rect 35420 5740 35476 5796
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34860 5180 34916 5236
rect 35196 5292 35252 5348
rect 34636 5068 34692 5124
rect 34524 4956 34580 5012
rect 36092 6524 36148 6580
rect 35644 5010 35700 5012
rect 35644 4958 35646 5010
rect 35646 4958 35698 5010
rect 35698 4958 35700 5010
rect 35644 4956 35700 4958
rect 35420 4898 35476 4900
rect 35420 4846 35422 4898
rect 35422 4846 35474 4898
rect 35474 4846 35476 4898
rect 35420 4844 35476 4846
rect 35980 5292 36036 5348
rect 35868 5010 35924 5012
rect 35868 4958 35870 5010
rect 35870 4958 35922 5010
rect 35922 4958 35924 5010
rect 35868 4956 35924 4958
rect 35756 4396 35812 4452
rect 27804 3388 27860 3444
rect 26236 3276 26292 3332
rect 27020 3330 27076 3332
rect 27020 3278 27022 3330
rect 27022 3278 27074 3330
rect 27074 3278 27076 3330
rect 27020 3276 27076 3278
rect 29372 3388 29428 3444
rect 32172 3554 32228 3556
rect 32172 3502 32174 3554
rect 32174 3502 32226 3554
rect 32226 3502 32228 3554
rect 32172 3500 32228 3502
rect 34748 4172 34804 4228
rect 34076 4060 34132 4116
rect 33740 3442 33796 3444
rect 33740 3390 33742 3442
rect 33742 3390 33794 3442
rect 33794 3390 33796 3442
rect 33740 3388 33796 3390
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35980 4226 36036 4228
rect 35980 4174 35982 4226
rect 35982 4174 36034 4226
rect 36034 4174 36036 4226
rect 35980 4172 36036 4174
rect 35980 3948 36036 4004
rect 35980 3724 36036 3780
rect 35196 3554 35252 3556
rect 35196 3502 35198 3554
rect 35198 3502 35250 3554
rect 35250 3502 35252 3554
rect 35196 3500 35252 3502
rect 37436 9996 37492 10052
rect 37548 10556 37604 10612
rect 37436 9548 37492 9604
rect 38220 11676 38276 11732
rect 38332 11340 38388 11396
rect 37660 10498 37716 10500
rect 37660 10446 37662 10498
rect 37662 10446 37714 10498
rect 37714 10446 37716 10498
rect 37660 10444 37716 10446
rect 38220 11116 38276 11172
rect 38780 11340 38836 11396
rect 39228 11676 39284 11732
rect 39116 11564 39172 11620
rect 38668 11228 38724 11284
rect 38780 11004 38836 11060
rect 39452 12908 39508 12964
rect 39788 12738 39844 12740
rect 39788 12686 39790 12738
rect 39790 12686 39842 12738
rect 39842 12686 39844 12738
rect 39788 12684 39844 12686
rect 39452 11394 39508 11396
rect 39452 11342 39454 11394
rect 39454 11342 39506 11394
rect 39506 11342 39508 11394
rect 39452 11340 39508 11342
rect 39340 11004 39396 11060
rect 39452 10834 39508 10836
rect 39452 10782 39454 10834
rect 39454 10782 39506 10834
rect 39506 10782 39508 10834
rect 39452 10780 39508 10782
rect 37884 9602 37940 9604
rect 37884 9550 37886 9602
rect 37886 9550 37938 9602
rect 37938 9550 37940 9602
rect 37884 9548 37940 9550
rect 37772 8988 37828 9044
rect 38332 8988 38388 9044
rect 37660 8876 37716 8932
rect 37884 8540 37940 8596
rect 37436 7644 37492 7700
rect 37324 7420 37380 7476
rect 36428 6860 36484 6916
rect 36316 6076 36372 6132
rect 37212 6412 37268 6468
rect 36204 5740 36260 5796
rect 36316 5234 36372 5236
rect 36316 5182 36318 5234
rect 36318 5182 36370 5234
rect 36370 5182 36372 5234
rect 36316 5180 36372 5182
rect 36204 5068 36260 5124
rect 36988 5122 37044 5124
rect 36988 5070 36990 5122
rect 36990 5070 37042 5122
rect 37042 5070 37044 5122
rect 36988 5068 37044 5070
rect 37100 4450 37156 4452
rect 37100 4398 37102 4450
rect 37102 4398 37154 4450
rect 37154 4398 37156 4450
rect 37100 4396 37156 4398
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 36428 3388 36484 3444
rect 37772 6578 37828 6580
rect 37772 6526 37774 6578
rect 37774 6526 37826 6578
rect 37826 6526 37828 6578
rect 37772 6524 37828 6526
rect 39564 10610 39620 10612
rect 39564 10558 39566 10610
rect 39566 10558 39618 10610
rect 39618 10558 39620 10610
rect 39564 10556 39620 10558
rect 38892 9996 38948 10052
rect 39004 10108 39060 10164
rect 38892 9826 38948 9828
rect 38892 9774 38894 9826
rect 38894 9774 38946 9826
rect 38946 9774 38948 9826
rect 38892 9772 38948 9774
rect 39004 9436 39060 9492
rect 38892 8482 38948 8484
rect 38892 8430 38894 8482
rect 38894 8430 38946 8482
rect 38946 8430 38948 8482
rect 38892 8428 38948 8430
rect 38780 8258 38836 8260
rect 38780 8206 38782 8258
rect 38782 8206 38834 8258
rect 38834 8206 38836 8258
rect 38780 8204 38836 8206
rect 38556 7868 38612 7924
rect 39452 9884 39508 9940
rect 40684 12962 40740 12964
rect 40684 12910 40686 12962
rect 40686 12910 40738 12962
rect 40738 12910 40740 12962
rect 40684 12908 40740 12910
rect 41916 13804 41972 13860
rect 41468 13746 41524 13748
rect 41468 13694 41470 13746
rect 41470 13694 41522 13746
rect 41522 13694 41524 13746
rect 41468 13692 41524 13694
rect 41804 13692 41860 13748
rect 41692 13580 41748 13636
rect 40124 11452 40180 11508
rect 39676 9660 39732 9716
rect 40236 11340 40292 11396
rect 39564 9548 39620 9604
rect 39116 8988 39172 9044
rect 39004 7756 39060 7812
rect 39340 9266 39396 9268
rect 39340 9214 39342 9266
rect 39342 9214 39394 9266
rect 39394 9214 39396 9266
rect 39340 9212 39396 9214
rect 39900 10892 39956 10948
rect 40012 9996 40068 10052
rect 39900 9772 39956 9828
rect 40348 10556 40404 10612
rect 40124 9772 40180 9828
rect 40012 9660 40068 9716
rect 40460 9826 40516 9828
rect 40460 9774 40462 9826
rect 40462 9774 40514 9826
rect 40514 9774 40516 9826
rect 40460 9772 40516 9774
rect 39788 8930 39844 8932
rect 39788 8878 39790 8930
rect 39790 8878 39842 8930
rect 39842 8878 39844 8930
rect 39788 8876 39844 8878
rect 40236 9212 40292 9268
rect 40012 8876 40068 8932
rect 40124 8764 40180 8820
rect 39228 7532 39284 7588
rect 39676 8204 39732 8260
rect 39788 7868 39844 7924
rect 37996 6972 38052 7028
rect 37884 5404 37940 5460
rect 37772 5292 37828 5348
rect 37660 5068 37716 5124
rect 38332 4732 38388 4788
rect 38444 6972 38500 7028
rect 39564 7420 39620 7476
rect 39340 7362 39396 7364
rect 39340 7310 39342 7362
rect 39342 7310 39394 7362
rect 39394 7310 39396 7362
rect 39340 7308 39396 7310
rect 39228 7250 39284 7252
rect 39228 7198 39230 7250
rect 39230 7198 39282 7250
rect 39282 7198 39284 7250
rect 39228 7196 39284 7198
rect 38892 6972 38948 7028
rect 39452 6300 39508 6356
rect 39228 5740 39284 5796
rect 39452 5964 39508 6020
rect 38780 4844 38836 4900
rect 39228 4844 39284 4900
rect 38892 4732 38948 4788
rect 38892 3948 38948 4004
rect 39228 3948 39284 4004
rect 39900 7586 39956 7588
rect 39900 7534 39902 7586
rect 39902 7534 39954 7586
rect 39954 7534 39956 7586
rect 39900 7532 39956 7534
rect 39788 6636 39844 6692
rect 41020 11116 41076 11172
rect 40796 10780 40852 10836
rect 41244 11676 41300 11732
rect 41356 11506 41412 11508
rect 41356 11454 41358 11506
rect 41358 11454 41410 11506
rect 41410 11454 41412 11506
rect 41356 11452 41412 11454
rect 41580 11788 41636 11844
rect 42364 13746 42420 13748
rect 42364 13694 42366 13746
rect 42366 13694 42418 13746
rect 42418 13694 42420 13746
rect 42364 13692 42420 13694
rect 42140 13468 42196 13524
rect 42476 12962 42532 12964
rect 42476 12910 42478 12962
rect 42478 12910 42530 12962
rect 42530 12910 42532 12962
rect 42476 12908 42532 12910
rect 41916 11676 41972 11732
rect 40796 9660 40852 9716
rect 40684 9602 40740 9604
rect 40684 9550 40686 9602
rect 40686 9550 40738 9602
rect 40738 9550 40740 9602
rect 40684 9548 40740 9550
rect 40908 8764 40964 8820
rect 41132 9436 41188 9492
rect 41916 11394 41972 11396
rect 41916 11342 41918 11394
rect 41918 11342 41970 11394
rect 41970 11342 41972 11394
rect 41916 11340 41972 11342
rect 42028 11116 42084 11172
rect 42140 10556 42196 10612
rect 42028 9884 42084 9940
rect 42476 11394 42532 11396
rect 42476 11342 42478 11394
rect 42478 11342 42530 11394
rect 42530 11342 42532 11394
rect 42476 11340 42532 11342
rect 42364 11116 42420 11172
rect 42252 10220 42308 10276
rect 42364 10780 42420 10836
rect 42924 14364 42980 14420
rect 43036 13580 43092 13636
rect 43372 15260 43428 15316
rect 43148 13356 43204 13412
rect 42812 13020 42868 13076
rect 43148 12962 43204 12964
rect 43148 12910 43150 12962
rect 43150 12910 43202 12962
rect 43202 12910 43204 12962
rect 43148 12908 43204 12910
rect 42700 11228 42756 11284
rect 42588 10610 42644 10612
rect 42588 10558 42590 10610
rect 42590 10558 42642 10610
rect 42642 10558 42644 10610
rect 42588 10556 42644 10558
rect 44044 15986 44100 15988
rect 44044 15934 44046 15986
rect 44046 15934 44098 15986
rect 44098 15934 44100 15986
rect 44044 15932 44100 15934
rect 43708 15260 43764 15316
rect 45164 21308 45220 21364
rect 46172 21980 46228 22036
rect 45388 21698 45444 21700
rect 45388 21646 45390 21698
rect 45390 21646 45442 21698
rect 45442 21646 45444 21698
rect 45388 21644 45444 21646
rect 46060 21586 46116 21588
rect 46060 21534 46062 21586
rect 46062 21534 46114 21586
rect 46114 21534 46116 21586
rect 46060 21532 46116 21534
rect 46284 21532 46340 21588
rect 45276 19458 45332 19460
rect 45276 19406 45278 19458
rect 45278 19406 45330 19458
rect 45330 19406 45332 19458
rect 45276 19404 45332 19406
rect 45164 19234 45220 19236
rect 45164 19182 45166 19234
rect 45166 19182 45218 19234
rect 45218 19182 45220 19234
rect 45164 19180 45220 19182
rect 44828 19122 44884 19124
rect 44828 19070 44830 19122
rect 44830 19070 44882 19122
rect 44882 19070 44884 19122
rect 44828 19068 44884 19070
rect 45164 18396 45220 18452
rect 44940 18284 44996 18340
rect 45948 19292 46004 19348
rect 45836 19234 45892 19236
rect 45836 19182 45838 19234
rect 45838 19182 45890 19234
rect 45890 19182 45892 19234
rect 45836 19180 45892 19182
rect 45612 18226 45668 18228
rect 45612 18174 45614 18226
rect 45614 18174 45666 18226
rect 45666 18174 45668 18226
rect 45612 18172 45668 18174
rect 45388 18060 45444 18116
rect 44940 17778 44996 17780
rect 44940 17726 44942 17778
rect 44942 17726 44994 17778
rect 44994 17726 44996 17778
rect 44940 17724 44996 17726
rect 45388 17778 45444 17780
rect 45388 17726 45390 17778
rect 45390 17726 45442 17778
rect 45442 17726 45444 17778
rect 45388 17724 45444 17726
rect 44828 17164 44884 17220
rect 44828 16716 44884 16772
rect 46172 18338 46228 18340
rect 46172 18286 46174 18338
rect 46174 18286 46226 18338
rect 46226 18286 46228 18338
rect 46172 18284 46228 18286
rect 45836 17442 45892 17444
rect 45836 17390 45838 17442
rect 45838 17390 45890 17442
rect 45890 17390 45892 17442
rect 45836 17388 45892 17390
rect 45276 16210 45332 16212
rect 45276 16158 45278 16210
rect 45278 16158 45330 16210
rect 45330 16158 45332 16210
rect 45276 16156 45332 16158
rect 46172 18060 46228 18116
rect 46620 24444 46676 24500
rect 46844 21980 46900 22036
rect 46508 17724 46564 17780
rect 46060 17164 46116 17220
rect 44156 15484 44212 15540
rect 43708 14418 43764 14420
rect 43708 14366 43710 14418
rect 43710 14366 43762 14418
rect 43762 14366 43764 14418
rect 43708 14364 43764 14366
rect 43596 13356 43652 13412
rect 43484 13020 43540 13076
rect 43708 12962 43764 12964
rect 43708 12910 43710 12962
rect 43710 12910 43762 12962
rect 43762 12910 43764 12962
rect 43708 12908 43764 12910
rect 43484 12124 43540 12180
rect 43820 11676 43876 11732
rect 43372 11564 43428 11620
rect 43036 11394 43092 11396
rect 43036 11342 43038 11394
rect 43038 11342 43090 11394
rect 43090 11342 43092 11394
rect 43036 11340 43092 11342
rect 42812 9996 42868 10052
rect 42924 11116 42980 11172
rect 43260 11004 43316 11060
rect 41356 9436 41412 9492
rect 41804 9212 41860 9268
rect 41916 9602 41972 9604
rect 41916 9550 41918 9602
rect 41918 9550 41970 9602
rect 41970 9550 41972 9602
rect 41916 9548 41972 9550
rect 41468 8988 41524 9044
rect 40572 7308 40628 7364
rect 41244 8092 41300 8148
rect 41132 7868 41188 7924
rect 41020 7084 41076 7140
rect 40460 6748 40516 6804
rect 40460 6188 40516 6244
rect 40684 6412 40740 6468
rect 40908 6690 40964 6692
rect 40908 6638 40910 6690
rect 40910 6638 40962 6690
rect 40962 6638 40964 6690
rect 40908 6636 40964 6638
rect 41020 6524 41076 6580
rect 40348 6018 40404 6020
rect 40348 5966 40350 6018
rect 40350 5966 40402 6018
rect 40402 5966 40404 6018
rect 40348 5964 40404 5966
rect 40124 5852 40180 5908
rect 41020 6130 41076 6132
rect 41020 6078 41022 6130
rect 41022 6078 41074 6130
rect 41074 6078 41076 6130
rect 41020 6076 41076 6078
rect 41356 6860 41412 6916
rect 41468 7756 41524 7812
rect 40908 5964 40964 6020
rect 41692 7084 41748 7140
rect 41580 6636 41636 6692
rect 40796 5740 40852 5796
rect 40572 5292 40628 5348
rect 38444 3388 38500 3444
rect 38780 3612 38836 3668
rect 40012 4172 40068 4228
rect 42028 6972 42084 7028
rect 41916 6076 41972 6132
rect 41692 5906 41748 5908
rect 41692 5854 41694 5906
rect 41694 5854 41746 5906
rect 41746 5854 41748 5906
rect 41692 5852 41748 5854
rect 41916 4844 41972 4900
rect 40796 4172 40852 4228
rect 41580 4226 41636 4228
rect 41580 4174 41582 4226
rect 41582 4174 41634 4226
rect 41634 4174 41636 4226
rect 41580 4172 41636 4174
rect 40348 3836 40404 3892
rect 39564 3500 39620 3556
rect 39116 3442 39172 3444
rect 39116 3390 39118 3442
rect 39118 3390 39170 3442
rect 39170 3390 39172 3442
rect 39116 3388 39172 3390
rect 42140 6578 42196 6580
rect 42140 6526 42142 6578
rect 42142 6526 42194 6578
rect 42194 6526 42196 6578
rect 42140 6524 42196 6526
rect 42252 6188 42308 6244
rect 42364 6860 42420 6916
rect 42364 6412 42420 6468
rect 42140 5906 42196 5908
rect 42140 5854 42142 5906
rect 42142 5854 42194 5906
rect 42194 5854 42196 5906
rect 42140 5852 42196 5854
rect 42252 4956 42308 5012
rect 42476 4450 42532 4452
rect 42476 4398 42478 4450
rect 42478 4398 42530 4450
rect 42530 4398 42532 4450
rect 42476 4396 42532 4398
rect 43036 9100 43092 9156
rect 42924 8204 42980 8260
rect 42812 6860 42868 6916
rect 42812 6690 42868 6692
rect 42812 6638 42814 6690
rect 42814 6638 42866 6690
rect 42866 6638 42868 6690
rect 42812 6636 42868 6638
rect 42924 6578 42980 6580
rect 42924 6526 42926 6578
rect 42926 6526 42978 6578
rect 42978 6526 42980 6578
rect 42924 6524 42980 6526
rect 42812 5794 42868 5796
rect 42812 5742 42814 5794
rect 42814 5742 42866 5794
rect 42866 5742 42868 5794
rect 42812 5740 42868 5742
rect 43820 11394 43876 11396
rect 43820 11342 43822 11394
rect 43822 11342 43874 11394
rect 43874 11342 43876 11394
rect 43820 11340 43876 11342
rect 43260 8428 43316 8484
rect 44044 12908 44100 12964
rect 44716 12348 44772 12404
rect 44044 11228 44100 11284
rect 43596 9602 43652 9604
rect 43596 9550 43598 9602
rect 43598 9550 43650 9602
rect 43650 9550 43652 9602
rect 43596 9548 43652 9550
rect 43484 7308 43540 7364
rect 43708 6914 43764 6916
rect 43708 6862 43710 6914
rect 43710 6862 43762 6914
rect 43762 6862 43764 6914
rect 43708 6860 43764 6862
rect 43484 5234 43540 5236
rect 43484 5182 43486 5234
rect 43486 5182 43538 5234
rect 43538 5182 43540 5234
rect 43484 5180 43540 5182
rect 43372 5068 43428 5124
rect 42700 4172 42756 4228
rect 42812 3948 42868 4004
rect 42924 3836 42980 3892
rect 43260 4226 43316 4228
rect 43260 4174 43262 4226
rect 43262 4174 43314 4226
rect 43314 4174 43316 4226
rect 43260 4172 43316 4174
rect 43708 3554 43764 3556
rect 43708 3502 43710 3554
rect 43710 3502 43762 3554
rect 43762 3502 43764 3554
rect 43708 3500 43764 3502
rect 43932 9436 43988 9492
rect 43932 8428 43988 8484
rect 44268 8316 44324 8372
rect 43932 6972 43988 7028
rect 44044 7644 44100 7700
rect 44156 6914 44212 6916
rect 44156 6862 44158 6914
rect 44158 6862 44210 6914
rect 44210 6862 44212 6914
rect 44156 6860 44212 6862
rect 44044 6466 44100 6468
rect 44044 6414 44046 6466
rect 44046 6414 44098 6466
rect 44098 6414 44100 6466
rect 44044 6412 44100 6414
rect 44268 5122 44324 5124
rect 44268 5070 44270 5122
rect 44270 5070 44322 5122
rect 44322 5070 44324 5122
rect 44268 5068 44324 5070
rect 44492 12124 44548 12180
rect 44828 9602 44884 9604
rect 44828 9550 44830 9602
rect 44830 9550 44882 9602
rect 44882 9550 44884 9602
rect 44828 9548 44884 9550
rect 45948 15148 46004 15204
rect 45276 12908 45332 12964
rect 45164 12348 45220 12404
rect 45052 8258 45108 8260
rect 45052 8206 45054 8258
rect 45054 8206 45106 8258
rect 45106 8206 45108 8258
rect 45052 8204 45108 8206
rect 44716 7474 44772 7476
rect 44716 7422 44718 7474
rect 44718 7422 44770 7474
rect 44770 7422 44772 7474
rect 44716 7420 44772 7422
rect 45052 6802 45108 6804
rect 45052 6750 45054 6802
rect 45054 6750 45106 6802
rect 45106 6750 45108 6802
rect 45052 6748 45108 6750
rect 45388 8258 45444 8260
rect 45388 8206 45390 8258
rect 45390 8206 45442 8258
rect 45442 8206 45444 8258
rect 45388 8204 45444 8206
rect 45276 6972 45332 7028
rect 45500 6914 45556 6916
rect 45500 6862 45502 6914
rect 45502 6862 45554 6914
rect 45554 6862 45556 6914
rect 45500 6860 45556 6862
rect 45836 13132 45892 13188
rect 46284 16828 46340 16884
rect 46060 12460 46116 12516
rect 45836 10668 45892 10724
rect 45836 9602 45892 9604
rect 45836 9550 45838 9602
rect 45838 9550 45890 9602
rect 45890 9550 45892 9602
rect 45836 9548 45892 9550
rect 46172 9100 46228 9156
rect 44940 5740 44996 5796
rect 44380 4956 44436 5012
rect 44604 4060 44660 4116
rect 44828 5292 44884 5348
rect 45052 4396 45108 4452
rect 46060 8316 46116 8372
rect 45948 8258 46004 8260
rect 45948 8206 45950 8258
rect 45950 8206 46002 8258
rect 46002 8206 46004 8258
rect 45948 8204 46004 8206
rect 45948 6412 46004 6468
rect 46060 6300 46116 6356
rect 46284 7980 46340 8036
rect 45836 4844 45892 4900
rect 43372 2716 43428 2772
<< metal3 >>
rect 47200 45108 48000 45136
rect 42914 45052 42924 45108
rect 42980 45052 48000 45108
rect 47200 45024 48000 45052
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 14588 44492 20188 44548
rect 14588 44436 14644 44492
rect 20132 44436 20188 44492
rect 14578 44380 14588 44436
rect 14644 44380 14654 44436
rect 15586 44380 15596 44436
rect 15652 44380 18172 44436
rect 18228 44380 18238 44436
rect 20132 44380 20412 44436
rect 20468 44380 20478 44436
rect 21532 44380 21980 44436
rect 22036 44380 22046 44436
rect 39218 44380 39228 44436
rect 39284 44380 39294 44436
rect 43026 44380 43036 44436
rect 43092 44380 45164 44436
rect 45220 44380 45230 44436
rect 21532 44324 21588 44380
rect 39228 44324 39284 44380
rect 17490 44268 17500 44324
rect 17556 44268 21588 44324
rect 21746 44268 21756 44324
rect 21812 44268 22428 44324
rect 22484 44268 22764 44324
rect 22820 44268 22830 44324
rect 30566 44268 30604 44324
rect 30660 44268 30670 44324
rect 39228 44268 44156 44324
rect 44212 44268 44222 44324
rect 20178 44156 20188 44212
rect 20244 44156 21868 44212
rect 21924 44156 21934 44212
rect 33506 44156 33516 44212
rect 33572 44156 34860 44212
rect 34916 44156 34926 44212
rect 37090 44156 37100 44212
rect 37156 44156 41468 44212
rect 41524 44156 41534 44212
rect 41692 44156 43596 44212
rect 43652 44156 43662 44212
rect 41692 44100 41748 44156
rect 11890 44044 11900 44100
rect 11956 44044 13804 44100
rect 13860 44044 13870 44100
rect 19842 44044 19852 44100
rect 19908 44044 20244 44100
rect 20402 44044 20412 44100
rect 20468 44044 20860 44100
rect 20916 44044 20926 44100
rect 22082 44044 22092 44100
rect 22148 44044 23100 44100
rect 23156 44044 23166 44100
rect 34178 44044 34188 44100
rect 34244 44044 35868 44100
rect 35924 44044 35934 44100
rect 40450 44044 40460 44100
rect 40516 44044 41748 44100
rect 42354 44044 42364 44100
rect 42420 44044 44380 44100
rect 44436 44044 44446 44100
rect 45602 44044 45612 44100
rect 45668 44044 45678 44100
rect 20188 43988 20244 44044
rect 45612 43988 45668 44044
rect 20188 43932 22652 43988
rect 22708 43932 22718 43988
rect 33394 43932 33404 43988
rect 33460 43932 33964 43988
rect 34020 43932 39228 43988
rect 39284 43932 39900 43988
rect 39956 43932 39966 43988
rect 41346 43932 41356 43988
rect 41412 43932 45668 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 9538 43820 9548 43876
rect 9604 43820 10108 43876
rect 10164 43820 17948 43876
rect 18004 43820 18014 43876
rect 21970 43820 21980 43876
rect 22036 43820 28476 43876
rect 28532 43820 28542 43876
rect 36418 43820 36428 43876
rect 36484 43820 37324 43876
rect 37380 43820 40124 43876
rect 40180 43820 40190 43876
rect 42242 43820 42252 43876
rect 42308 43820 43708 43876
rect 43764 43820 43774 43876
rect 15138 43708 15148 43764
rect 15204 43708 19292 43764
rect 19348 43708 19358 43764
rect 22418 43708 22428 43764
rect 22484 43708 23212 43764
rect 23268 43708 23278 43764
rect 27794 43708 27804 43764
rect 27860 43708 29148 43764
rect 29204 43708 29214 43764
rect 31042 43708 31052 43764
rect 31108 43708 31836 43764
rect 31892 43708 31902 43764
rect 43138 43708 43148 43764
rect 43204 43708 44940 43764
rect 44996 43708 45006 43764
rect 21074 43596 21084 43652
rect 21140 43596 23548 43652
rect 23604 43596 23614 43652
rect 29474 43596 29484 43652
rect 29540 43596 30268 43652
rect 30324 43596 30334 43652
rect 32610 43596 32620 43652
rect 32676 43596 41692 43652
rect 41748 43596 45948 43652
rect 46004 43596 46014 43652
rect 24994 43484 25004 43540
rect 25060 43484 25676 43540
rect 25732 43484 25742 43540
rect 28690 43484 28700 43540
rect 28756 43484 29596 43540
rect 29652 43484 29662 43540
rect 39106 43484 39116 43540
rect 39172 43484 41244 43540
rect 41300 43484 41310 43540
rect 42130 43484 42140 43540
rect 42196 43484 43148 43540
rect 43204 43484 43214 43540
rect 43922 43484 43932 43540
rect 43988 43484 44268 43540
rect 44324 43484 44334 43540
rect 15922 43372 15932 43428
rect 15988 43372 16828 43428
rect 16884 43372 16894 43428
rect 19170 43372 19180 43428
rect 19236 43372 21644 43428
rect 21700 43372 22540 43428
rect 22596 43372 22606 43428
rect 26450 43372 26460 43428
rect 26516 43372 31388 43428
rect 31444 43372 31454 43428
rect 32834 43372 32844 43428
rect 32900 43372 35196 43428
rect 35252 43372 35262 43428
rect 35634 43372 35644 43428
rect 35700 43372 37100 43428
rect 37156 43372 37166 43428
rect 37986 43372 37996 43428
rect 38052 43372 39676 43428
rect 39732 43372 39742 43428
rect 41010 43372 41020 43428
rect 41076 43372 43596 43428
rect 43652 43372 44492 43428
rect 44548 43372 44558 43428
rect 41020 43316 41076 43372
rect 30146 43260 30156 43316
rect 30212 43260 30492 43316
rect 30548 43260 30716 43316
rect 30772 43260 31276 43316
rect 31332 43260 31342 43316
rect 39554 43260 39564 43316
rect 39620 43260 41076 43316
rect 41682 43260 41692 43316
rect 41748 43260 42476 43316
rect 42532 43260 42542 43316
rect 25778 43148 25788 43204
rect 25844 43148 31052 43204
rect 31108 43148 31118 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 10098 43036 10108 43092
rect 10164 43036 11732 43092
rect 36306 43036 36316 43092
rect 36372 43036 39452 43092
rect 39508 43036 39518 43092
rect 11676 42980 11732 43036
rect 6626 42924 6636 42980
rect 6692 42924 11004 42980
rect 11060 42924 11070 42980
rect 11666 42924 11676 42980
rect 11732 42924 13468 42980
rect 13524 42924 13534 42980
rect 20066 42924 20076 42980
rect 20132 42924 21868 42980
rect 21924 42924 21934 42980
rect 23426 42924 23436 42980
rect 23492 42924 26684 42980
rect 26740 42924 26750 42980
rect 34850 42924 34860 42980
rect 34916 42924 38444 42980
rect 38500 42924 38510 42980
rect 40114 42924 40124 42980
rect 40180 42924 42924 42980
rect 42980 42924 42990 42980
rect 29250 42812 29260 42868
rect 29316 42812 32284 42868
rect 32340 42812 32956 42868
rect 33012 42812 33022 42868
rect 42802 42812 42812 42868
rect 42868 42812 43484 42868
rect 43540 42812 45276 42868
rect 45332 42812 45342 42868
rect 9650 42700 9660 42756
rect 9716 42700 10892 42756
rect 10948 42700 11452 42756
rect 11508 42700 12460 42756
rect 12516 42700 12526 42756
rect 13906 42700 13916 42756
rect 13972 42700 14364 42756
rect 14420 42700 15148 42756
rect 15204 42700 15214 42756
rect 15810 42700 15820 42756
rect 15876 42700 18396 42756
rect 18452 42700 21980 42756
rect 22036 42700 22046 42756
rect 23202 42700 23212 42756
rect 23268 42700 26348 42756
rect 26404 42700 26414 42756
rect 29810 42700 29820 42756
rect 29876 42700 30044 42756
rect 30100 42700 30716 42756
rect 30772 42700 30782 42756
rect 33394 42700 33404 42756
rect 33460 42700 34188 42756
rect 34244 42700 34636 42756
rect 34692 42700 34702 42756
rect 36082 42700 36092 42756
rect 36148 42700 41132 42756
rect 41188 42700 41198 42756
rect 6626 42588 6636 42644
rect 6692 42588 9548 42644
rect 9604 42588 9614 42644
rect 12898 42588 12908 42644
rect 12964 42588 13692 42644
rect 13748 42588 14028 42644
rect 14084 42588 14094 42644
rect 24658 42588 24668 42644
rect 24724 42588 26124 42644
rect 26180 42588 26190 42644
rect 28466 42588 28476 42644
rect 28532 42588 32508 42644
rect 32564 42588 32574 42644
rect 34402 42588 34412 42644
rect 34468 42588 40124 42644
rect 40180 42588 40190 42644
rect 44258 42588 44268 42644
rect 44324 42588 44828 42644
rect 44884 42588 44894 42644
rect 18162 42476 18172 42532
rect 18228 42476 24220 42532
rect 24276 42476 24780 42532
rect 24836 42476 28140 42532
rect 28196 42476 28206 42532
rect 28914 42476 28924 42532
rect 28980 42476 30156 42532
rect 30212 42476 31500 42532
rect 31556 42476 31948 42532
rect 32004 42476 33068 42532
rect 33124 42476 34748 42532
rect 34804 42476 34814 42532
rect 37874 42476 37884 42532
rect 37940 42476 41692 42532
rect 41748 42476 41758 42532
rect 43810 42476 43820 42532
rect 43876 42476 44156 42532
rect 44212 42476 46060 42532
rect 46116 42476 46126 42532
rect 17266 42364 17276 42420
rect 17332 42364 19180 42420
rect 19236 42364 19246 42420
rect 26562 42364 26572 42420
rect 26628 42364 28700 42420
rect 28756 42364 28766 42420
rect 33394 42364 33404 42420
rect 33460 42364 33852 42420
rect 33908 42364 36316 42420
rect 36372 42364 36382 42420
rect 36642 42364 36652 42420
rect 36708 42364 37548 42420
rect 37604 42364 43148 42420
rect 43204 42364 44940 42420
rect 44996 42364 45006 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 30258 42252 30268 42308
rect 30324 42252 32396 42308
rect 32452 42252 33180 42308
rect 33236 42252 35532 42308
rect 35588 42252 35598 42308
rect 43474 42252 43484 42308
rect 43540 42252 43820 42308
rect 43876 42252 43886 42308
rect 44594 42252 44604 42308
rect 44660 42252 46284 42308
rect 46340 42252 46350 42308
rect 43698 42140 43708 42196
rect 43764 42140 45164 42196
rect 45220 42140 45230 42196
rect 45490 42140 45500 42196
rect 45556 42140 45566 42196
rect 45500 42084 45556 42140
rect 9314 42028 9324 42084
rect 9380 42028 10556 42084
rect 10612 42028 10622 42084
rect 16268 42028 16828 42084
rect 16884 42028 17500 42084
rect 17556 42028 17566 42084
rect 35634 42028 35644 42084
rect 35700 42028 36204 42084
rect 36260 42028 36270 42084
rect 43586 42028 43596 42084
rect 43652 42028 44604 42084
rect 44660 42028 44670 42084
rect 44940 42028 45556 42084
rect 13682 41804 13692 41860
rect 13748 41804 14924 41860
rect 14980 41804 14990 41860
rect 16268 41748 16324 42028
rect 18050 41916 18060 41972
rect 18116 41916 24444 41972
rect 24500 41916 24510 41972
rect 29922 41916 29932 41972
rect 29988 41916 31164 41972
rect 31220 41916 31230 41972
rect 37090 41916 37100 41972
rect 37156 41916 40012 41972
rect 40068 41916 40078 41972
rect 41906 41916 41916 41972
rect 41972 41916 44716 41972
rect 44772 41916 44782 41972
rect 44940 41860 44996 42028
rect 33170 41804 33180 41860
rect 33236 41804 35196 41860
rect 35252 41804 35262 41860
rect 36418 41804 36428 41860
rect 36484 41804 36988 41860
rect 37044 41804 38556 41860
rect 38612 41804 38622 41860
rect 40338 41804 40348 41860
rect 40404 41804 43484 41860
rect 43540 41804 44996 41860
rect 16258 41692 16268 41748
rect 16324 41692 16334 41748
rect 18050 41692 18060 41748
rect 18116 41692 19292 41748
rect 19348 41692 19358 41748
rect 33058 41692 33068 41748
rect 33124 41692 34972 41748
rect 35028 41692 35038 41748
rect 15474 41580 15484 41636
rect 15540 41580 17388 41636
rect 17444 41580 18396 41636
rect 18452 41580 18462 41636
rect 43922 41580 43932 41636
rect 43988 41580 45388 41636
rect 45444 41580 45454 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 16156 41524 16212 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 16146 41468 16156 41524
rect 16212 41468 16222 41524
rect 17826 41356 17836 41412
rect 17892 41356 18396 41412
rect 18452 41356 18462 41412
rect 25330 41356 25340 41412
rect 25396 41356 27132 41412
rect 27188 41356 27198 41412
rect 30034 41356 30044 41412
rect 30100 41356 30716 41412
rect 30772 41356 30782 41412
rect 31378 41356 31388 41412
rect 31444 41356 32172 41412
rect 32228 41356 32732 41412
rect 32788 41356 33292 41412
rect 33348 41356 33358 41412
rect 43922 41356 43932 41412
rect 43988 41356 45164 41412
rect 45220 41356 45230 41412
rect 12786 41244 12796 41300
rect 12852 41244 14700 41300
rect 14756 41244 18060 41300
rect 18116 41244 18126 41300
rect 28130 41244 28140 41300
rect 28196 41244 30268 41300
rect 30324 41244 30334 41300
rect 35970 41244 35980 41300
rect 36036 41244 36540 41300
rect 36596 41244 37212 41300
rect 37268 41244 37278 41300
rect 41458 41244 41468 41300
rect 41524 41244 45836 41300
rect 45892 41244 45902 41300
rect 6066 41132 6076 41188
rect 6132 41132 10108 41188
rect 10164 41132 10668 41188
rect 10724 41132 11788 41188
rect 11844 41132 11854 41188
rect 15586 41132 15596 41188
rect 15652 41132 16492 41188
rect 16548 41132 16558 41188
rect 18162 41132 18172 41188
rect 18228 41132 20412 41188
rect 20468 41132 20478 41188
rect 24210 41132 24220 41188
rect 24276 41132 24556 41188
rect 24612 41132 25340 41188
rect 25396 41132 28028 41188
rect 28084 41132 28094 41188
rect 30492 41132 33852 41188
rect 33908 41132 33918 41188
rect 38210 41132 38220 41188
rect 38276 41132 44828 41188
rect 44884 41132 44894 41188
rect 45938 41132 45948 41188
rect 46004 41132 46014 41188
rect 30492 41076 30548 41132
rect 45948 41076 46004 41132
rect 11442 41020 11452 41076
rect 11508 41020 14028 41076
rect 14084 41020 14094 41076
rect 21410 41020 21420 41076
rect 21476 41020 23436 41076
rect 23492 41020 23502 41076
rect 26852 41020 30548 41076
rect 30706 41020 30716 41076
rect 30772 41020 31948 41076
rect 32004 41020 32014 41076
rect 44706 41020 44716 41076
rect 44772 41020 45612 41076
rect 45668 41020 46004 41076
rect 20850 40908 20860 40964
rect 20916 40908 22876 40964
rect 22932 40908 22942 40964
rect 26852 40852 26908 41020
rect 27682 40908 27692 40964
rect 27748 40908 28476 40964
rect 28532 40908 28542 40964
rect 29698 40908 29708 40964
rect 29764 40908 31276 40964
rect 31332 40908 31342 40964
rect 34150 40908 34188 40964
rect 34244 40908 34254 40964
rect 38882 40908 38892 40964
rect 38948 40908 45948 40964
rect 46004 40908 46014 40964
rect 22978 40796 22988 40852
rect 23044 40796 26908 40852
rect 30492 40796 31164 40852
rect 31220 40796 31230 40852
rect 35186 40796 35196 40852
rect 35252 40796 43708 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 30492 40740 30548 40796
rect 43652 40740 43708 40796
rect 22866 40684 22876 40740
rect 22932 40684 24332 40740
rect 24388 40684 24398 40740
rect 28466 40684 28476 40740
rect 28532 40684 30492 40740
rect 30548 40684 30558 40740
rect 30706 40684 30716 40740
rect 30772 40684 31612 40740
rect 31668 40684 31678 40740
rect 40002 40684 40012 40740
rect 40068 40684 40572 40740
rect 40628 40684 42588 40740
rect 42644 40684 42654 40740
rect 43474 40684 43484 40740
rect 43540 40684 43550 40740
rect 43652 40684 44940 40740
rect 44996 40684 45836 40740
rect 45892 40684 45902 40740
rect 43484 40628 43540 40684
rect 20178 40572 20188 40628
rect 20244 40572 20468 40628
rect 21634 40572 21644 40628
rect 21700 40572 23548 40628
rect 23604 40572 23614 40628
rect 26002 40572 26012 40628
rect 26068 40572 26908 40628
rect 29474 40572 29484 40628
rect 29540 40572 31948 40628
rect 32004 40572 32014 40628
rect 32274 40572 32284 40628
rect 32340 40572 33180 40628
rect 33236 40572 33246 40628
rect 35074 40572 35084 40628
rect 35140 40572 41356 40628
rect 41412 40572 41422 40628
rect 43484 40572 44604 40628
rect 44660 40572 44670 40628
rect 45602 40572 45612 40628
rect 45668 40572 45678 40628
rect 20412 40516 20468 40572
rect 26852 40516 26908 40572
rect 45612 40516 45668 40572
rect 15026 40460 15036 40516
rect 15092 40460 15708 40516
rect 15764 40460 15774 40516
rect 17602 40460 17612 40516
rect 17668 40460 20188 40516
rect 20244 40460 20254 40516
rect 20412 40460 23212 40516
rect 23268 40460 23278 40516
rect 26852 40460 29372 40516
rect 29428 40460 29438 40516
rect 29698 40460 29708 40516
rect 29764 40460 30492 40516
rect 30548 40460 30558 40516
rect 30706 40460 30716 40516
rect 30772 40460 30810 40516
rect 31714 40460 31724 40516
rect 31780 40460 35532 40516
rect 35588 40460 36316 40516
rect 36372 40460 36382 40516
rect 36754 40460 36764 40516
rect 36820 40460 37884 40516
rect 37940 40460 38780 40516
rect 38836 40460 40684 40516
rect 40740 40460 40750 40516
rect 43474 40460 43484 40516
rect 43540 40460 45668 40516
rect 47200 40404 48000 40432
rect 9090 40348 9100 40404
rect 9156 40348 10332 40404
rect 10388 40348 17500 40404
rect 17556 40348 20188 40404
rect 20244 40348 20254 40404
rect 27346 40348 27356 40404
rect 27412 40348 28588 40404
rect 28644 40348 28654 40404
rect 32386 40348 32396 40404
rect 32452 40348 33180 40404
rect 33236 40348 33246 40404
rect 34262 40348 34300 40404
rect 34356 40348 34366 40404
rect 36194 40348 36204 40404
rect 36260 40348 37660 40404
rect 37716 40348 38164 40404
rect 38322 40348 38332 40404
rect 38388 40348 38892 40404
rect 38948 40348 38958 40404
rect 40226 40348 40236 40404
rect 40292 40348 41020 40404
rect 41076 40348 42700 40404
rect 42756 40348 42766 40404
rect 45154 40348 45164 40404
rect 45220 40348 45724 40404
rect 45780 40348 45790 40404
rect 46844 40348 48000 40404
rect 38108 40292 38164 40348
rect 12562 40236 12572 40292
rect 12628 40236 13468 40292
rect 13524 40236 13534 40292
rect 19282 40236 19292 40292
rect 19348 40236 23548 40292
rect 23604 40236 23614 40292
rect 31378 40236 31388 40292
rect 31444 40236 31948 40292
rect 32004 40236 32014 40292
rect 36866 40236 36876 40292
rect 36932 40236 37772 40292
rect 37828 40236 37838 40292
rect 38098 40236 38108 40292
rect 38164 40236 40348 40292
rect 40404 40236 40414 40292
rect 46844 40180 46900 40348
rect 47200 40320 48000 40348
rect 17714 40124 17724 40180
rect 17780 40124 23660 40180
rect 23716 40124 23726 40180
rect 24322 40124 24332 40180
rect 24388 40124 28700 40180
rect 28756 40124 28766 40180
rect 30828 40124 35868 40180
rect 35924 40124 38332 40180
rect 38388 40124 38398 40180
rect 38994 40124 39004 40180
rect 39060 40124 41916 40180
rect 41972 40124 44156 40180
rect 44212 40124 44222 40180
rect 46834 40124 46844 40180
rect 46900 40124 46910 40180
rect 30828 40068 30884 40124
rect 28914 40012 28924 40068
rect 28980 40012 29484 40068
rect 29540 40012 30884 40068
rect 31266 40012 31276 40068
rect 31332 40012 31724 40068
rect 31780 40012 31790 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 30258 39900 30268 39956
rect 30324 39900 30828 39956
rect 30884 39900 30894 39956
rect 33926 39900 33964 39956
rect 34020 39900 34030 39956
rect 6850 39788 6860 39844
rect 6916 39788 8428 39844
rect 10098 39788 10108 39844
rect 10164 39788 11788 39844
rect 11844 39788 18956 39844
rect 19012 39788 20076 39844
rect 20132 39788 20142 39844
rect 32274 39788 32284 39844
rect 32340 39788 32564 39844
rect 43138 39788 43148 39844
rect 43204 39788 43708 39844
rect 8372 39732 8428 39788
rect 32508 39732 32564 39788
rect 43652 39732 43708 39788
rect 8372 39676 11116 39732
rect 11172 39676 11182 39732
rect 29698 39676 29708 39732
rect 29764 39676 30492 39732
rect 30548 39676 30558 39732
rect 31714 39676 31724 39732
rect 31780 39676 32508 39732
rect 32564 39676 32574 39732
rect 32946 39676 32956 39732
rect 33012 39676 33516 39732
rect 33572 39676 33582 39732
rect 43652 39676 43820 39732
rect 43876 39676 43886 39732
rect 12898 39564 12908 39620
rect 12964 39564 14140 39620
rect 14196 39564 14364 39620
rect 14420 39564 14430 39620
rect 15474 39564 15484 39620
rect 15540 39564 16940 39620
rect 16996 39564 17006 39620
rect 18722 39564 18732 39620
rect 18788 39564 20524 39620
rect 20580 39564 20590 39620
rect 29810 39564 29820 39620
rect 29876 39564 30380 39620
rect 30436 39564 30446 39620
rect 31574 39564 31612 39620
rect 31668 39564 31678 39620
rect 33058 39564 33068 39620
rect 33124 39564 35756 39620
rect 35812 39564 35822 39620
rect 36082 39564 36092 39620
rect 36148 39564 38668 39620
rect 44258 39564 44268 39620
rect 44324 39564 45052 39620
rect 45108 39564 45118 39620
rect 38612 39508 38668 39564
rect 11666 39452 11676 39508
rect 11732 39452 13468 39508
rect 13524 39452 13534 39508
rect 13794 39452 13804 39508
rect 13860 39452 14588 39508
rect 14644 39452 14654 39508
rect 15260 39452 16604 39508
rect 16660 39452 16670 39508
rect 21298 39452 21308 39508
rect 21364 39452 23212 39508
rect 23268 39452 23278 39508
rect 28914 39452 28924 39508
rect 28980 39452 32732 39508
rect 32788 39452 32798 39508
rect 33170 39452 33180 39508
rect 33236 39452 33628 39508
rect 33684 39452 33694 39508
rect 35858 39452 35868 39508
rect 35924 39452 37212 39508
rect 37268 39452 37278 39508
rect 38612 39452 38780 39508
rect 38836 39452 38846 39508
rect 39106 39452 39116 39508
rect 39172 39452 41244 39508
rect 41300 39452 41310 39508
rect 13468 39396 13524 39452
rect 15260 39396 15316 39452
rect 37212 39396 37268 39452
rect 7074 39340 7084 39396
rect 7140 39340 7756 39396
rect 7812 39340 7822 39396
rect 8372 39340 8764 39396
rect 8820 39340 8830 39396
rect 8978 39340 8988 39396
rect 9044 39340 9772 39396
rect 9828 39340 11900 39396
rect 11956 39340 11966 39396
rect 13468 39340 14028 39396
rect 14084 39340 14094 39396
rect 14466 39340 14476 39396
rect 14532 39340 15260 39396
rect 15316 39340 15326 39396
rect 16706 39340 16716 39396
rect 16772 39340 20188 39396
rect 20244 39340 20254 39396
rect 26852 39340 29148 39396
rect 29204 39340 29214 39396
rect 29670 39340 29708 39396
rect 29764 39340 29774 39396
rect 30706 39340 30716 39396
rect 30772 39340 31948 39396
rect 32004 39340 32014 39396
rect 34412 39340 35084 39396
rect 35140 39340 35150 39396
rect 37212 39340 45164 39396
rect 45220 39340 45948 39396
rect 46004 39340 46014 39396
rect 46162 39340 46172 39396
rect 46228 39340 46844 39396
rect 46900 39340 46910 39396
rect 8372 39284 8428 39340
rect 26852 39284 26908 39340
rect 6066 39228 6076 39284
rect 6132 39228 8428 39284
rect 26562 39228 26572 39284
rect 26628 39228 26908 39284
rect 27346 39228 27356 39284
rect 27412 39228 30828 39284
rect 30884 39228 30894 39284
rect 33842 39228 33852 39284
rect 33908 39228 34076 39284
rect 34132 39228 34142 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 34412 39172 34468 39340
rect 39330 39228 39340 39284
rect 39396 39228 41916 39284
rect 41972 39228 41982 39284
rect 13122 39116 13132 39172
rect 13188 39116 19292 39172
rect 19348 39116 19358 39172
rect 25106 39116 25116 39172
rect 25172 39116 27468 39172
rect 27524 39116 28028 39172
rect 28084 39116 28094 39172
rect 29138 39116 29148 39172
rect 29204 39116 29820 39172
rect 29876 39116 32172 39172
rect 32228 39116 33908 39172
rect 34178 39116 34188 39172
rect 34244 39116 34468 39172
rect 34626 39116 34636 39172
rect 34692 39116 34972 39172
rect 35028 39116 35038 39172
rect 38612 39116 43708 39172
rect 33852 39060 33908 39116
rect 38612 39060 38668 39116
rect 18274 39004 18284 39060
rect 18340 39004 20188 39060
rect 20290 39004 20300 39060
rect 20356 39004 21532 39060
rect 21588 39004 22876 39060
rect 22932 39004 22942 39060
rect 23090 39004 23100 39060
rect 23156 39004 23660 39060
rect 23716 39004 23726 39060
rect 24098 39004 24108 39060
rect 24164 39004 26348 39060
rect 26404 39004 26684 39060
rect 26740 39004 26750 39060
rect 26898 39004 26908 39060
rect 26964 39004 27002 39060
rect 27794 39004 27804 39060
rect 27860 39004 28476 39060
rect 28532 39004 28542 39060
rect 31154 39004 31164 39060
rect 31220 39004 33628 39060
rect 33684 39004 33694 39060
rect 33852 39004 38668 39060
rect 43652 39060 43708 39116
rect 43652 39004 45612 39060
rect 45668 39004 45678 39060
rect 20132 38948 20188 39004
rect 2818 38892 2828 38948
rect 2884 38892 3500 38948
rect 3556 38892 3566 38948
rect 6402 38892 6412 38948
rect 6468 38892 8988 38948
rect 9044 38892 9054 38948
rect 18050 38892 18060 38948
rect 18116 38892 19404 38948
rect 19460 38892 19470 38948
rect 20132 38892 21364 38948
rect 23314 38892 23324 38948
rect 23380 38892 27916 38948
rect 27972 38892 27982 38948
rect 28578 38892 28588 38948
rect 28644 38892 29372 38948
rect 29428 38892 29596 38948
rect 29652 38892 30268 38948
rect 30324 38892 30334 38948
rect 31714 38892 31724 38948
rect 31780 38892 42140 38948
rect 42196 38892 42206 38948
rect 21308 38836 21364 38892
rect 5058 38780 5068 38836
rect 5124 38780 8652 38836
rect 8708 38780 8718 38836
rect 15586 38780 15596 38836
rect 15652 38780 16492 38836
rect 16548 38780 16558 38836
rect 17714 38780 17724 38836
rect 17780 38780 18620 38836
rect 18676 38780 18686 38836
rect 20066 38780 20076 38836
rect 20132 38780 20860 38836
rect 20916 38780 20926 38836
rect 21298 38780 21308 38836
rect 21364 38780 21374 38836
rect 24434 38780 24444 38836
rect 24500 38780 25116 38836
rect 25172 38780 27020 38836
rect 27076 38780 27086 38836
rect 29250 38780 29260 38836
rect 29316 38780 33852 38836
rect 33908 38780 33918 38836
rect 34066 38780 34076 38836
rect 34132 38780 34412 38836
rect 34468 38780 34478 38836
rect 34626 38780 34636 38836
rect 34692 38780 34972 38836
rect 35028 38780 35038 38836
rect 38210 38780 38220 38836
rect 38276 38780 39340 38836
rect 39396 38780 40236 38836
rect 40292 38780 40302 38836
rect 45154 38780 45164 38836
rect 45220 38780 46508 38836
rect 46564 38780 46574 38836
rect 3042 38668 3052 38724
rect 3108 38668 3948 38724
rect 4004 38668 4014 38724
rect 7746 38668 7756 38724
rect 7812 38668 8428 38724
rect 9426 38668 9436 38724
rect 9492 38668 11900 38724
rect 11956 38668 11966 38724
rect 14354 38668 14364 38724
rect 14420 38668 15148 38724
rect 15204 38668 15214 38724
rect 16156 38668 18396 38724
rect 18452 38668 20412 38724
rect 20468 38668 20478 38724
rect 24322 38668 24332 38724
rect 24388 38668 25228 38724
rect 25284 38668 25294 38724
rect 26114 38668 26124 38724
rect 26180 38668 26908 38724
rect 26964 38668 26974 38724
rect 27570 38668 27580 38724
rect 27636 38668 28028 38724
rect 28084 38668 28700 38724
rect 28756 38668 28766 38724
rect 30604 38668 31724 38724
rect 31780 38668 31790 38724
rect 34290 38668 34300 38724
rect 34356 38668 35084 38724
rect 35140 38668 35150 38724
rect 8372 38612 8428 38668
rect 16156 38612 16212 38668
rect 8372 38556 9940 38612
rect 16146 38556 16156 38612
rect 16212 38556 16222 38612
rect 29138 38556 29148 38612
rect 29204 38556 29932 38612
rect 29988 38556 29998 38612
rect 9884 38500 9940 38556
rect 30604 38500 30660 38668
rect 9874 38444 9884 38500
rect 9940 38444 9950 38500
rect 17126 38444 17164 38500
rect 17220 38444 17230 38500
rect 26786 38444 26796 38500
rect 26852 38444 30604 38500
rect 30660 38444 30670 38500
rect 34598 38444 34636 38500
rect 34692 38444 34702 38500
rect 43362 38444 43372 38500
rect 43428 38444 44716 38500
rect 44772 38444 44782 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 31042 38332 31052 38388
rect 31108 38332 34972 38388
rect 35028 38332 35038 38388
rect 40786 38332 40796 38388
rect 40852 38332 45948 38388
rect 46004 38332 46014 38388
rect 3602 38220 3612 38276
rect 3668 38220 4284 38276
rect 4340 38220 4350 38276
rect 9986 38220 9996 38276
rect 10052 38220 11116 38276
rect 11172 38220 11182 38276
rect 11554 38220 11564 38276
rect 11620 38220 13132 38276
rect 13188 38220 13198 38276
rect 13356 38220 15148 38276
rect 18162 38220 18172 38276
rect 18228 38220 19404 38276
rect 19460 38220 20300 38276
rect 20356 38220 20366 38276
rect 20738 38220 20748 38276
rect 20804 38220 21756 38276
rect 21812 38220 21822 38276
rect 22530 38220 22540 38276
rect 22596 38220 23884 38276
rect 23940 38220 23950 38276
rect 26852 38220 30716 38276
rect 30772 38220 32508 38276
rect 32564 38220 34300 38276
rect 34356 38220 34366 38276
rect 38332 38220 39788 38276
rect 39844 38220 40908 38276
rect 40964 38220 40974 38276
rect 13356 38164 13412 38220
rect 15092 38164 15148 38220
rect 26852 38164 26908 38220
rect 9874 38108 9884 38164
rect 9940 38108 13412 38164
rect 13906 38108 13916 38164
rect 13972 38108 13982 38164
rect 15092 38108 26908 38164
rect 28802 38108 28812 38164
rect 28868 38108 30156 38164
rect 30212 38108 30222 38164
rect 31938 38108 31948 38164
rect 32004 38108 32732 38164
rect 32788 38108 34188 38164
rect 34244 38108 34254 38164
rect 13916 38052 13972 38108
rect 38332 38052 38388 38220
rect 38612 38108 44940 38164
rect 44996 38108 45006 38164
rect 7410 37996 7420 38052
rect 7476 37996 10108 38052
rect 10164 37996 14700 38052
rect 14756 37996 14766 38052
rect 17938 37996 17948 38052
rect 18004 37996 19068 38052
rect 19124 37996 19134 38052
rect 19618 37996 19628 38052
rect 19684 37996 21308 38052
rect 21364 37996 21374 38052
rect 22194 37996 22204 38052
rect 22260 37996 22540 38052
rect 22596 37996 22606 38052
rect 25442 37996 25452 38052
rect 25508 37996 27692 38052
rect 27748 37996 28364 38052
rect 28420 37996 28430 38052
rect 29362 37996 29372 38052
rect 29428 37996 30492 38052
rect 30548 37996 30558 38052
rect 31826 37996 31836 38052
rect 31892 37996 35980 38052
rect 36036 37996 36046 38052
rect 38322 37996 38332 38052
rect 38388 37996 38398 38052
rect 38612 37940 38668 38108
rect 41346 37996 41356 38052
rect 41412 37996 43484 38052
rect 43540 37996 45052 38052
rect 45108 37996 45118 38052
rect 3490 37884 3500 37940
rect 3556 37884 4172 37940
rect 4228 37884 4238 37940
rect 11890 37884 11900 37940
rect 11956 37884 12796 37940
rect 12852 37884 12862 37940
rect 13682 37884 13692 37940
rect 13748 37884 14252 37940
rect 14308 37884 14318 37940
rect 26786 37884 26796 37940
rect 26852 37884 27244 37940
rect 27300 37884 27310 37940
rect 28242 37884 28252 37940
rect 28308 37884 29148 37940
rect 29204 37884 29214 37940
rect 33926 37884 33964 37940
rect 34020 37884 34030 37940
rect 36418 37884 36428 37940
rect 36484 37884 38668 37940
rect 38882 37884 38892 37940
rect 38948 37884 43596 37940
rect 43652 37884 44156 37940
rect 44212 37884 44222 37940
rect 12338 37772 12348 37828
rect 12404 37772 15148 37828
rect 16706 37772 16716 37828
rect 16772 37772 17500 37828
rect 17556 37772 17566 37828
rect 28130 37772 28140 37828
rect 28196 37772 30268 37828
rect 30324 37772 30334 37828
rect 32386 37772 32396 37828
rect 32452 37772 33516 37828
rect 33572 37772 33582 37828
rect 36082 37772 36092 37828
rect 36148 37772 37212 37828
rect 37268 37772 37884 37828
rect 37940 37772 39564 37828
rect 39620 37772 39630 37828
rect 43026 37772 43036 37828
rect 43092 37772 44380 37828
rect 44436 37772 44446 37828
rect 15092 37716 15148 37772
rect 10882 37660 10892 37716
rect 10948 37660 12684 37716
rect 12740 37660 12750 37716
rect 15092 37660 17780 37716
rect 8754 37548 8764 37604
rect 8820 37548 9604 37604
rect 5170 37436 5180 37492
rect 5236 37436 8988 37492
rect 9044 37436 9054 37492
rect 9548 37380 9604 37548
rect 12684 37492 12740 37660
rect 17724 37604 17780 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 17714 37548 17724 37604
rect 17780 37548 17790 37604
rect 27682 37548 27692 37604
rect 27748 37548 28140 37604
rect 28196 37548 28206 37604
rect 33282 37548 33292 37604
rect 33348 37548 33852 37604
rect 33908 37548 33918 37604
rect 39330 37548 39340 37604
rect 39396 37548 40236 37604
rect 40292 37548 44044 37604
rect 44100 37548 44110 37604
rect 12684 37436 30940 37492
rect 30996 37436 32620 37492
rect 32676 37436 32686 37492
rect 35252 37436 36876 37492
rect 36932 37436 36942 37492
rect 38434 37436 38444 37492
rect 38500 37436 38892 37492
rect 38948 37436 39116 37492
rect 39172 37436 39182 37492
rect 39666 37436 39676 37492
rect 39732 37436 41468 37492
rect 41524 37436 43260 37492
rect 43316 37436 43326 37492
rect 8194 37324 8204 37380
rect 8260 37324 8876 37380
rect 8932 37324 8942 37380
rect 9538 37324 9548 37380
rect 9604 37324 24108 37380
rect 24164 37324 24174 37380
rect 35252 37268 35308 37436
rect 36876 37380 36932 37436
rect 36876 37324 41020 37380
rect 41076 37324 41086 37380
rect 1810 37212 1820 37268
rect 1876 37212 4620 37268
rect 4676 37212 5740 37268
rect 5796 37212 5806 37268
rect 9314 37212 9324 37268
rect 9380 37212 9884 37268
rect 9940 37212 9950 37268
rect 11778 37212 11788 37268
rect 11844 37212 12684 37268
rect 12740 37212 12750 37268
rect 16930 37212 16940 37268
rect 16996 37212 20300 37268
rect 20356 37212 20636 37268
rect 20692 37212 20702 37268
rect 24658 37212 24668 37268
rect 24724 37212 31948 37268
rect 32004 37212 32014 37268
rect 34524 37212 35308 37268
rect 1698 37100 1708 37156
rect 1764 37100 3388 37156
rect 3444 37100 3948 37156
rect 4004 37100 4014 37156
rect 12338 37100 12348 37156
rect 12404 37100 12414 37156
rect 16370 37100 16380 37156
rect 16436 37100 18508 37156
rect 18564 37100 18574 37156
rect 32386 37100 32396 37156
rect 32452 37100 33180 37156
rect 33236 37100 33246 37156
rect 4946 36988 4956 37044
rect 5012 36988 11452 37044
rect 11508 36988 11518 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 12348 36596 12404 37100
rect 34524 37044 34580 37212
rect 36866 37100 36876 37156
rect 36932 37100 39228 37156
rect 39284 37100 39294 37156
rect 43362 37100 43372 37156
rect 43428 37100 43932 37156
rect 43988 37100 43998 37156
rect 13122 36988 13132 37044
rect 13188 36988 25452 37044
rect 25508 36988 25518 37044
rect 32946 36988 32956 37044
rect 33012 36988 34524 37044
rect 34580 36988 34590 37044
rect 34962 36988 34972 37044
rect 35028 36988 39564 37044
rect 39620 36988 39630 37044
rect 42466 36988 42476 37044
rect 42532 36988 43484 37044
rect 43540 36988 43550 37044
rect 19170 36876 19180 36932
rect 19236 36876 23212 36932
rect 23268 36876 23548 36932
rect 23604 36876 23614 36932
rect 31826 36876 31836 36932
rect 31892 36876 32172 36932
rect 32228 36876 32238 36932
rect 36194 36876 36204 36932
rect 36260 36876 39676 36932
rect 39732 36876 39742 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 43698 36764 43708 36820
rect 43764 36764 44940 36820
rect 44996 36764 45006 36820
rect 44940 36708 44996 36764
rect 17014 36652 17052 36708
rect 17108 36652 17118 36708
rect 44940 36652 45556 36708
rect 12348 36540 15148 36596
rect 32498 36540 32508 36596
rect 32564 36540 33628 36596
rect 33684 36540 33852 36596
rect 33908 36540 33918 36596
rect 34822 36540 34860 36596
rect 34916 36540 34926 36596
rect 2818 36428 2828 36484
rect 2884 36428 2894 36484
rect 3266 36428 3276 36484
rect 3332 36428 3388 36484
rect 3444 36428 3454 36484
rect 2828 36372 2884 36428
rect 15092 36372 15148 36540
rect 17350 36428 17388 36484
rect 17444 36428 17454 36484
rect 17602 36428 17612 36484
rect 17668 36428 18284 36484
rect 18340 36428 18350 36484
rect 29362 36428 29372 36484
rect 29428 36428 33068 36484
rect 33124 36428 35644 36484
rect 35700 36428 35710 36484
rect 37202 36428 37212 36484
rect 37268 36428 39452 36484
rect 39508 36428 39518 36484
rect 2828 36316 3388 36372
rect 5842 36316 5852 36372
rect 5908 36316 7756 36372
rect 7812 36316 7822 36372
rect 12562 36316 12572 36372
rect 12628 36316 13468 36372
rect 13524 36316 13534 36372
rect 15092 36316 17500 36372
rect 17556 36316 17566 36372
rect 18386 36316 18396 36372
rect 18452 36316 19180 36372
rect 19236 36316 19246 36372
rect 19506 36316 19516 36372
rect 19572 36316 26348 36372
rect 26404 36316 26414 36372
rect 29586 36316 29596 36372
rect 29652 36316 29932 36372
rect 29988 36316 29998 36372
rect 30258 36316 30268 36372
rect 30324 36316 30940 36372
rect 30996 36316 31006 36372
rect 41906 36316 41916 36372
rect 41972 36316 44828 36372
rect 44884 36316 44894 36372
rect 3332 36260 3388 36316
rect 3332 36204 3836 36260
rect 3892 36204 3902 36260
rect 6962 36204 6972 36260
rect 7028 36204 8988 36260
rect 9044 36204 9054 36260
rect 14578 36204 14588 36260
rect 14644 36204 20412 36260
rect 20468 36204 20478 36260
rect 21298 36204 21308 36260
rect 21364 36204 22876 36260
rect 22932 36204 22942 36260
rect 28242 36204 28252 36260
rect 28308 36204 30156 36260
rect 30212 36204 30222 36260
rect 34626 36204 34636 36260
rect 34692 36204 38780 36260
rect 38836 36204 38846 36260
rect 44930 36204 44940 36260
rect 44996 36204 45276 36260
rect 45332 36204 45342 36260
rect 15586 36092 15596 36148
rect 15652 36092 16828 36148
rect 16884 36092 17836 36148
rect 17892 36092 17902 36148
rect 28354 36092 28364 36148
rect 28420 36092 29820 36148
rect 29876 36092 29886 36148
rect 32050 36092 32060 36148
rect 32116 36092 33516 36148
rect 33572 36092 41580 36148
rect 41636 36092 41646 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 45500 36036 45556 36652
rect 16370 35980 16380 36036
rect 16436 35980 16940 36036
rect 16996 35980 17006 36036
rect 17154 35980 17164 36036
rect 17220 35980 17258 36036
rect 17378 35980 17388 36036
rect 17444 35980 17482 36036
rect 17938 35980 17948 36036
rect 18004 35980 18014 36036
rect 23212 35980 27132 36036
rect 27188 35980 27198 36036
rect 30594 35980 30604 36036
rect 30660 35980 31388 36036
rect 31444 35980 31454 36036
rect 32610 35980 32620 36036
rect 32676 35980 33292 36036
rect 33348 35980 33358 36036
rect 35298 35980 35308 36036
rect 35364 35980 37100 36036
rect 37156 35980 40908 36036
rect 40964 35980 40974 36036
rect 45378 35980 45388 36036
rect 45444 35980 45556 36036
rect 17948 35924 18004 35980
rect 23212 35924 23268 35980
rect 17014 35868 17052 35924
rect 17108 35868 17118 35924
rect 17266 35868 17276 35924
rect 17332 35868 18004 35924
rect 23202 35868 23212 35924
rect 23268 35868 23278 35924
rect 23762 35868 23772 35924
rect 23828 35868 25228 35924
rect 25284 35868 25294 35924
rect 29250 35868 29260 35924
rect 29316 35868 30044 35924
rect 30100 35868 31276 35924
rect 31332 35868 31342 35924
rect 32172 35868 35420 35924
rect 35476 35868 35486 35924
rect 36978 35868 36988 35924
rect 37044 35868 41804 35924
rect 41860 35868 41870 35924
rect 42242 35868 42252 35924
rect 42308 35868 43036 35924
rect 43092 35868 43102 35924
rect 32172 35812 32228 35868
rect 3826 35756 3836 35812
rect 3892 35756 4732 35812
rect 4788 35756 5740 35812
rect 5796 35756 5806 35812
rect 16818 35756 16828 35812
rect 16884 35756 17948 35812
rect 18004 35756 18396 35812
rect 18452 35756 18462 35812
rect 22530 35756 22540 35812
rect 22596 35756 27244 35812
rect 27300 35756 27310 35812
rect 31126 35756 31164 35812
rect 31220 35756 32228 35812
rect 36642 35756 36652 35812
rect 36708 35756 38668 35812
rect 38724 35756 39004 35812
rect 39060 35756 39070 35812
rect 47200 35700 48000 35728
rect 5618 35644 5628 35700
rect 5684 35644 6748 35700
rect 6804 35644 9436 35700
rect 9492 35644 9502 35700
rect 15698 35644 15708 35700
rect 15764 35644 19404 35700
rect 19460 35644 19470 35700
rect 29922 35644 29932 35700
rect 29988 35644 30940 35700
rect 30996 35644 31006 35700
rect 46274 35644 46284 35700
rect 46340 35644 46620 35700
rect 46676 35644 48000 35700
rect 47200 35616 48000 35644
rect 5954 35532 5964 35588
rect 6020 35532 6860 35588
rect 6916 35532 6926 35588
rect 8866 35532 8876 35588
rect 8932 35532 9772 35588
rect 9828 35532 9838 35588
rect 12674 35532 12684 35588
rect 12740 35532 25452 35588
rect 25508 35532 25518 35588
rect 32162 35532 32172 35588
rect 32228 35532 34076 35588
rect 34132 35532 34142 35588
rect 17714 35420 17724 35476
rect 17780 35420 25676 35476
rect 25732 35420 25742 35476
rect 26450 35420 26460 35476
rect 26516 35420 29148 35476
rect 29204 35420 29214 35476
rect 32498 35420 32508 35476
rect 32564 35420 34188 35476
rect 34244 35420 35980 35476
rect 36036 35420 36046 35476
rect 39666 35420 39676 35476
rect 39732 35420 42028 35476
rect 42084 35420 42094 35476
rect 13010 35308 13020 35364
rect 13076 35308 15932 35364
rect 15988 35308 17612 35364
rect 17668 35308 17678 35364
rect 25106 35308 25116 35364
rect 25172 35308 27468 35364
rect 27524 35308 30268 35364
rect 30324 35308 30716 35364
rect 30772 35308 33068 35364
rect 33124 35308 33134 35364
rect 41010 35308 41020 35364
rect 41076 35308 42364 35364
rect 42420 35308 42430 35364
rect 45798 35308 45836 35364
rect 45892 35308 45902 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 5282 35196 5292 35252
rect 5348 35196 6524 35252
rect 6580 35196 7196 35252
rect 7252 35196 7262 35252
rect 8194 35196 8204 35252
rect 8260 35196 10108 35252
rect 10164 35196 10174 35252
rect 18050 35196 18060 35252
rect 18116 35196 20412 35252
rect 20468 35196 20478 35252
rect 21746 35196 21756 35252
rect 21812 35196 22988 35252
rect 23044 35196 23054 35252
rect 32050 35196 32060 35252
rect 32116 35196 32396 35252
rect 32452 35196 32462 35252
rect 36418 35196 36428 35252
rect 36484 35196 37772 35252
rect 37828 35196 37838 35252
rect 7858 35084 7868 35140
rect 7924 35084 8764 35140
rect 8820 35084 9884 35140
rect 9940 35084 9950 35140
rect 34850 35084 34860 35140
rect 34916 35084 34972 35140
rect 35028 35084 35038 35140
rect 37538 35084 37548 35140
rect 37604 35084 38444 35140
rect 38500 35084 38510 35140
rect 41234 35084 41244 35140
rect 41300 35084 43148 35140
rect 43204 35084 43214 35140
rect 43698 35084 43708 35140
rect 43764 35084 45836 35140
rect 45892 35084 45902 35140
rect 4834 34972 4844 35028
rect 4900 34972 6356 35028
rect 6514 34972 6524 35028
rect 6580 34972 7756 35028
rect 7812 34972 9660 35028
rect 9716 34972 9726 35028
rect 13682 34972 13692 35028
rect 13748 34972 16940 35028
rect 16996 34972 17006 35028
rect 17826 34972 17836 35028
rect 17892 34972 20524 35028
rect 20580 34972 20590 35028
rect 36306 34972 36316 35028
rect 36372 34972 37772 35028
rect 37828 34972 37838 35028
rect 43810 34972 43820 35028
rect 43876 34972 46172 35028
rect 46228 34972 46238 35028
rect 6300 34916 6356 34972
rect 2818 34860 2828 34916
rect 2884 34860 3276 34916
rect 3332 34860 4396 34916
rect 4452 34860 5068 34916
rect 5124 34860 5134 34916
rect 6290 34860 6300 34916
rect 6356 34860 7868 34916
rect 7924 34860 7934 34916
rect 16594 34860 16604 34916
rect 16660 34860 20636 34916
rect 20692 34860 21868 34916
rect 21924 34860 21934 34916
rect 35634 34860 35644 34916
rect 35700 34860 37212 34916
rect 37268 34860 37278 34916
rect 40226 34860 40236 34916
rect 40292 34860 41132 34916
rect 41188 34860 41198 34916
rect 7298 34748 7308 34804
rect 7364 34748 9996 34804
rect 10052 34748 10062 34804
rect 19954 34748 19964 34804
rect 20020 34748 21420 34804
rect 21476 34748 21486 34804
rect 35522 34748 35532 34804
rect 35588 34748 36988 34804
rect 37044 34748 37054 34804
rect 42130 34748 42140 34804
rect 42196 34748 44828 34804
rect 44884 34748 44894 34804
rect 17266 34636 17276 34692
rect 17332 34636 18508 34692
rect 18564 34636 19068 34692
rect 19124 34636 19134 34692
rect 21522 34636 21532 34692
rect 21588 34636 21868 34692
rect 21924 34636 21934 34692
rect 26898 34636 26908 34692
rect 26964 34636 27356 34692
rect 27412 34636 28588 34692
rect 28644 34636 41356 34692
rect 41412 34636 41422 34692
rect 43362 34636 43372 34692
rect 43428 34636 45052 34692
rect 45108 34636 45118 34692
rect 11890 34524 11900 34580
rect 11956 34524 12572 34580
rect 12628 34524 15148 34580
rect 20850 34524 20860 34580
rect 20916 34524 23212 34580
rect 23268 34524 23278 34580
rect 10322 34412 10332 34468
rect 10388 34412 10780 34468
rect 10836 34412 12012 34468
rect 12068 34412 12078 34468
rect 13794 34412 13804 34468
rect 13860 34412 14924 34468
rect 14980 34412 14990 34468
rect 9874 34300 9884 34356
rect 9940 34300 10444 34356
rect 10500 34300 10510 34356
rect 11106 34300 11116 34356
rect 11172 34300 11788 34356
rect 11844 34300 11854 34356
rect 13010 34300 13020 34356
rect 13076 34300 14700 34356
rect 14756 34300 14766 34356
rect 3332 34188 4396 34244
rect 4452 34188 5180 34244
rect 5236 34188 5246 34244
rect 6850 34188 6860 34244
rect 6916 34188 7812 34244
rect 9650 34188 9660 34244
rect 9716 34188 11452 34244
rect 11508 34188 11518 34244
rect 11666 34188 11676 34244
rect 11732 34188 13580 34244
rect 13636 34188 13646 34244
rect 3332 34132 3388 34188
rect 7756 34132 7812 34188
rect 2706 34076 2716 34132
rect 2772 34076 3052 34132
rect 3108 34076 3388 34132
rect 4498 34076 4508 34132
rect 4564 34076 5292 34132
rect 5348 34076 5358 34132
rect 6402 34076 6412 34132
rect 6468 34076 6972 34132
rect 7028 34076 7038 34132
rect 7746 34076 7756 34132
rect 7812 34076 8092 34132
rect 8148 34076 8158 34132
rect 11890 34076 11900 34132
rect 11956 34076 13356 34132
rect 13412 34076 13422 34132
rect 14700 34020 14756 34300
rect 15092 34244 15148 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 16482 34412 16492 34468
rect 16548 34412 19516 34468
rect 19572 34412 19582 34468
rect 25330 34412 25340 34468
rect 25396 34412 26908 34468
rect 26964 34412 27804 34468
rect 27860 34412 29148 34468
rect 29204 34412 29214 34468
rect 17042 34300 17052 34356
rect 17108 34300 17500 34356
rect 17556 34300 18956 34356
rect 19012 34300 19022 34356
rect 22642 34300 22652 34356
rect 22708 34300 23772 34356
rect 23828 34300 35644 34356
rect 35700 34300 35710 34356
rect 37202 34300 37212 34356
rect 37268 34300 39116 34356
rect 39172 34300 39182 34356
rect 43698 34300 43708 34356
rect 43764 34300 44828 34356
rect 44884 34300 46060 34356
rect 46116 34300 46126 34356
rect 15092 34188 18228 34244
rect 18610 34188 18620 34244
rect 18676 34188 20860 34244
rect 20916 34188 20926 34244
rect 23090 34188 23100 34244
rect 23156 34188 24444 34244
rect 24500 34188 25228 34244
rect 25284 34188 25294 34244
rect 32274 34188 32284 34244
rect 32340 34188 33516 34244
rect 33572 34188 34076 34244
rect 34132 34188 34142 34244
rect 34850 34188 34860 34244
rect 34916 34188 34926 34244
rect 36530 34188 36540 34244
rect 36596 34188 37324 34244
rect 37380 34188 37390 34244
rect 38210 34188 38220 34244
rect 38276 34188 39340 34244
rect 39396 34188 39406 34244
rect 41682 34188 41692 34244
rect 41748 34188 43484 34244
rect 43540 34188 43550 34244
rect 45490 34188 45500 34244
rect 45556 34188 45836 34244
rect 45892 34188 45902 34244
rect 2146 33964 2156 34020
rect 2212 33964 2940 34020
rect 2996 33964 3006 34020
rect 3378 33964 3388 34020
rect 3444 33964 4844 34020
rect 4900 33964 8204 34020
rect 8260 33964 8270 34020
rect 10994 33964 11004 34020
rect 11060 33964 11788 34020
rect 11844 33964 11854 34020
rect 12786 33964 12796 34020
rect 12852 33964 13692 34020
rect 13748 33964 13758 34020
rect 14700 33964 15260 34020
rect 15316 33964 15326 34020
rect 12002 33852 12012 33908
rect 12068 33852 13916 33908
rect 13972 33852 14476 33908
rect 14532 33852 14542 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 18172 33684 18228 34188
rect 21970 34076 21980 34132
rect 22036 34076 24108 34132
rect 24164 34076 24174 34132
rect 31826 34076 31836 34132
rect 31892 34076 32396 34132
rect 32452 34076 32844 34132
rect 32900 34076 32910 34132
rect 33618 34076 33628 34132
rect 33684 34076 34636 34132
rect 34692 34076 34702 34132
rect 34860 34020 34916 34188
rect 35858 34076 35868 34132
rect 35924 34076 37660 34132
rect 37716 34076 40460 34132
rect 40516 34076 40908 34132
rect 40964 34076 40974 34132
rect 19954 33964 19964 34020
rect 20020 33964 22316 34020
rect 22372 33964 22382 34020
rect 28354 33964 28364 34020
rect 28420 33964 29260 34020
rect 29316 33964 29326 34020
rect 34178 33964 34188 34020
rect 34244 33964 34916 34020
rect 21410 33852 21420 33908
rect 21476 33852 23100 33908
rect 23156 33852 23166 33908
rect 23874 33852 23884 33908
rect 23940 33852 25340 33908
rect 25396 33852 25406 33908
rect 25554 33852 25564 33908
rect 25620 33852 25900 33908
rect 25956 33852 25966 33908
rect 32050 33852 32060 33908
rect 32116 33852 35868 33908
rect 35924 33852 35934 33908
rect 23100 33796 23156 33852
rect 23100 33740 23996 33796
rect 24052 33740 24062 33796
rect 25638 33740 25676 33796
rect 25732 33740 25742 33796
rect 30482 33740 30492 33796
rect 30548 33740 34748 33796
rect 34804 33740 34814 33796
rect 38658 33740 38668 33796
rect 38724 33740 39788 33796
rect 39844 33740 43932 33796
rect 43988 33740 45724 33796
rect 45780 33740 45790 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 5282 33628 5292 33684
rect 5348 33628 5358 33684
rect 17042 33628 17052 33684
rect 17108 33628 17500 33684
rect 17556 33628 17566 33684
rect 18162 33628 18172 33684
rect 18228 33628 18238 33684
rect 24322 33628 24332 33684
rect 24388 33628 26124 33684
rect 26180 33628 26190 33684
rect 30594 33628 30604 33684
rect 30660 33628 31500 33684
rect 31556 33628 34412 33684
rect 34468 33628 34478 33684
rect 5292 33572 5348 33628
rect 4610 33516 4620 33572
rect 4676 33516 7532 33572
rect 7588 33516 7598 33572
rect 11778 33516 11788 33572
rect 11844 33516 16940 33572
rect 16996 33516 17006 33572
rect 19394 33516 19404 33572
rect 19460 33516 21980 33572
rect 22036 33516 23212 33572
rect 23268 33516 23278 33572
rect 28690 33516 28700 33572
rect 28756 33516 29148 33572
rect 29204 33516 29214 33572
rect 31154 33516 31164 33572
rect 31220 33516 31948 33572
rect 32004 33516 32014 33572
rect 33170 33516 33180 33572
rect 33236 33516 34300 33572
rect 34356 33516 34366 33572
rect 34850 33516 34860 33572
rect 34916 33516 35196 33572
rect 35252 33516 35262 33572
rect 42466 33516 42476 33572
rect 42532 33516 45836 33572
rect 45892 33516 45902 33572
rect 17490 33404 17500 33460
rect 17556 33404 17948 33460
rect 18004 33404 18014 33460
rect 18610 33404 18620 33460
rect 18676 33404 19628 33460
rect 19684 33404 19694 33460
rect 26002 33404 26012 33460
rect 26068 33404 28252 33460
rect 28308 33404 28318 33460
rect 30034 33404 30044 33460
rect 30100 33404 34188 33460
rect 34244 33404 34254 33460
rect 34962 33404 34972 33460
rect 35028 33404 35084 33460
rect 35140 33404 35150 33460
rect 45154 33404 45164 33460
rect 45220 33404 46172 33460
rect 46228 33404 46238 33460
rect 9986 33292 9996 33348
rect 10052 33292 11900 33348
rect 11956 33292 11966 33348
rect 28578 33292 28588 33348
rect 28644 33292 30156 33348
rect 30212 33292 30222 33348
rect 31042 33292 31052 33348
rect 31108 33292 31612 33348
rect 31668 33292 31678 33348
rect 41794 33292 41804 33348
rect 41860 33292 42252 33348
rect 42308 33292 42812 33348
rect 42868 33292 42878 33348
rect 14242 33180 14252 33236
rect 14308 33180 15372 33236
rect 15428 33180 15438 33236
rect 20402 33180 20412 33236
rect 20468 33180 22764 33236
rect 22820 33180 23436 33236
rect 23492 33180 23502 33236
rect 28130 33180 28140 33236
rect 28196 33180 29708 33236
rect 29764 33180 31164 33236
rect 31220 33180 31230 33236
rect 34290 33180 34300 33236
rect 34356 33180 36204 33236
rect 36260 33180 39788 33236
rect 39844 33180 44940 33236
rect 44996 33180 45006 33236
rect 12898 33068 12908 33124
rect 12964 33068 14028 33124
rect 14084 33068 14094 33124
rect 17462 33068 17500 33124
rect 17556 33068 17566 33124
rect 25442 33068 25452 33124
rect 25508 33068 28364 33124
rect 28420 33068 28430 33124
rect 29922 33068 29932 33124
rect 29988 33068 35084 33124
rect 35140 33068 35150 33124
rect 29932 33012 29988 33068
rect 21970 32956 21980 33012
rect 22036 32956 22876 33012
rect 22932 32956 26908 33012
rect 27234 32956 27244 33012
rect 27300 32956 29988 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 26852 32900 26908 32956
rect 26852 32844 30492 32900
rect 30548 32844 33404 32900
rect 33460 32844 33470 32900
rect 41906 32844 41916 32900
rect 41972 32844 42476 32900
rect 42532 32844 42542 32900
rect 15092 32732 16828 32788
rect 16884 32732 19740 32788
rect 19796 32732 19806 32788
rect 20850 32732 20860 32788
rect 20916 32732 21420 32788
rect 21476 32732 21486 32788
rect 26534 32732 26572 32788
rect 26628 32732 26638 32788
rect 31266 32732 31276 32788
rect 31332 32732 32396 32788
rect 32452 32732 32462 32788
rect 38882 32732 38892 32788
rect 38948 32732 41804 32788
rect 41860 32732 44156 32788
rect 44212 32732 44222 32788
rect 15092 32564 15148 32732
rect 16706 32620 16716 32676
rect 16772 32620 17388 32676
rect 17444 32620 17454 32676
rect 23324 32620 25228 32676
rect 25284 32620 26348 32676
rect 26404 32620 26414 32676
rect 29586 32620 29596 32676
rect 29652 32620 31164 32676
rect 31220 32620 31230 32676
rect 31826 32620 31836 32676
rect 31892 32620 38108 32676
rect 38164 32620 38668 32676
rect 39442 32620 39452 32676
rect 39508 32620 42028 32676
rect 42084 32620 42094 32676
rect 23324 32564 23380 32620
rect 38612 32564 38668 32620
rect 11106 32508 11116 32564
rect 11172 32508 11788 32564
rect 11844 32508 11854 32564
rect 14802 32508 14812 32564
rect 14868 32508 15148 32564
rect 16594 32508 16604 32564
rect 16660 32508 18396 32564
rect 18452 32508 19068 32564
rect 19124 32508 19516 32564
rect 19572 32508 19582 32564
rect 20738 32508 20748 32564
rect 20804 32508 22988 32564
rect 23044 32508 23054 32564
rect 23314 32508 23324 32564
rect 23380 32508 23390 32564
rect 24098 32508 24108 32564
rect 24164 32508 24556 32564
rect 24612 32508 26908 32564
rect 26964 32508 28140 32564
rect 28196 32508 28206 32564
rect 31042 32508 31052 32564
rect 31108 32508 31612 32564
rect 31668 32508 31678 32564
rect 32274 32508 32284 32564
rect 32340 32508 34524 32564
rect 34580 32508 34590 32564
rect 35970 32508 35980 32564
rect 36036 32508 38444 32564
rect 38500 32508 38510 32564
rect 38612 32508 39004 32564
rect 39060 32508 44492 32564
rect 44548 32508 44558 32564
rect 10322 32396 10332 32452
rect 10388 32396 11564 32452
rect 11620 32396 11630 32452
rect 16258 32396 16268 32452
rect 16324 32396 17948 32452
rect 18004 32396 18014 32452
rect 24434 32396 24444 32452
rect 24500 32396 26908 32452
rect 27682 32396 27692 32452
rect 27748 32396 29484 32452
rect 29540 32396 29550 32452
rect 32162 32396 32172 32452
rect 32228 32396 32620 32452
rect 32676 32396 34300 32452
rect 34356 32396 34366 32452
rect 36082 32396 36092 32452
rect 36148 32396 37996 32452
rect 38052 32396 38062 32452
rect 38220 32396 39228 32452
rect 39284 32396 39294 32452
rect 41458 32396 41468 32452
rect 41524 32396 41534 32452
rect 9538 32284 9548 32340
rect 9604 32284 10444 32340
rect 10500 32284 10510 32340
rect 20178 32284 20188 32340
rect 20244 32284 22428 32340
rect 22484 32284 22494 32340
rect 23426 32284 23436 32340
rect 23492 32284 25844 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 25788 32116 25844 32284
rect 26852 32228 26908 32396
rect 38220 32340 38276 32396
rect 41468 32340 41524 32396
rect 30146 32284 30156 32340
rect 30212 32284 30940 32340
rect 30996 32284 31006 32340
rect 37874 32284 37884 32340
rect 37940 32284 38276 32340
rect 38434 32284 38444 32340
rect 38500 32284 41524 32340
rect 42466 32284 42476 32340
rect 42532 32284 43484 32340
rect 43540 32284 43550 32340
rect 26852 32172 28364 32228
rect 28420 32172 28430 32228
rect 35858 32172 35868 32228
rect 35924 32172 42812 32228
rect 42868 32172 42878 32228
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 16370 32060 16380 32116
rect 16436 32060 16940 32116
rect 16996 32060 18060 32116
rect 18116 32060 18126 32116
rect 24434 32060 24444 32116
rect 24500 32060 25452 32116
rect 25508 32060 25518 32116
rect 25788 32060 31724 32116
rect 31780 32060 31790 32116
rect 37650 32060 37660 32116
rect 37716 32060 41020 32116
rect 41076 32060 41086 32116
rect 12226 31948 12236 32004
rect 12292 31948 15372 32004
rect 15428 31948 16268 32004
rect 16324 31948 16334 32004
rect 24546 31948 24556 32004
rect 24612 31948 26572 32004
rect 26628 31948 27468 32004
rect 27524 31948 28028 32004
rect 28084 31948 28094 32004
rect 33394 31948 33404 32004
rect 33460 31948 34076 32004
rect 34132 31948 36988 32004
rect 37044 31948 37054 32004
rect 4610 31836 4620 31892
rect 4676 31836 5740 31892
rect 5796 31836 5806 31892
rect 13906 31836 13916 31892
rect 13972 31836 14588 31892
rect 14644 31836 14654 31892
rect 19842 31836 19852 31892
rect 19908 31836 20412 31892
rect 20468 31836 21420 31892
rect 21476 31836 21486 31892
rect 24770 31836 24780 31892
rect 24836 31836 25564 31892
rect 25620 31836 25630 31892
rect 27570 31836 27580 31892
rect 27636 31836 30380 31892
rect 30436 31836 30446 31892
rect 34402 31836 34412 31892
rect 34468 31836 35756 31892
rect 35812 31836 37100 31892
rect 37156 31836 37166 31892
rect 39330 31836 39340 31892
rect 39396 31836 40460 31892
rect 40516 31836 40526 31892
rect 41570 31836 41580 31892
rect 41636 31836 42924 31892
rect 42980 31836 43820 31892
rect 43876 31836 43886 31892
rect 44930 31836 44940 31892
rect 44996 31836 45388 31892
rect 45444 31836 45454 31892
rect 7634 31724 7644 31780
rect 7700 31724 8428 31780
rect 8484 31724 15260 31780
rect 15316 31724 17276 31780
rect 17332 31724 21308 31780
rect 21364 31724 21374 31780
rect 27010 31724 27020 31780
rect 27076 31724 29036 31780
rect 29092 31724 29102 31780
rect 35522 31724 35532 31780
rect 35588 31724 37324 31780
rect 37380 31724 37390 31780
rect 41794 31724 41804 31780
rect 41860 31724 43036 31780
rect 43092 31724 45724 31780
rect 45780 31724 45790 31780
rect 7410 31612 7420 31668
rect 7476 31612 9548 31668
rect 9604 31612 9614 31668
rect 10210 31612 10220 31668
rect 10276 31612 13468 31668
rect 13524 31612 13534 31668
rect 23202 31612 23212 31668
rect 23268 31612 23660 31668
rect 23716 31612 24108 31668
rect 24164 31612 24174 31668
rect 28578 31612 28588 31668
rect 28644 31612 28654 31668
rect 37538 31612 37548 31668
rect 37604 31612 40012 31668
rect 40068 31612 40078 31668
rect 28588 31556 28644 31612
rect 5506 31500 5516 31556
rect 5572 31500 6188 31556
rect 6244 31500 6254 31556
rect 11890 31500 11900 31556
rect 11956 31500 13804 31556
rect 13860 31500 13870 31556
rect 17826 31500 17836 31556
rect 17892 31500 20412 31556
rect 20468 31500 20478 31556
rect 28588 31500 42588 31556
rect 42644 31500 42654 31556
rect 43922 31500 43932 31556
rect 43988 31500 45948 31556
rect 46004 31500 46396 31556
rect 46452 31500 46462 31556
rect 5842 31388 5852 31444
rect 5908 31388 6300 31444
rect 6356 31388 7756 31444
rect 7812 31388 7822 31444
rect 12562 31388 12572 31444
rect 12628 31388 13020 31444
rect 13076 31388 14140 31444
rect 14196 31388 14812 31444
rect 14868 31388 15484 31444
rect 15540 31388 15550 31444
rect 18610 31388 18620 31444
rect 18676 31388 19404 31444
rect 19460 31388 19470 31444
rect 28354 31388 28364 31444
rect 28420 31388 29708 31444
rect 29764 31388 29774 31444
rect 30818 31388 30828 31444
rect 30884 31388 37212 31444
rect 37268 31388 38332 31444
rect 38388 31388 38398 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 14578 31276 14588 31332
rect 14644 31276 18172 31332
rect 18228 31276 18238 31332
rect 28466 31276 28476 31332
rect 28532 31276 33852 31332
rect 33908 31276 34860 31332
rect 34916 31276 34926 31332
rect 36194 31276 36204 31332
rect 36260 31276 37660 31332
rect 37716 31276 37726 31332
rect 7186 31164 7196 31220
rect 7252 31164 8092 31220
rect 8148 31164 8158 31220
rect 35858 31164 35868 31220
rect 35924 31164 40236 31220
rect 40292 31164 40302 31220
rect 41794 31164 41804 31220
rect 41860 31164 41870 31220
rect 41804 31108 41860 31164
rect 7858 31052 7868 31108
rect 7924 31052 8428 31108
rect 8484 31052 8494 31108
rect 14690 31052 14700 31108
rect 14756 31052 15708 31108
rect 15764 31052 15774 31108
rect 19282 31052 19292 31108
rect 19348 31052 21084 31108
rect 21140 31052 23548 31108
rect 23650 31052 23660 31108
rect 23716 31052 24668 31108
rect 24724 31052 26684 31108
rect 26740 31052 26750 31108
rect 26852 31052 27916 31108
rect 27972 31052 27982 31108
rect 28802 31052 28812 31108
rect 28868 31052 41860 31108
rect 42354 31052 42364 31108
rect 42420 31052 44380 31108
rect 44436 31052 44446 31108
rect 9090 30940 9100 30996
rect 9156 30940 9884 30996
rect 9940 30940 10668 30996
rect 10724 30940 10734 30996
rect 10882 30940 10892 30996
rect 10948 30940 13356 30996
rect 13412 30940 14028 30996
rect 14084 30940 14094 30996
rect 20290 30940 20300 30996
rect 20356 30940 21756 30996
rect 21812 30940 23324 30996
rect 23380 30940 23390 30996
rect 23492 30884 23548 31052
rect 26852 30884 26908 31052
rect 47200 30996 48000 31024
rect 39554 30940 39564 30996
rect 39620 30940 41580 30996
rect 41636 30940 41646 30996
rect 46162 30940 46172 30996
rect 46228 30940 48000 30996
rect 47200 30912 48000 30940
rect 23492 30828 26908 30884
rect 30146 30828 30156 30884
rect 30212 30828 30716 30884
rect 30772 30828 31724 30884
rect 31780 30828 32508 30884
rect 32564 30828 32574 30884
rect 33954 30828 33964 30884
rect 34020 30828 34748 30884
rect 34804 30828 35980 30884
rect 36036 30828 36046 30884
rect 3332 30716 5236 30772
rect 18498 30716 18508 30772
rect 18564 30716 19404 30772
rect 19460 30716 19470 30772
rect 21410 30716 21420 30772
rect 21476 30716 23324 30772
rect 23380 30716 23390 30772
rect 26114 30716 26124 30772
rect 26180 30716 26684 30772
rect 26740 30716 31164 30772
rect 31220 30716 35084 30772
rect 35140 30716 35150 30772
rect 38322 30716 38332 30772
rect 38388 30716 40124 30772
rect 40180 30716 40190 30772
rect 3332 30324 3388 30716
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 5180 30548 5236 30716
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 5170 30492 5180 30548
rect 5236 30492 5740 30548
rect 5796 30492 5806 30548
rect 17378 30492 17388 30548
rect 17444 30492 19068 30548
rect 19124 30492 19134 30548
rect 43026 30492 43036 30548
rect 43092 30492 44268 30548
rect 44324 30492 45836 30548
rect 45892 30492 45902 30548
rect 4386 30380 4396 30436
rect 4452 30380 6972 30436
rect 7028 30380 7038 30436
rect 7298 30380 7308 30436
rect 7364 30380 8428 30436
rect 8484 30380 8494 30436
rect 3154 30268 3164 30324
rect 3220 30268 3388 30324
rect 4610 30268 4620 30324
rect 4676 30268 5628 30324
rect 5684 30268 5694 30324
rect 6738 30268 6748 30324
rect 6804 30268 7420 30324
rect 7476 30268 7868 30324
rect 7924 30268 7934 30324
rect 10322 30268 10332 30324
rect 10388 30268 10892 30324
rect 10948 30268 10958 30324
rect 18162 30268 18172 30324
rect 18228 30268 19516 30324
rect 19572 30268 19582 30324
rect 20514 30268 20524 30324
rect 20580 30268 22316 30324
rect 22372 30268 22382 30324
rect 26786 30268 26796 30324
rect 26852 30268 27244 30324
rect 27300 30268 27310 30324
rect 29250 30268 29260 30324
rect 29316 30268 30380 30324
rect 30436 30268 30446 30324
rect 3266 30156 3276 30212
rect 3332 30156 5852 30212
rect 5908 30156 5918 30212
rect 6178 30156 6188 30212
rect 6244 30156 7084 30212
rect 7140 30156 7150 30212
rect 15250 30156 15260 30212
rect 15316 30156 16380 30212
rect 16436 30156 16446 30212
rect 17602 30156 17612 30212
rect 17668 30156 19292 30212
rect 19348 30156 19628 30212
rect 19684 30156 19694 30212
rect 20402 30156 20412 30212
rect 20468 30156 21532 30212
rect 21588 30156 21598 30212
rect 22726 30156 22764 30212
rect 22820 30156 22830 30212
rect 24658 30156 24668 30212
rect 24724 30156 25340 30212
rect 25396 30156 25406 30212
rect 31378 30156 31388 30212
rect 31444 30156 33404 30212
rect 33460 30156 33470 30212
rect 35970 30156 35980 30212
rect 36036 30156 37548 30212
rect 37604 30156 37614 30212
rect 39778 30156 39788 30212
rect 39844 30156 40348 30212
rect 40404 30156 42252 30212
rect 42308 30156 44940 30212
rect 44996 30156 45388 30212
rect 45444 30156 45454 30212
rect 3826 30044 3836 30100
rect 3892 30044 5740 30100
rect 5796 30044 5806 30100
rect 8082 30044 8092 30100
rect 8148 30044 9548 30100
rect 9604 30044 9614 30100
rect 21532 29988 21588 30156
rect 33404 30100 33460 30156
rect 24882 30044 24892 30100
rect 24948 30044 25900 30100
rect 25956 30044 26348 30100
rect 26404 30044 27804 30100
rect 27860 30044 27870 30100
rect 29586 30044 29596 30100
rect 29652 30044 30268 30100
rect 30324 30044 30334 30100
rect 33404 30044 36092 30100
rect 36148 30044 36158 30100
rect 42578 30044 42588 30100
rect 42644 30044 44156 30100
rect 44212 30044 44222 30100
rect 2482 29932 2492 29988
rect 2548 29932 6636 29988
rect 6692 29932 6702 29988
rect 10658 29932 10668 29988
rect 10724 29932 12460 29988
rect 12516 29932 12526 29988
rect 17938 29932 17948 29988
rect 18004 29932 19628 29988
rect 19684 29932 20076 29988
rect 20132 29932 20142 29988
rect 21532 29932 22428 29988
rect 22484 29932 22494 29988
rect 22754 29932 22764 29988
rect 22820 29932 25676 29988
rect 25732 29932 25742 29988
rect 26852 29876 26908 29988
rect 26964 29932 26974 29988
rect 27682 29932 27692 29988
rect 27748 29932 29932 29988
rect 29988 29932 29998 29988
rect 31266 29932 31276 29988
rect 31332 29932 33404 29988
rect 33460 29932 33470 29988
rect 36418 29932 36428 29988
rect 36484 29932 39676 29988
rect 39732 29932 39742 29988
rect 21298 29820 21308 29876
rect 21364 29820 21756 29876
rect 21812 29820 21822 29876
rect 25330 29820 25340 29876
rect 25396 29820 26908 29876
rect 27570 29820 27580 29876
rect 27636 29820 29484 29876
rect 29540 29820 29550 29876
rect 30146 29820 30156 29876
rect 30212 29820 31052 29876
rect 31108 29820 32172 29876
rect 32228 29820 32238 29876
rect 32946 29820 32956 29876
rect 33012 29820 34860 29876
rect 34916 29820 37212 29876
rect 37268 29820 37278 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 1810 29708 1820 29764
rect 1876 29708 1886 29764
rect 16370 29708 16380 29764
rect 16436 29708 17836 29764
rect 17892 29708 18508 29764
rect 18564 29708 18574 29764
rect 24322 29708 24332 29764
rect 24388 29708 26460 29764
rect 26516 29708 26526 29764
rect 36092 29708 39788 29764
rect 39844 29708 39854 29764
rect 1820 29316 1876 29708
rect 6850 29596 6860 29652
rect 6916 29596 8652 29652
rect 8708 29596 8718 29652
rect 15810 29596 15820 29652
rect 15876 29596 17724 29652
rect 17780 29596 17790 29652
rect 24546 29596 24556 29652
rect 24612 29596 25228 29652
rect 25284 29596 25294 29652
rect 25442 29596 25452 29652
rect 25508 29596 30716 29652
rect 30772 29596 31276 29652
rect 31332 29596 31342 29652
rect 32274 29596 32284 29652
rect 32340 29596 33180 29652
rect 33236 29596 33246 29652
rect 33394 29596 33404 29652
rect 33460 29596 35756 29652
rect 35812 29596 35822 29652
rect 36092 29540 36148 29708
rect 40786 29596 40796 29652
rect 40852 29596 42812 29652
rect 42868 29596 45388 29652
rect 45444 29596 45454 29652
rect 3332 29484 5516 29540
rect 5572 29484 5582 29540
rect 6514 29484 6524 29540
rect 6580 29484 8876 29540
rect 8932 29484 8942 29540
rect 11218 29484 11228 29540
rect 11284 29484 11676 29540
rect 11732 29484 20636 29540
rect 20692 29484 20702 29540
rect 22866 29484 22876 29540
rect 22932 29484 30156 29540
rect 30212 29484 30222 29540
rect 30482 29484 30492 29540
rect 30548 29484 31612 29540
rect 31668 29484 34972 29540
rect 35028 29484 36092 29540
rect 36148 29484 36158 29540
rect 3332 29428 3388 29484
rect 5516 29428 5572 29484
rect 3042 29372 3052 29428
rect 3108 29372 3388 29428
rect 3714 29372 3724 29428
rect 3780 29372 4844 29428
rect 4900 29372 4910 29428
rect 5516 29372 7308 29428
rect 7364 29372 8540 29428
rect 8596 29372 8988 29428
rect 9044 29372 9054 29428
rect 22418 29372 22428 29428
rect 22484 29372 24444 29428
rect 24500 29372 27132 29428
rect 27188 29372 27198 29428
rect 32274 29372 32284 29428
rect 32340 29372 32620 29428
rect 32676 29372 32686 29428
rect 33282 29372 33292 29428
rect 33348 29372 33628 29428
rect 33684 29372 33694 29428
rect 3724 29316 3780 29372
rect 1810 29260 1820 29316
rect 1876 29260 3780 29316
rect 14466 29260 14476 29316
rect 14532 29260 15820 29316
rect 15876 29260 17164 29316
rect 17220 29260 17230 29316
rect 18946 29260 18956 29316
rect 19012 29260 21532 29316
rect 21588 29260 21598 29316
rect 23314 29260 23324 29316
rect 23380 29260 25452 29316
rect 25508 29260 25518 29316
rect 2034 29148 2044 29204
rect 2100 29148 5628 29204
rect 5684 29148 5694 29204
rect 15250 29148 15260 29204
rect 15316 29148 15484 29204
rect 15540 29148 20300 29204
rect 20356 29148 20366 29204
rect 22418 29148 22428 29204
rect 22484 29148 22876 29204
rect 22932 29148 22942 29204
rect 25554 29148 25564 29204
rect 25620 29148 29148 29204
rect 29204 29148 29214 29204
rect 18722 29036 18732 29092
rect 18788 29036 25788 29092
rect 25844 29036 25854 29092
rect 26002 29036 26012 29092
rect 26068 29036 26572 29092
rect 26628 29036 26638 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 25788 28980 25844 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 21644 28924 23996 28980
rect 24052 28924 24062 28980
rect 25788 28924 31612 28980
rect 31668 28924 31678 28980
rect 39778 28924 39788 28980
rect 39844 28924 41020 28980
rect 41076 28924 41916 28980
rect 41972 28924 42476 28980
rect 42532 28924 42542 28980
rect 21644 28868 21700 28924
rect 12226 28812 12236 28868
rect 12292 28812 20860 28868
rect 20916 28812 21644 28868
rect 21700 28812 21710 28868
rect 21970 28812 21980 28868
rect 22036 28812 23212 28868
rect 23268 28812 23278 28868
rect 25442 28812 25452 28868
rect 25508 28812 26572 28868
rect 26628 28812 26638 28868
rect 26786 28812 26796 28868
rect 26852 28812 30828 28868
rect 30884 28812 30894 28868
rect 33842 28812 33852 28868
rect 33908 28812 38444 28868
rect 38500 28812 39900 28868
rect 39956 28812 39966 28868
rect 40338 28812 40348 28868
rect 40404 28812 42364 28868
rect 42420 28812 43484 28868
rect 43540 28812 43550 28868
rect 6626 28700 6636 28756
rect 6692 28700 7420 28756
rect 7476 28700 7486 28756
rect 11106 28700 11116 28756
rect 11172 28700 11564 28756
rect 11620 28700 11630 28756
rect 13010 28700 13020 28756
rect 13076 28700 14476 28756
rect 14532 28700 14542 28756
rect 17938 28700 17948 28756
rect 18004 28700 20188 28756
rect 20244 28700 20254 28756
rect 24882 28700 24892 28756
rect 24948 28700 25340 28756
rect 25396 28700 26236 28756
rect 26292 28700 26302 28756
rect 28130 28700 28140 28756
rect 28196 28700 28308 28756
rect 28466 28700 28476 28756
rect 28532 28700 29596 28756
rect 29652 28700 32060 28756
rect 32116 28700 32126 28756
rect 33170 28700 33180 28756
rect 33236 28700 33740 28756
rect 33796 28700 34076 28756
rect 34132 28700 34142 28756
rect 41682 28700 41692 28756
rect 41748 28700 44940 28756
rect 44996 28700 45006 28756
rect 28252 28644 28308 28700
rect 8306 28588 8316 28644
rect 8372 28588 9548 28644
rect 9604 28588 9614 28644
rect 10770 28588 10780 28644
rect 10836 28588 11732 28644
rect 16930 28588 16940 28644
rect 16996 28588 19628 28644
rect 19684 28588 20748 28644
rect 20804 28588 20814 28644
rect 22614 28588 22652 28644
rect 22708 28588 22718 28644
rect 27794 28588 27804 28644
rect 27860 28588 27870 28644
rect 28252 28588 29260 28644
rect 29316 28588 29326 28644
rect 29474 28588 29484 28644
rect 29540 28588 30940 28644
rect 30996 28588 32452 28644
rect 33394 28588 33404 28644
rect 33460 28588 35980 28644
rect 36036 28588 36046 28644
rect 38434 28588 38444 28644
rect 38500 28588 39116 28644
rect 39172 28588 39182 28644
rect 39890 28588 39900 28644
rect 39956 28588 42252 28644
rect 42308 28588 42318 28644
rect 43474 28588 43484 28644
rect 43540 28588 44828 28644
rect 44884 28588 44894 28644
rect 11676 28532 11732 28588
rect 1698 28476 1708 28532
rect 1764 28476 2604 28532
rect 2660 28476 2670 28532
rect 11666 28476 11676 28532
rect 11732 28476 11742 28532
rect 21522 28476 21532 28532
rect 21588 28476 23324 28532
rect 23380 28476 23390 28532
rect 24546 28476 24556 28532
rect 24612 28476 25788 28532
rect 25844 28476 25854 28532
rect 27804 28420 27860 28588
rect 32396 28532 32452 28588
rect 32386 28476 32396 28532
rect 32452 28476 32462 28532
rect 43362 28476 43372 28532
rect 43428 28476 44156 28532
rect 44212 28476 46060 28532
rect 46116 28476 46126 28532
rect 2034 28364 2044 28420
rect 2100 28364 4956 28420
rect 5012 28364 5740 28420
rect 5796 28364 5806 28420
rect 11554 28364 11564 28420
rect 11620 28364 13468 28420
rect 13524 28364 13534 28420
rect 16930 28364 16940 28420
rect 16996 28364 18396 28420
rect 18452 28364 18462 28420
rect 19058 28364 19068 28420
rect 19124 28364 19404 28420
rect 19460 28364 20076 28420
rect 20132 28364 20142 28420
rect 26198 28364 26236 28420
rect 26292 28364 26302 28420
rect 26562 28364 26572 28420
rect 26628 28364 29148 28420
rect 29204 28364 29214 28420
rect 29922 28364 29932 28420
rect 29988 28364 32508 28420
rect 32564 28364 32574 28420
rect 37426 28364 37436 28420
rect 37492 28364 39564 28420
rect 39620 28364 40124 28420
rect 40180 28364 40572 28420
rect 40628 28364 40638 28420
rect 45826 28364 45836 28420
rect 45892 28364 46508 28420
rect 46564 28364 46574 28420
rect 10434 28252 10444 28308
rect 10500 28252 11004 28308
rect 11060 28252 11788 28308
rect 11844 28252 12124 28308
rect 12180 28252 12190 28308
rect 20178 28252 20188 28308
rect 20244 28252 33292 28308
rect 33348 28252 34188 28308
rect 34244 28252 34254 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 6402 28140 6412 28196
rect 6468 28140 7756 28196
rect 7812 28140 7822 28196
rect 8754 28140 8764 28196
rect 8820 28140 9660 28196
rect 9716 28140 11676 28196
rect 11732 28140 11742 28196
rect 28130 28140 28140 28196
rect 28196 28140 28476 28196
rect 28532 28140 28542 28196
rect 31602 28140 31612 28196
rect 31668 28140 32060 28196
rect 32116 28140 32126 28196
rect 20290 28028 20300 28084
rect 20356 28028 27244 28084
rect 27300 28028 27310 28084
rect 28140 27972 28196 28140
rect 28354 28028 28364 28084
rect 28420 28028 29260 28084
rect 29316 28028 29326 28084
rect 32274 28028 32284 28084
rect 32340 28028 32508 28084
rect 32564 28028 33516 28084
rect 33572 28028 33582 28084
rect 2818 27916 2828 27972
rect 2884 27916 3500 27972
rect 3556 27916 3566 27972
rect 5282 27916 5292 27972
rect 5348 27916 6188 27972
rect 6244 27916 6254 27972
rect 14690 27916 14700 27972
rect 14756 27916 17836 27972
rect 17892 27916 17902 27972
rect 19506 27916 19516 27972
rect 19572 27916 20188 27972
rect 20244 27916 20254 27972
rect 21746 27916 21756 27972
rect 21812 27916 22988 27972
rect 23044 27916 23054 27972
rect 26114 27916 26124 27972
rect 26180 27916 28196 27972
rect 28914 27916 28924 27972
rect 28980 27916 36092 27972
rect 36148 27916 36158 27972
rect 36978 27916 36988 27972
rect 37044 27916 38892 27972
rect 38948 27916 39284 27972
rect 39228 27860 39284 27916
rect 3938 27804 3948 27860
rect 4004 27804 5516 27860
rect 5572 27804 5582 27860
rect 5954 27804 5964 27860
rect 6020 27804 7644 27860
rect 7700 27804 7710 27860
rect 7970 27804 7980 27860
rect 8036 27804 8540 27860
rect 8596 27804 8606 27860
rect 12450 27804 12460 27860
rect 12516 27804 13580 27860
rect 13636 27804 13646 27860
rect 14018 27804 14028 27860
rect 14084 27804 15484 27860
rect 15540 27804 15550 27860
rect 32498 27804 32508 27860
rect 32564 27804 35980 27860
rect 36036 27804 36046 27860
rect 37314 27804 37324 27860
rect 37380 27804 37548 27860
rect 37604 27804 38780 27860
rect 38836 27804 38846 27860
rect 39218 27804 39228 27860
rect 39284 27804 39294 27860
rect 41206 27804 41244 27860
rect 41300 27804 42140 27860
rect 42196 27804 44828 27860
rect 44884 27804 44894 27860
rect 13346 27692 13356 27748
rect 13412 27692 14476 27748
rect 14532 27692 14542 27748
rect 17490 27692 17500 27748
rect 17556 27692 18732 27748
rect 18788 27692 18798 27748
rect 29138 27692 29148 27748
rect 29204 27692 29484 27748
rect 29540 27692 29550 27748
rect 32162 27692 32172 27748
rect 32228 27692 33068 27748
rect 33124 27692 33134 27748
rect 39778 27692 39788 27748
rect 39844 27692 41020 27748
rect 41076 27692 43260 27748
rect 43316 27692 43326 27748
rect 2594 27580 2604 27636
rect 2660 27580 3276 27636
rect 3332 27580 4732 27636
rect 4788 27580 4798 27636
rect 12114 27580 12124 27636
rect 12180 27580 14588 27636
rect 14644 27580 14654 27636
rect 16258 27580 16268 27636
rect 16324 27580 17388 27636
rect 17444 27580 17454 27636
rect 20626 27580 20636 27636
rect 20692 27580 23660 27636
rect 23716 27580 23726 27636
rect 41878 27580 41916 27636
rect 41972 27580 41982 27636
rect 20636 27524 20692 27580
rect 16818 27468 16828 27524
rect 16884 27468 20692 27524
rect 20748 27468 28700 27524
rect 28756 27468 28766 27524
rect 40786 27468 40796 27524
rect 40852 27468 42924 27524
rect 42980 27468 42990 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 20748 27412 20804 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 15922 27356 15932 27412
rect 15988 27356 20804 27412
rect 24658 27356 24668 27412
rect 24724 27356 26908 27412
rect 26964 27356 31668 27412
rect 22642 27244 22652 27300
rect 22708 27244 27580 27300
rect 27636 27244 28476 27300
rect 28532 27244 28542 27300
rect 29250 27244 29260 27300
rect 29316 27244 30380 27300
rect 30436 27244 30446 27300
rect 13234 27132 13244 27188
rect 13300 27132 13916 27188
rect 13972 27132 15036 27188
rect 15092 27132 15102 27188
rect 18274 27132 18284 27188
rect 18340 27132 24556 27188
rect 24612 27132 24622 27188
rect 31612 27076 31668 27356
rect 33282 27244 33292 27300
rect 33348 27244 33852 27300
rect 33908 27244 33918 27300
rect 34066 27244 34076 27300
rect 34132 27244 37996 27300
rect 38052 27244 38780 27300
rect 38836 27244 38846 27300
rect 43922 27244 43932 27300
rect 43988 27244 44716 27300
rect 44772 27244 44782 27300
rect 32498 27132 32508 27188
rect 32564 27132 34860 27188
rect 34916 27132 36428 27188
rect 36484 27132 36494 27188
rect 37314 27132 37324 27188
rect 37380 27132 37884 27188
rect 37940 27132 37950 27188
rect 40338 27132 40348 27188
rect 40404 27132 40414 27188
rect 41794 27132 41804 27188
rect 41860 27132 45052 27188
rect 45108 27132 45118 27188
rect 40348 27076 40404 27132
rect 13570 27020 13580 27076
rect 13636 27020 14252 27076
rect 14308 27020 14318 27076
rect 18386 27020 18396 27076
rect 18452 27020 18956 27076
rect 19012 27020 19022 27076
rect 26450 27020 26460 27076
rect 26516 27020 27692 27076
rect 27748 27020 28364 27076
rect 28420 27020 28430 27076
rect 31612 27020 35308 27076
rect 35364 27020 35374 27076
rect 40002 27020 40012 27076
rect 40068 27020 41020 27076
rect 41076 27020 41086 27076
rect 41234 27020 41244 27076
rect 41300 27020 44044 27076
rect 44100 27020 44110 27076
rect 44370 27020 44380 27076
rect 44436 27020 45612 27076
rect 45668 27020 45678 27076
rect 41244 26964 41300 27020
rect 19058 26908 19068 26964
rect 19124 26908 20412 26964
rect 20468 26908 25228 26964
rect 25284 26908 25294 26964
rect 40348 26908 41300 26964
rect 3154 26796 3164 26852
rect 3220 26796 3836 26852
rect 3892 26796 3902 26852
rect 19292 26796 19740 26852
rect 19796 26796 19806 26852
rect 20066 26796 20076 26852
rect 20132 26796 21308 26852
rect 21364 26796 21374 26852
rect 21858 26796 21868 26852
rect 21924 26796 22652 26852
rect 22708 26796 25452 26852
rect 25508 26796 25518 26852
rect 26114 26796 26124 26852
rect 26180 26796 30268 26852
rect 30324 26796 30334 26852
rect 19292 26740 19348 26796
rect 40348 26740 40404 26908
rect 40562 26796 40572 26852
rect 40628 26796 41244 26852
rect 41300 26796 41580 26852
rect 41636 26796 41646 26852
rect 43138 26796 43148 26852
rect 43204 26796 46060 26852
rect 46116 26796 46126 26852
rect 3042 26684 3052 26740
rect 3108 26684 5852 26740
rect 5908 26684 5918 26740
rect 19282 26684 19292 26740
rect 19348 26684 19358 26740
rect 26450 26684 26460 26740
rect 26516 26684 26572 26740
rect 26628 26684 26638 26740
rect 40338 26684 40348 26740
rect 40404 26684 40414 26740
rect 41458 26684 41468 26740
rect 41524 26684 46284 26740
rect 46340 26684 46350 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 2482 26572 2492 26628
rect 2548 26572 3948 26628
rect 4004 26572 4014 26628
rect 9202 26572 9212 26628
rect 9268 26572 17612 26628
rect 17668 26572 17678 26628
rect 22194 26572 22204 26628
rect 22260 26572 22988 26628
rect 23044 26572 23054 26628
rect 39554 26572 39564 26628
rect 39620 26572 41692 26628
rect 41748 26572 41758 26628
rect 41906 26572 41916 26628
rect 41972 26572 42140 26628
rect 42196 26572 42206 26628
rect 42690 26572 42700 26628
rect 42756 26572 43260 26628
rect 43316 26572 43326 26628
rect 3154 26460 3164 26516
rect 3220 26460 4620 26516
rect 4676 26460 4686 26516
rect 9650 26460 9660 26516
rect 9716 26460 10668 26516
rect 10724 26460 23212 26516
rect 23268 26460 23436 26516
rect 23492 26460 23502 26516
rect 35970 26460 35980 26516
rect 36036 26460 37884 26516
rect 37940 26460 38444 26516
rect 38500 26460 41804 26516
rect 41860 26460 45276 26516
rect 45332 26460 45342 26516
rect 22642 26348 22652 26404
rect 22708 26348 22764 26404
rect 22820 26348 26012 26404
rect 26068 26348 26078 26404
rect 26226 26348 26236 26404
rect 26292 26348 26330 26404
rect 30258 26348 30268 26404
rect 30324 26348 30828 26404
rect 30884 26348 30894 26404
rect 32386 26348 32396 26404
rect 32452 26348 32956 26404
rect 33012 26348 33022 26404
rect 47200 26292 48000 26320
rect 5730 26236 5740 26292
rect 5796 26236 9436 26292
rect 9492 26236 9502 26292
rect 10770 26236 10780 26292
rect 10836 26236 13916 26292
rect 13972 26236 13982 26292
rect 16818 26236 16828 26292
rect 16884 26236 18284 26292
rect 18340 26236 19292 26292
rect 19348 26236 19358 26292
rect 21746 26236 21756 26292
rect 21812 26236 23548 26292
rect 23604 26236 23614 26292
rect 45938 26236 45948 26292
rect 46004 26236 48000 26292
rect 47200 26208 48000 26236
rect 14690 26124 14700 26180
rect 14756 26124 20412 26180
rect 20468 26124 20478 26180
rect 36306 26124 36316 26180
rect 36372 26124 36764 26180
rect 36820 26124 36830 26180
rect 37650 26124 37660 26180
rect 37716 26124 38892 26180
rect 38948 26124 38958 26180
rect 40226 26124 40236 26180
rect 40292 26124 41468 26180
rect 41524 26124 41534 26180
rect 21410 26012 21420 26068
rect 21476 26012 22428 26068
rect 22484 26012 22494 26068
rect 31154 26012 31164 26068
rect 31220 26012 32172 26068
rect 32228 26012 32238 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 17490 25788 17500 25844
rect 17556 25788 18732 25844
rect 18788 25788 31276 25844
rect 31332 25788 31836 25844
rect 31892 25788 33180 25844
rect 33236 25788 33246 25844
rect 4498 25676 4508 25732
rect 4564 25676 5740 25732
rect 5796 25676 5806 25732
rect 18946 25676 18956 25732
rect 19012 25676 19404 25732
rect 19460 25676 25564 25732
rect 25620 25676 25630 25732
rect 34178 25676 34188 25732
rect 34244 25676 36316 25732
rect 36372 25676 36382 25732
rect 43026 25676 43036 25732
rect 43092 25676 44828 25732
rect 44884 25676 44894 25732
rect 8306 25564 8316 25620
rect 8372 25564 12796 25620
rect 12852 25564 16380 25620
rect 16436 25564 16446 25620
rect 20178 25564 20188 25620
rect 20244 25564 21196 25620
rect 21252 25564 22652 25620
rect 22708 25564 22718 25620
rect 22876 25564 28924 25620
rect 28980 25564 28990 25620
rect 30706 25564 30716 25620
rect 30772 25564 31164 25620
rect 31220 25564 31230 25620
rect 38210 25564 38220 25620
rect 38276 25564 38556 25620
rect 38612 25564 38622 25620
rect 40226 25564 40236 25620
rect 40292 25564 40796 25620
rect 40852 25564 41132 25620
rect 41188 25564 41198 25620
rect 42690 25564 42700 25620
rect 42756 25564 43372 25620
rect 43428 25564 45612 25620
rect 45668 25564 45678 25620
rect 22876 25508 22932 25564
rect 18050 25452 18060 25508
rect 18116 25452 20300 25508
rect 20356 25452 20972 25508
rect 21028 25452 22932 25508
rect 26796 25452 30996 25508
rect 31490 25452 31500 25508
rect 31556 25452 32508 25508
rect 32564 25452 32574 25508
rect 32722 25452 32732 25508
rect 32788 25452 37324 25508
rect 37380 25452 37390 25508
rect 37538 25452 37548 25508
rect 37604 25452 38780 25508
rect 38836 25452 42028 25508
rect 42084 25452 42094 25508
rect 43250 25452 43260 25508
rect 43316 25452 46060 25508
rect 46116 25452 46126 25508
rect 26796 25396 26852 25452
rect 9426 25340 9436 25396
rect 9492 25340 11004 25396
rect 11060 25340 11070 25396
rect 16482 25340 16492 25396
rect 16548 25340 21084 25396
rect 21140 25340 21150 25396
rect 24546 25340 24556 25396
rect 24612 25340 25452 25396
rect 25508 25340 26796 25396
rect 26852 25340 26862 25396
rect 30940 25284 30996 25452
rect 31154 25340 31164 25396
rect 31220 25340 31948 25396
rect 32004 25340 32014 25396
rect 36082 25340 36092 25396
rect 36148 25340 37436 25396
rect 37492 25340 37502 25396
rect 7196 25228 7756 25284
rect 7812 25228 8540 25284
rect 8596 25228 8606 25284
rect 9762 25228 9772 25284
rect 9828 25228 14252 25284
rect 14308 25228 14318 25284
rect 16818 25228 16828 25284
rect 16884 25228 18620 25284
rect 18676 25228 18686 25284
rect 23090 25228 23100 25284
rect 23156 25228 23166 25284
rect 24098 25228 24108 25284
rect 24164 25228 25340 25284
rect 25396 25228 25406 25284
rect 26114 25228 26124 25284
rect 26180 25228 29148 25284
rect 29204 25228 29214 25284
rect 30940 25228 32284 25284
rect 32340 25228 32956 25284
rect 33012 25228 33628 25284
rect 33684 25228 33694 25284
rect 35186 25228 35196 25284
rect 35252 25228 36652 25284
rect 36708 25228 36718 25284
rect 38322 25228 38332 25284
rect 38388 25228 38780 25284
rect 38836 25228 38846 25284
rect 38994 25228 39004 25284
rect 39060 25228 39508 25284
rect 39666 25228 39676 25284
rect 39732 25228 40684 25284
rect 40740 25228 40750 25284
rect 41458 25228 41468 25284
rect 41524 25228 44268 25284
rect 44324 25228 46060 25284
rect 46116 25228 46126 25284
rect 7196 25172 7252 25228
rect 23100 25172 23156 25228
rect 3154 25116 3164 25172
rect 3220 25116 3948 25172
rect 4004 25116 4014 25172
rect 7186 25116 7196 25172
rect 7252 25116 7262 25172
rect 20514 25116 20524 25172
rect 20580 25116 22316 25172
rect 22372 25116 23156 25172
rect 25666 25116 25676 25172
rect 25732 25116 37100 25172
rect 37156 25116 37166 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 39452 25060 39508 25228
rect 40898 25116 40908 25172
rect 40964 25116 44940 25172
rect 44996 25116 45006 25172
rect 6514 25004 6524 25060
rect 6580 25004 7084 25060
rect 7140 25004 7150 25060
rect 22642 25004 22652 25060
rect 22708 25004 23324 25060
rect 23380 25004 23390 25060
rect 39452 25004 39900 25060
rect 39956 25004 39966 25060
rect 41458 25004 41468 25060
rect 41524 25004 42812 25060
rect 42868 25004 43260 25060
rect 43316 25004 43326 25060
rect 1698 24892 1708 24948
rect 1764 24892 3276 24948
rect 3332 24892 4956 24948
rect 5012 24892 5404 24948
rect 5460 24892 5470 24948
rect 22530 24892 22540 24948
rect 22596 24892 23996 24948
rect 24052 24892 24062 24948
rect 27234 24892 27244 24948
rect 27300 24892 28364 24948
rect 28420 24892 28430 24948
rect 38070 24892 38108 24948
rect 38164 24892 38174 24948
rect 41122 24892 41132 24948
rect 41188 24892 43148 24948
rect 43204 24892 43214 24948
rect 6514 24780 6524 24836
rect 6580 24780 8540 24836
rect 8596 24780 8606 24836
rect 26786 24780 26796 24836
rect 26852 24780 35868 24836
rect 35924 24780 35934 24836
rect 36306 24780 36316 24836
rect 36372 24780 36764 24836
rect 36820 24780 36830 24836
rect 40114 24780 40124 24836
rect 40180 24780 41020 24836
rect 41076 24780 42364 24836
rect 42420 24780 42430 24836
rect 2370 24668 2380 24724
rect 2436 24668 3164 24724
rect 3220 24668 4620 24724
rect 4676 24668 4686 24724
rect 4946 24668 4956 24724
rect 5012 24668 6188 24724
rect 6244 24668 6254 24724
rect 8306 24668 8316 24724
rect 8372 24668 9772 24724
rect 9828 24668 9838 24724
rect 13570 24668 13580 24724
rect 13636 24668 15764 24724
rect 16370 24668 16380 24724
rect 16436 24668 17724 24724
rect 17780 24668 17790 24724
rect 34962 24668 34972 24724
rect 35028 24668 38108 24724
rect 38164 24668 38174 24724
rect 39442 24668 39452 24724
rect 39508 24668 40460 24724
rect 40516 24668 40526 24724
rect 41570 24668 41580 24724
rect 41636 24668 42252 24724
rect 42308 24668 42318 24724
rect 42466 24668 42476 24724
rect 42532 24668 43148 24724
rect 43204 24668 43214 24724
rect 15708 24612 15764 24668
rect 12674 24556 12684 24612
rect 12740 24556 14700 24612
rect 14756 24556 14766 24612
rect 15698 24556 15708 24612
rect 15764 24556 21532 24612
rect 21588 24556 22316 24612
rect 22372 24556 22382 24612
rect 31714 24556 31724 24612
rect 31780 24556 32508 24612
rect 32564 24556 34188 24612
rect 34244 24556 34254 24612
rect 38770 24556 38780 24612
rect 38836 24556 39004 24612
rect 39060 24556 40124 24612
rect 40180 24556 40908 24612
rect 40964 24556 40974 24612
rect 42914 24556 42924 24612
rect 42980 24556 44828 24612
rect 44884 24556 44894 24612
rect 3826 24444 3836 24500
rect 3892 24444 5404 24500
rect 5460 24444 5470 24500
rect 23202 24444 23212 24500
rect 23268 24444 24444 24500
rect 24500 24444 24510 24500
rect 31826 24444 31836 24500
rect 31892 24444 35868 24500
rect 35924 24444 35934 24500
rect 41682 24444 41692 24500
rect 41748 24444 46620 24500
rect 46676 24444 46686 24500
rect 6066 24332 6076 24388
rect 6132 24332 23548 24388
rect 23604 24332 23614 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 11778 24220 11788 24276
rect 11844 24220 14812 24276
rect 14868 24220 14878 24276
rect 35858 24220 35868 24276
rect 35924 24220 36204 24276
rect 36260 24220 36540 24276
rect 36596 24220 36606 24276
rect 7074 24108 7084 24164
rect 7140 24108 7756 24164
rect 7812 24108 7822 24164
rect 11442 24108 11452 24164
rect 11508 24108 12348 24164
rect 12404 24108 12414 24164
rect 25666 24108 25676 24164
rect 25732 24108 26572 24164
rect 26628 24108 29484 24164
rect 29540 24108 29550 24164
rect 29698 24108 29708 24164
rect 29764 24108 31164 24164
rect 31220 24108 31230 24164
rect 37650 24108 37660 24164
rect 37716 24108 38332 24164
rect 38388 24108 38398 24164
rect 44146 24108 44156 24164
rect 44212 24108 46060 24164
rect 46116 24108 46126 24164
rect 6626 23996 6636 24052
rect 6692 23996 8092 24052
rect 8148 23996 8652 24052
rect 8708 23996 8718 24052
rect 6066 23884 6076 23940
rect 6132 23884 7980 23940
rect 8036 23884 8046 23940
rect 12898 23884 12908 23940
rect 12964 23884 13244 23940
rect 13300 23884 13804 23940
rect 13860 23884 13870 23940
rect 21522 23884 21532 23940
rect 21588 23884 22204 23940
rect 22260 23884 22270 23940
rect 22838 23884 22876 23940
rect 22932 23884 22942 23940
rect 33954 23884 33964 23940
rect 34020 23884 34636 23940
rect 34692 23884 34702 23940
rect 36194 23884 36204 23940
rect 36260 23884 37940 23940
rect 40114 23884 40124 23940
rect 40180 23884 41132 23940
rect 41188 23884 41198 23940
rect 42354 23884 42364 23940
rect 42420 23884 42924 23940
rect 42980 23884 42990 23940
rect 43334 23884 43372 23940
rect 43428 23884 43438 23940
rect 6076 23828 6132 23884
rect 4732 23772 6132 23828
rect 7298 23772 7308 23828
rect 7364 23772 8204 23828
rect 8260 23772 8270 23828
rect 9762 23772 9772 23828
rect 9828 23772 10780 23828
rect 10836 23772 10846 23828
rect 12002 23772 12012 23828
rect 12068 23772 12460 23828
rect 12516 23772 16156 23828
rect 16212 23772 16222 23828
rect 20738 23772 20748 23828
rect 20804 23772 25340 23828
rect 25396 23772 32956 23828
rect 33012 23772 33740 23828
rect 33796 23772 33806 23828
rect 35186 23772 35196 23828
rect 35252 23772 36988 23828
rect 37044 23772 37054 23828
rect 4732 23716 4788 23772
rect 37884 23716 37940 23884
rect 40450 23772 40460 23828
rect 40516 23772 41468 23828
rect 41524 23772 41534 23828
rect 42130 23772 42140 23828
rect 42196 23772 43260 23828
rect 43316 23772 43326 23828
rect 2482 23660 2492 23716
rect 2548 23660 3612 23716
rect 3668 23660 3678 23716
rect 4722 23660 4732 23716
rect 4788 23660 4798 23716
rect 5730 23660 5740 23716
rect 5796 23660 6524 23716
rect 6580 23660 6590 23716
rect 7074 23660 7084 23716
rect 7140 23660 7980 23716
rect 8036 23660 8046 23716
rect 13570 23660 13580 23716
rect 13636 23660 14924 23716
rect 14980 23660 14990 23716
rect 17724 23660 20412 23716
rect 20468 23660 20478 23716
rect 21858 23660 21868 23716
rect 21924 23660 22988 23716
rect 23044 23660 26796 23716
rect 26852 23660 26862 23716
rect 37874 23660 37884 23716
rect 37940 23660 38108 23716
rect 38164 23660 38174 23716
rect 38434 23660 38444 23716
rect 38500 23660 41020 23716
rect 41076 23660 41086 23716
rect 41794 23660 41804 23716
rect 41860 23660 41870 23716
rect 42578 23660 42588 23716
rect 42644 23660 44044 23716
rect 44100 23660 44110 23716
rect 6402 23548 6412 23604
rect 6468 23548 8428 23604
rect 8484 23548 8494 23604
rect 14130 23548 14140 23604
rect 14196 23548 15708 23604
rect 15764 23548 15774 23604
rect 3490 23324 3500 23380
rect 3556 23324 5516 23380
rect 5572 23324 5582 23380
rect 13010 23324 13020 23380
rect 13076 23324 13692 23380
rect 13748 23324 13758 23380
rect 17724 23268 17780 23660
rect 41804 23604 41860 23660
rect 20514 23548 20524 23604
rect 20580 23548 20590 23604
rect 22082 23548 22092 23604
rect 22148 23548 23436 23604
rect 23492 23548 27580 23604
rect 27636 23548 27646 23604
rect 41804 23548 44380 23604
rect 44436 23548 45052 23604
rect 45108 23548 45118 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 20524 23380 20580 23548
rect 22502 23436 22540 23492
rect 22596 23436 22606 23492
rect 26226 23436 26236 23492
rect 26292 23436 26684 23492
rect 26740 23436 26908 23492
rect 26964 23436 26974 23492
rect 27458 23436 27468 23492
rect 27524 23436 28700 23492
rect 28756 23436 34076 23492
rect 34132 23436 34142 23492
rect 40226 23436 40236 23492
rect 40292 23436 42700 23492
rect 42756 23436 42766 23492
rect 20524 23324 22428 23380
rect 22484 23324 22988 23380
rect 23044 23324 23054 23380
rect 24546 23324 24556 23380
rect 24612 23324 25900 23380
rect 25956 23324 25966 23380
rect 26114 23324 26124 23380
rect 26180 23324 27580 23380
rect 27636 23324 27646 23380
rect 28130 23324 28140 23380
rect 28196 23324 28812 23380
rect 28868 23324 28878 23380
rect 30380 23324 33628 23380
rect 33684 23324 34188 23380
rect 34244 23324 34254 23380
rect 38322 23324 38332 23380
rect 38388 23324 38398 23380
rect 40338 23324 40348 23380
rect 40404 23324 41356 23380
rect 41412 23324 41422 23380
rect 41570 23324 41580 23380
rect 41636 23324 42252 23380
rect 42308 23324 44156 23380
rect 44212 23324 44222 23380
rect 28140 23268 28196 23324
rect 30380 23268 30436 23324
rect 38332 23268 38388 23324
rect 4610 23212 4620 23268
rect 4676 23212 5740 23268
rect 5796 23212 5806 23268
rect 6860 23212 8428 23268
rect 8484 23212 10556 23268
rect 10612 23212 10622 23268
rect 14690 23212 14700 23268
rect 14756 23212 17780 23268
rect 21298 23212 21308 23268
rect 21364 23212 23100 23268
rect 23156 23212 24220 23268
rect 24276 23212 24286 23268
rect 26002 23212 26012 23268
rect 26068 23212 28196 23268
rect 28578 23212 28588 23268
rect 28644 23212 30436 23268
rect 31686 23212 31724 23268
rect 31780 23212 31790 23268
rect 33730 23212 33740 23268
rect 33796 23212 34972 23268
rect 35028 23212 35868 23268
rect 35924 23212 36204 23268
rect 36260 23212 36270 23268
rect 37426 23212 37436 23268
rect 37492 23212 39116 23268
rect 39172 23212 39182 23268
rect 6860 23156 6916 23212
rect 4386 23100 4396 23156
rect 4452 23100 5852 23156
rect 5908 23100 5918 23156
rect 6850 23100 6860 23156
rect 6916 23100 6926 23156
rect 8194 23100 8204 23156
rect 8260 23100 8764 23156
rect 8820 23100 8830 23156
rect 9874 23100 9884 23156
rect 9940 23100 10332 23156
rect 10388 23100 10398 23156
rect 16818 23100 16828 23156
rect 16884 23100 18284 23156
rect 18340 23100 19068 23156
rect 19124 23100 19134 23156
rect 20626 23100 20636 23156
rect 20692 23100 20702 23156
rect 23650 23100 23660 23156
rect 23716 23100 25228 23156
rect 25284 23100 25564 23156
rect 25620 23100 25630 23156
rect 25778 23100 25788 23156
rect 25844 23100 27244 23156
rect 27300 23100 27310 23156
rect 28466 23100 28476 23156
rect 28532 23100 29708 23156
rect 29764 23100 29774 23156
rect 31154 23100 31164 23156
rect 31220 23100 32396 23156
rect 32452 23100 32462 23156
rect 34626 23100 34636 23156
rect 34692 23100 35756 23156
rect 35812 23100 35822 23156
rect 38546 23100 38556 23156
rect 38612 23100 39228 23156
rect 39284 23100 39294 23156
rect 42018 23100 42028 23156
rect 42084 23100 46060 23156
rect 46116 23100 46126 23156
rect 20636 23044 20692 23100
rect 16370 22988 16380 23044
rect 16436 22988 20692 23044
rect 21746 22988 21756 23044
rect 21812 22988 26572 23044
rect 26628 22988 26638 23044
rect 26908 22988 30828 23044
rect 30884 22988 30940 23044
rect 30996 22988 31006 23044
rect 31714 22988 31724 23044
rect 31780 22988 37772 23044
rect 37828 22988 37838 23044
rect 26908 22932 26964 22988
rect 5954 22876 5964 22932
rect 6020 22876 7084 22932
rect 7140 22876 7150 22932
rect 17714 22876 17724 22932
rect 17780 22876 21308 22932
rect 21364 22876 21374 22932
rect 23650 22876 23660 22932
rect 23716 22876 26964 22932
rect 28354 22876 28364 22932
rect 28420 22876 30044 22932
rect 30100 22876 30110 22932
rect 37986 22876 37996 22932
rect 38052 22876 38108 22932
rect 38164 22876 38174 22932
rect 42354 22876 42364 22932
rect 42420 22876 42924 22932
rect 42980 22876 43820 22932
rect 43876 22876 43886 22932
rect 20290 22764 20300 22820
rect 20356 22764 21532 22820
rect 21588 22764 23100 22820
rect 23156 22764 23166 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8754 22652 8764 22708
rect 8820 22652 16380 22708
rect 16436 22652 16446 22708
rect 22642 22652 22652 22708
rect 22708 22652 25788 22708
rect 25844 22652 25854 22708
rect 19730 22540 19740 22596
rect 19796 22540 20524 22596
rect 20580 22540 23884 22596
rect 23940 22540 23950 22596
rect 4722 22428 4732 22484
rect 4788 22428 7756 22484
rect 7812 22428 7822 22484
rect 12898 22428 12908 22484
rect 12964 22428 13692 22484
rect 13748 22428 13758 22484
rect 19170 22428 19180 22484
rect 19236 22428 21980 22484
rect 22036 22428 22046 22484
rect 30370 22428 30380 22484
rect 30436 22428 31836 22484
rect 31892 22428 39228 22484
rect 39284 22428 39294 22484
rect 43138 22428 43148 22484
rect 43204 22428 43708 22484
rect 43764 22428 43774 22484
rect 2818 22316 2828 22372
rect 2884 22316 4396 22372
rect 4452 22316 4462 22372
rect 9986 22316 9996 22372
rect 10052 22316 11452 22372
rect 11508 22316 11518 22372
rect 17154 22316 17164 22372
rect 17220 22316 17724 22372
rect 17780 22316 30044 22372
rect 30100 22316 30492 22372
rect 30548 22316 30558 22372
rect 42242 22316 42252 22372
rect 42308 22316 42700 22372
rect 42756 22316 42766 22372
rect 4050 22204 4060 22260
rect 4116 22204 5740 22260
rect 5796 22204 5806 22260
rect 14018 22204 14028 22260
rect 14084 22204 16268 22260
rect 16324 22204 16334 22260
rect 31378 22204 31388 22260
rect 31444 22204 33852 22260
rect 33908 22204 34524 22260
rect 34580 22204 34590 22260
rect 35634 22204 35644 22260
rect 35700 22204 37324 22260
rect 37380 22204 37390 22260
rect 41794 22204 41804 22260
rect 41860 22204 46172 22260
rect 46228 22204 46238 22260
rect 3938 22092 3948 22148
rect 4004 22092 5516 22148
rect 5572 22092 5582 22148
rect 12786 22092 12796 22148
rect 12852 22092 13804 22148
rect 13860 22092 13870 22148
rect 24322 22092 24332 22148
rect 24388 22092 25452 22148
rect 25508 22092 25518 22148
rect 35298 22092 35308 22148
rect 35364 22092 36988 22148
rect 37044 22092 37054 22148
rect 38882 22092 38892 22148
rect 38948 22092 38958 22148
rect 42242 22092 42252 22148
rect 42308 22092 45276 22148
rect 45332 22092 45342 22148
rect 30930 21980 30940 22036
rect 30996 21980 31948 22036
rect 32004 21980 32014 22036
rect 38434 21980 38444 22036
rect 38500 21980 38510 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 7074 21868 7084 21924
rect 7140 21868 8316 21924
rect 8372 21868 8382 21924
rect 14130 21868 14140 21924
rect 14196 21868 14812 21924
rect 14868 21868 14878 21924
rect 21980 21868 22652 21924
rect 22708 21868 22718 21924
rect 31276 21868 31612 21924
rect 31668 21868 31678 21924
rect 21980 21812 22036 21868
rect 31276 21812 31332 21868
rect 38444 21812 38500 21980
rect 38892 21924 38948 22092
rect 46162 21980 46172 22036
rect 46228 21980 46844 22036
rect 46900 21980 46910 22036
rect 38892 21868 45052 21924
rect 45108 21868 45118 21924
rect 5282 21756 5292 21812
rect 5348 21756 6300 21812
rect 6356 21756 6366 21812
rect 6962 21756 6972 21812
rect 7028 21756 7868 21812
rect 7924 21756 8540 21812
rect 8596 21756 8606 21812
rect 10770 21756 10780 21812
rect 10836 21756 13244 21812
rect 13300 21756 13310 21812
rect 15922 21756 15932 21812
rect 15988 21756 17948 21812
rect 18004 21756 18396 21812
rect 18452 21756 18462 21812
rect 21970 21756 21980 21812
rect 22036 21756 22046 21812
rect 22418 21756 22428 21812
rect 22484 21756 22876 21812
rect 22932 21756 22942 21812
rect 23202 21756 23212 21812
rect 23268 21756 24332 21812
rect 24388 21756 24398 21812
rect 26450 21756 26460 21812
rect 26516 21756 27244 21812
rect 27300 21756 27310 21812
rect 30370 21756 30380 21812
rect 30436 21756 31332 21812
rect 31490 21756 31500 21812
rect 31556 21756 32060 21812
rect 32116 21756 32126 21812
rect 38444 21756 39676 21812
rect 39732 21756 40236 21812
rect 40292 21756 40302 21812
rect 2706 21644 2716 21700
rect 2772 21644 4956 21700
rect 5012 21644 5852 21700
rect 5908 21644 5918 21700
rect 20962 21644 20972 21700
rect 21028 21644 22988 21700
rect 23044 21644 23054 21700
rect 24098 21644 24108 21700
rect 24164 21644 26124 21700
rect 26180 21644 26190 21700
rect 36530 21644 36540 21700
rect 36596 21644 38108 21700
rect 38164 21644 38174 21700
rect 44146 21644 44156 21700
rect 44212 21644 45388 21700
rect 45444 21644 45454 21700
rect 47200 21588 48000 21616
rect 8082 21532 8092 21588
rect 8148 21532 9772 21588
rect 9828 21532 9838 21588
rect 22866 21532 22876 21588
rect 22932 21532 23996 21588
rect 24052 21532 24062 21588
rect 25554 21532 25564 21588
rect 25620 21532 26908 21588
rect 26964 21532 26974 21588
rect 29474 21532 29484 21588
rect 29540 21532 30044 21588
rect 30100 21532 31388 21588
rect 31444 21532 31454 21588
rect 39666 21532 39676 21588
rect 39732 21532 40908 21588
rect 40964 21532 40974 21588
rect 44258 21532 44268 21588
rect 44324 21532 46060 21588
rect 46116 21532 46126 21588
rect 46274 21532 46284 21588
rect 46340 21532 48000 21588
rect 47200 21504 48000 21532
rect 2482 21420 2492 21476
rect 2548 21420 3612 21476
rect 3668 21420 3678 21476
rect 8390 21420 8428 21476
rect 8484 21420 8494 21476
rect 21298 21420 21308 21476
rect 21364 21420 23100 21476
rect 23156 21420 23166 21476
rect 23762 21420 23772 21476
rect 23828 21420 25788 21476
rect 25844 21420 25854 21476
rect 26226 21420 26236 21476
rect 26292 21420 28588 21476
rect 28644 21420 28654 21476
rect 39554 21420 39564 21476
rect 39620 21420 40348 21476
rect 40404 21420 40414 21476
rect 44146 21420 44156 21476
rect 44212 21420 44940 21476
rect 44996 21420 45006 21476
rect 18498 21308 18508 21364
rect 18564 21308 26572 21364
rect 26628 21308 29036 21364
rect 29092 21308 30604 21364
rect 30660 21308 30670 21364
rect 41570 21308 41580 21364
rect 41636 21308 42700 21364
rect 42756 21308 45164 21364
rect 45220 21308 45230 21364
rect 16706 21196 16716 21252
rect 16772 21196 21084 21252
rect 21140 21196 26348 21252
rect 26404 21196 26414 21252
rect 37874 21196 37884 21252
rect 37940 21196 39340 21252
rect 39396 21196 39406 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 38546 21084 38556 21140
rect 38612 21084 40460 21140
rect 40516 21084 42476 21140
rect 42532 21084 42542 21140
rect 12898 20972 12908 21028
rect 12964 20972 14252 21028
rect 14308 20972 15708 21028
rect 15764 20972 15774 21028
rect 35298 20972 35308 21028
rect 35364 20972 36988 21028
rect 37044 20972 44044 21028
rect 44100 20972 44940 21028
rect 44996 20972 45006 21028
rect 32162 20860 32172 20916
rect 32228 20860 33068 20916
rect 33124 20860 33134 20916
rect 33618 20860 33628 20916
rect 33684 20860 34188 20916
rect 34244 20860 39676 20916
rect 39732 20860 39742 20916
rect 40338 20860 40348 20916
rect 40404 20860 41356 20916
rect 41412 20860 42140 20916
rect 42196 20860 42206 20916
rect 12674 20748 12684 20804
rect 12740 20748 13356 20804
rect 13412 20748 14028 20804
rect 14084 20748 15372 20804
rect 15428 20748 15438 20804
rect 18162 20748 18172 20804
rect 18228 20748 19180 20804
rect 19236 20748 19246 20804
rect 19842 20748 19852 20804
rect 19908 20748 21756 20804
rect 21812 20748 21822 20804
rect 29698 20748 29708 20804
rect 29764 20748 30156 20804
rect 30212 20748 30222 20804
rect 38098 20748 38108 20804
rect 38164 20748 40908 20804
rect 40964 20748 43596 20804
rect 43652 20748 43662 20804
rect 3042 20636 3052 20692
rect 3108 20636 3500 20692
rect 3556 20636 3566 20692
rect 7746 20636 7756 20692
rect 7812 20636 9436 20692
rect 9492 20636 10668 20692
rect 10724 20636 10734 20692
rect 21186 20636 21196 20692
rect 21252 20636 24220 20692
rect 24276 20636 24286 20692
rect 27234 20636 27244 20692
rect 27300 20636 29596 20692
rect 29652 20636 29662 20692
rect 30706 20636 30716 20692
rect 30772 20636 31724 20692
rect 31780 20636 31790 20692
rect 37986 20636 37996 20692
rect 38052 20636 38668 20692
rect 38770 20636 38780 20692
rect 38836 20636 41804 20692
rect 41860 20636 41870 20692
rect 43474 20636 43484 20692
rect 43540 20636 44828 20692
rect 44884 20636 44894 20692
rect 2258 20524 2268 20580
rect 2324 20524 3948 20580
rect 4004 20524 4014 20580
rect 6290 20524 6300 20580
rect 6356 20524 6366 20580
rect 10322 20524 10332 20580
rect 10388 20524 11004 20580
rect 11060 20524 11788 20580
rect 11844 20524 11854 20580
rect 16482 20524 16492 20580
rect 16548 20524 18508 20580
rect 18564 20524 18574 20580
rect 18946 20524 18956 20580
rect 19012 20524 22764 20580
rect 22820 20524 22830 20580
rect 28242 20524 28252 20580
rect 28308 20524 28476 20580
rect 28532 20524 30044 20580
rect 30100 20524 30110 20580
rect 30258 20524 30268 20580
rect 30324 20524 30828 20580
rect 30884 20524 34972 20580
rect 35028 20524 35038 20580
rect 6300 20356 6356 20524
rect 30268 20468 30324 20524
rect 20290 20412 20300 20468
rect 20356 20412 20860 20468
rect 20916 20412 20926 20468
rect 29474 20412 29484 20468
rect 29540 20412 30324 20468
rect 38612 20468 38668 20636
rect 38612 20412 44156 20468
rect 44212 20412 44222 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 2034 20300 2044 20356
rect 2100 20300 3276 20356
rect 3332 20300 4620 20356
rect 4676 20300 4686 20356
rect 6300 20300 16716 20356
rect 16772 20300 17388 20356
rect 17444 20300 17454 20356
rect 6412 20020 6468 20300
rect 17154 20188 17164 20244
rect 17220 20188 18172 20244
rect 18228 20188 19068 20244
rect 19124 20188 19134 20244
rect 19282 20188 19292 20244
rect 19348 20188 20188 20244
rect 20244 20188 20254 20244
rect 22978 20188 22988 20244
rect 23044 20188 24332 20244
rect 24388 20188 24398 20244
rect 28242 20188 28252 20244
rect 28308 20188 28588 20244
rect 28644 20188 29372 20244
rect 29428 20188 29438 20244
rect 31686 20188 31724 20244
rect 31780 20188 31790 20244
rect 33730 20188 33740 20244
rect 33796 20188 34468 20244
rect 34412 20132 34468 20188
rect 8082 20076 8092 20132
rect 8148 20076 8876 20132
rect 8932 20076 8942 20132
rect 10098 20076 10108 20132
rect 10164 20076 15260 20132
rect 15316 20076 15326 20132
rect 17042 20076 17052 20132
rect 17108 20076 17836 20132
rect 17892 20076 18620 20132
rect 18676 20076 18956 20132
rect 19012 20076 19022 20132
rect 20514 20076 20524 20132
rect 20580 20076 22092 20132
rect 22148 20076 23436 20132
rect 23492 20076 25340 20132
rect 25396 20076 25406 20132
rect 26002 20076 26012 20132
rect 26068 20076 27356 20132
rect 27412 20076 29148 20132
rect 29204 20076 29214 20132
rect 32386 20076 32396 20132
rect 32452 20076 33068 20132
rect 33124 20076 34188 20132
rect 34244 20076 34254 20132
rect 34412 20076 36092 20132
rect 36148 20076 36158 20132
rect 38546 20076 38556 20132
rect 38612 20076 39116 20132
rect 39172 20076 39182 20132
rect 39330 20076 39340 20132
rect 39396 20076 39406 20132
rect 39340 20020 39396 20076
rect 2594 19964 2604 20020
rect 2660 19964 5516 20020
rect 5572 19964 5582 20020
rect 6290 19964 6300 20020
rect 6356 19964 6468 20020
rect 23314 19964 23324 20020
rect 23380 19964 23772 20020
rect 23828 19964 23838 20020
rect 26786 19964 26796 20020
rect 26852 19964 27580 20020
rect 27636 19964 27646 20020
rect 31826 19964 31836 20020
rect 31892 19964 33516 20020
rect 33572 19964 33740 20020
rect 33796 19964 34524 20020
rect 34580 19964 34590 20020
rect 36642 19964 36652 20020
rect 36708 19964 38220 20020
rect 38276 19964 38286 20020
rect 38770 19964 38780 20020
rect 38836 19964 39396 20020
rect 4610 19852 4620 19908
rect 4676 19852 6188 19908
rect 6244 19852 6254 19908
rect 8194 19852 8204 19908
rect 8260 19852 9772 19908
rect 9828 19852 13020 19908
rect 13076 19852 13086 19908
rect 16706 19852 16716 19908
rect 16772 19852 17948 19908
rect 18004 19852 18014 19908
rect 24546 19852 24556 19908
rect 24612 19852 27692 19908
rect 27748 19852 27758 19908
rect 30370 19852 30380 19908
rect 30436 19852 33292 19908
rect 33348 19852 33358 19908
rect 34402 19852 34412 19908
rect 34468 19852 35644 19908
rect 35700 19852 35710 19908
rect 37090 19852 37100 19908
rect 37156 19852 43372 19908
rect 43428 19852 43438 19908
rect 3042 19740 3052 19796
rect 3108 19740 4508 19796
rect 4564 19740 4574 19796
rect 5282 19740 5292 19796
rect 5348 19740 8540 19796
rect 8596 19740 8606 19796
rect 27010 19740 27020 19796
rect 27076 19740 28700 19796
rect 28756 19740 28766 19796
rect 33730 19740 33740 19796
rect 33796 19740 34524 19796
rect 34580 19740 34590 19796
rect 35186 19740 35196 19796
rect 35252 19740 35700 19796
rect 35644 19684 35700 19740
rect 35634 19628 35644 19684
rect 35700 19628 35710 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4722 19404 4732 19460
rect 4788 19404 6076 19460
rect 6132 19404 6142 19460
rect 11218 19404 11228 19460
rect 11284 19404 13580 19460
rect 13636 19404 13646 19460
rect 20066 19404 20076 19460
rect 20132 19404 20748 19460
rect 20804 19404 21532 19460
rect 21588 19404 21598 19460
rect 36194 19404 36204 19460
rect 36260 19404 37772 19460
rect 37828 19404 39172 19460
rect 40786 19404 40796 19460
rect 40852 19404 45276 19460
rect 45332 19404 45342 19460
rect 39116 19348 39172 19404
rect 2818 19292 2828 19348
rect 2884 19292 3500 19348
rect 3556 19292 4620 19348
rect 4676 19292 5740 19348
rect 5796 19292 5806 19348
rect 12002 19292 12012 19348
rect 12068 19292 13804 19348
rect 13860 19292 13870 19348
rect 18162 19292 18172 19348
rect 18228 19292 20412 19348
rect 20468 19292 20478 19348
rect 25330 19292 25340 19348
rect 25396 19292 26348 19348
rect 26404 19292 26414 19348
rect 32050 19292 32060 19348
rect 32116 19292 32844 19348
rect 32900 19292 38780 19348
rect 38836 19292 38846 19348
rect 39106 19292 39116 19348
rect 39172 19292 39676 19348
rect 39732 19292 40908 19348
rect 40964 19292 40974 19348
rect 41346 19292 41356 19348
rect 41412 19292 41804 19348
rect 41860 19292 45948 19348
rect 46004 19292 46014 19348
rect 7746 19180 7756 19236
rect 7812 19180 8652 19236
rect 8708 19180 8718 19236
rect 12226 19180 12236 19236
rect 12292 19180 14140 19236
rect 14196 19180 14206 19236
rect 34738 19180 34748 19236
rect 34804 19180 37548 19236
rect 37604 19180 39004 19236
rect 39060 19180 39564 19236
rect 39620 19180 39630 19236
rect 45154 19180 45164 19236
rect 45220 19180 45836 19236
rect 45892 19180 45902 19236
rect 2482 19068 2492 19124
rect 2548 19068 4284 19124
rect 4340 19068 4350 19124
rect 12898 19068 12908 19124
rect 12964 19068 14476 19124
rect 14532 19068 14542 19124
rect 15474 19068 15484 19124
rect 15540 19068 20412 19124
rect 20468 19068 20972 19124
rect 21028 19068 21038 19124
rect 43474 19068 43484 19124
rect 43540 19068 44828 19124
rect 44884 19068 44894 19124
rect 3826 18956 3836 19012
rect 3892 18956 5852 19012
rect 5908 18956 5918 19012
rect 7522 18956 7532 19012
rect 7588 18956 8540 19012
rect 8596 18956 9100 19012
rect 9156 18956 9166 19012
rect 20738 18956 20748 19012
rect 20804 18956 21420 19012
rect 21476 18956 21980 19012
rect 22036 18956 23100 19012
rect 23156 18956 23166 19012
rect 29250 18956 29260 19012
rect 29316 18956 29326 19012
rect 29260 18900 29316 18956
rect 5730 18844 5740 18900
rect 5796 18844 6188 18900
rect 6244 18844 6254 18900
rect 29026 18844 29036 18900
rect 29092 18844 29316 18900
rect 38322 18844 38332 18900
rect 38388 18844 39340 18900
rect 39396 18844 40236 18900
rect 40292 18844 40302 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 18834 18732 18844 18788
rect 18900 18732 19516 18788
rect 19572 18732 19582 18788
rect 19516 18676 19572 18732
rect 19516 18620 20076 18676
rect 20132 18620 20142 18676
rect 33394 18620 33404 18676
rect 33460 18620 35084 18676
rect 35140 18620 35150 18676
rect 35746 18620 35756 18676
rect 35812 18620 36652 18676
rect 36708 18620 37212 18676
rect 37268 18620 37278 18676
rect 38612 18564 38668 18676
rect 38724 18620 38734 18676
rect 39218 18620 39228 18676
rect 39284 18620 39788 18676
rect 39844 18620 40460 18676
rect 40516 18620 42588 18676
rect 42644 18620 42654 18676
rect 1810 18508 1820 18564
rect 1876 18508 3388 18564
rect 3444 18508 5292 18564
rect 5348 18508 5852 18564
rect 5908 18508 5918 18564
rect 13010 18508 13020 18564
rect 13076 18508 13524 18564
rect 16258 18508 16268 18564
rect 16324 18508 17500 18564
rect 17556 18508 17566 18564
rect 19506 18508 19516 18564
rect 19572 18508 20188 18564
rect 20244 18508 20254 18564
rect 26674 18508 26684 18564
rect 26740 18508 28252 18564
rect 28308 18508 28318 18564
rect 30034 18508 30044 18564
rect 30100 18508 30716 18564
rect 30772 18508 30782 18564
rect 33954 18508 33964 18564
rect 34020 18508 38668 18564
rect 10770 18396 10780 18452
rect 10836 18396 11900 18452
rect 11956 18396 11966 18452
rect 13468 18340 13524 18508
rect 14130 18396 14140 18452
rect 14196 18396 15372 18452
rect 15428 18396 15438 18452
rect 19282 18396 19292 18452
rect 19348 18396 19964 18452
rect 20020 18396 20030 18452
rect 20402 18396 20412 18452
rect 20468 18396 21756 18452
rect 21812 18396 22316 18452
rect 22372 18396 22382 18452
rect 23314 18396 23324 18452
rect 23380 18396 24332 18452
rect 24388 18396 24398 18452
rect 29138 18396 29148 18452
rect 29204 18396 30156 18452
rect 30212 18396 30828 18452
rect 30884 18396 30894 18452
rect 31490 18396 31500 18452
rect 31556 18396 32396 18452
rect 32452 18396 33292 18452
rect 33348 18396 33358 18452
rect 34402 18396 34412 18452
rect 34468 18396 34860 18452
rect 34916 18396 34926 18452
rect 37986 18396 37996 18452
rect 38052 18396 38444 18452
rect 38500 18396 38510 18452
rect 42690 18396 42700 18452
rect 42756 18396 43820 18452
rect 43876 18396 45164 18452
rect 45220 18396 45230 18452
rect 37996 18340 38052 18396
rect 13468 18284 15932 18340
rect 15988 18284 15998 18340
rect 21634 18284 21644 18340
rect 21700 18284 22876 18340
rect 22932 18284 22942 18340
rect 27906 18284 27916 18340
rect 27972 18284 29932 18340
rect 29988 18284 29998 18340
rect 30706 18284 30716 18340
rect 30772 18284 38052 18340
rect 44930 18284 44940 18340
rect 44996 18284 46172 18340
rect 46228 18284 46238 18340
rect 19618 18172 19628 18228
rect 19684 18172 22428 18228
rect 22484 18172 22494 18228
rect 24210 18172 24220 18228
rect 24276 18172 26012 18228
rect 26068 18172 26078 18228
rect 33702 18172 33740 18228
rect 33796 18172 33806 18228
rect 38770 18172 38780 18228
rect 38836 18172 39452 18228
rect 39508 18172 44380 18228
rect 44436 18172 45612 18228
rect 45668 18172 45678 18228
rect 14466 18060 14476 18116
rect 14532 18060 15260 18116
rect 15316 18060 17388 18116
rect 17444 18060 18284 18116
rect 18340 18060 19404 18116
rect 19460 18060 19470 18116
rect 21522 18060 21532 18116
rect 21588 18060 22988 18116
rect 23044 18060 23054 18116
rect 45378 18060 45388 18116
rect 45444 18060 46172 18116
rect 46228 18060 46238 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 22530 17948 22540 18004
rect 22596 17948 31388 18004
rect 31444 17948 31948 18004
rect 32004 17948 32014 18004
rect 31714 17836 31724 17892
rect 31780 17836 33628 17892
rect 33684 17836 37884 17892
rect 37940 17836 37950 17892
rect 15922 17724 15932 17780
rect 15988 17724 19852 17780
rect 19908 17724 20636 17780
rect 20692 17724 24668 17780
rect 24724 17724 24734 17780
rect 40786 17724 40796 17780
rect 40852 17724 44940 17780
rect 44996 17724 45006 17780
rect 45378 17724 45388 17780
rect 45444 17724 46508 17780
rect 46564 17724 46574 17780
rect 45388 17668 45444 17724
rect 12562 17612 12572 17668
rect 12628 17612 14252 17668
rect 14308 17612 15036 17668
rect 15092 17612 15102 17668
rect 31490 17612 31500 17668
rect 31556 17612 32396 17668
rect 32452 17612 34188 17668
rect 34244 17612 34254 17668
rect 41346 17612 41356 17668
rect 41412 17612 45444 17668
rect 23314 17500 23324 17556
rect 23380 17500 28588 17556
rect 28644 17500 29484 17556
rect 29540 17500 31836 17556
rect 31892 17500 34300 17556
rect 34356 17500 34366 17556
rect 37202 17500 37212 17556
rect 37268 17500 38668 17556
rect 38612 17444 38668 17500
rect 20178 17388 20188 17444
rect 20244 17388 20524 17444
rect 20580 17388 20590 17444
rect 34738 17388 34748 17444
rect 34804 17388 35196 17444
rect 35252 17388 35262 17444
rect 35634 17388 35644 17444
rect 35700 17388 37100 17444
rect 37156 17388 37166 17444
rect 38612 17388 45836 17444
rect 45892 17388 45902 17444
rect 42700 17276 43484 17332
rect 43540 17276 43550 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 42700 17220 42756 17276
rect 34962 17164 34972 17220
rect 35028 17164 36092 17220
rect 36148 17164 36158 17220
rect 36642 17164 36652 17220
rect 36708 17164 38668 17220
rect 38724 17164 41580 17220
rect 41636 17164 42700 17220
rect 42756 17164 42766 17220
rect 43362 17164 43372 17220
rect 43428 17164 44828 17220
rect 44884 17164 46060 17220
rect 46116 17164 46126 17220
rect 10098 17052 10108 17108
rect 10164 17052 10780 17108
rect 10836 17052 13244 17108
rect 13300 17052 13310 17108
rect 16034 17052 16044 17108
rect 16100 17052 20524 17108
rect 20580 17052 20590 17108
rect 24658 17052 24668 17108
rect 24724 17052 25452 17108
rect 25508 17052 25518 17108
rect 26338 17052 26348 17108
rect 26404 17052 26908 17108
rect 26964 17052 27692 17108
rect 27748 17052 31388 17108
rect 31444 17052 33068 17108
rect 33124 17052 33134 17108
rect 34066 17052 34076 17108
rect 34132 17052 37212 17108
rect 37268 17052 37278 17108
rect 38322 17052 38332 17108
rect 38388 17052 41132 17108
rect 41188 17052 42252 17108
rect 42308 17052 43036 17108
rect 43092 17052 43102 17108
rect 33068 16996 33124 17052
rect 11554 16940 11564 16996
rect 11620 16940 12796 16996
rect 12852 16940 15596 16996
rect 15652 16940 15662 16996
rect 17490 16940 17500 16996
rect 17556 16940 20412 16996
rect 20468 16940 20478 16996
rect 27570 16940 27580 16996
rect 27636 16940 28140 16996
rect 28196 16940 31724 16996
rect 31780 16940 31790 16996
rect 33068 16940 34972 16996
rect 35028 16940 35980 16996
rect 36036 16940 36046 16996
rect 38210 16940 38220 16996
rect 38276 16940 39900 16996
rect 39956 16940 39966 16996
rect 47200 16884 48000 16912
rect 9650 16828 9660 16884
rect 9716 16828 11116 16884
rect 11172 16828 11182 16884
rect 18386 16828 18396 16884
rect 18452 16828 19180 16884
rect 19236 16828 19246 16884
rect 24322 16828 24332 16884
rect 24388 16828 25452 16884
rect 25508 16828 25518 16884
rect 32274 16828 32284 16884
rect 32340 16828 32620 16884
rect 32676 16828 33516 16884
rect 33572 16828 33582 16884
rect 34626 16828 34636 16884
rect 34692 16828 36540 16884
rect 36596 16828 37436 16884
rect 37492 16828 37502 16884
rect 38546 16828 38556 16884
rect 38612 16828 40012 16884
rect 40068 16828 40078 16884
rect 46274 16828 46284 16884
rect 46340 16828 48000 16884
rect 47200 16800 48000 16828
rect 4610 16716 4620 16772
rect 4676 16716 5516 16772
rect 5572 16716 5582 16772
rect 6850 16716 6860 16772
rect 6916 16716 10556 16772
rect 10612 16716 10622 16772
rect 11218 16716 11228 16772
rect 11284 16716 12908 16772
rect 12964 16716 12974 16772
rect 14578 16716 14588 16772
rect 14644 16716 15932 16772
rect 15988 16716 15998 16772
rect 16482 16716 16492 16772
rect 16548 16716 16828 16772
rect 16884 16716 16894 16772
rect 19954 16716 19964 16772
rect 20020 16716 20748 16772
rect 20804 16716 20814 16772
rect 30258 16716 30268 16772
rect 30324 16716 31948 16772
rect 32004 16716 32014 16772
rect 35522 16716 35532 16772
rect 35588 16716 36988 16772
rect 37044 16716 37054 16772
rect 40226 16716 40236 16772
rect 40292 16716 41468 16772
rect 41524 16716 41534 16772
rect 42578 16716 42588 16772
rect 42644 16716 44828 16772
rect 44884 16716 44894 16772
rect 15026 16604 15036 16660
rect 15092 16604 16156 16660
rect 16212 16604 16222 16660
rect 20290 16604 20300 16660
rect 20356 16604 20524 16660
rect 20580 16604 20590 16660
rect 28354 16492 28364 16548
rect 28420 16492 31724 16548
rect 31780 16492 31790 16548
rect 32386 16492 32396 16548
rect 32452 16492 33404 16548
rect 33460 16492 34300 16548
rect 34356 16492 34366 16548
rect 40338 16492 40348 16548
rect 40404 16492 41468 16548
rect 41524 16492 41534 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 30044 16380 30492 16436
rect 30548 16380 30558 16436
rect 32050 16380 32060 16436
rect 32116 16380 33180 16436
rect 33236 16380 33246 16436
rect 43586 16380 43596 16436
rect 2482 16268 2492 16324
rect 2548 16268 4732 16324
rect 4788 16268 4798 16324
rect 14354 16268 14364 16324
rect 14420 16268 15596 16324
rect 15652 16268 15662 16324
rect 17938 16156 17948 16212
rect 18004 16156 18732 16212
rect 18788 16156 19404 16212
rect 19460 16156 19470 16212
rect 26114 16156 26124 16212
rect 26180 16156 26796 16212
rect 26852 16156 27692 16212
rect 27748 16156 27758 16212
rect 28578 16156 28588 16212
rect 28644 16156 29484 16212
rect 29540 16156 29550 16212
rect 8866 16044 8876 16100
rect 8932 16044 9548 16100
rect 9604 16044 11228 16100
rect 11284 16044 11294 16100
rect 17714 16044 17724 16100
rect 17780 16044 18284 16100
rect 18340 16044 18956 16100
rect 19012 16044 19022 16100
rect 23090 16044 23100 16100
rect 23156 16044 23884 16100
rect 23940 16044 23950 16100
rect 30044 15988 30100 16380
rect 38882 16268 38892 16324
rect 38948 16268 40348 16324
rect 40404 16268 40414 16324
rect 43652 16212 43708 16436
rect 32050 16156 32060 16212
rect 32116 16156 34188 16212
rect 34244 16156 34254 16212
rect 43652 16156 45276 16212
rect 45332 16156 45342 16212
rect 33170 16044 33180 16100
rect 33236 16044 36092 16100
rect 36148 16044 36158 16100
rect 41794 16044 41804 16100
rect 41860 16044 43596 16100
rect 43652 16044 43662 16100
rect 9650 15932 9660 15988
rect 9716 15932 10444 15988
rect 10500 15932 10510 15988
rect 15250 15932 15260 15988
rect 15316 15932 16380 15988
rect 16436 15932 16446 15988
rect 17826 15932 17836 15988
rect 17892 15932 20300 15988
rect 20356 15932 20366 15988
rect 27346 15932 27356 15988
rect 27412 15932 27804 15988
rect 27860 15932 27870 15988
rect 30006 15932 30044 15988
rect 30100 15932 30110 15988
rect 34962 15932 34972 15988
rect 35028 15932 35084 15988
rect 35140 15932 35150 15988
rect 42914 15932 42924 15988
rect 42980 15932 44044 15988
rect 44100 15932 44110 15988
rect 9202 15820 9212 15876
rect 9268 15820 10108 15876
rect 10164 15820 10668 15876
rect 10724 15820 10734 15876
rect 18162 15820 18172 15876
rect 18228 15820 21868 15876
rect 21924 15820 21934 15876
rect 5618 15708 5628 15764
rect 5684 15708 15036 15764
rect 15092 15708 15102 15764
rect 17602 15708 17612 15764
rect 17668 15708 18732 15764
rect 18788 15708 19180 15764
rect 19236 15708 19246 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 3490 15596 3500 15652
rect 3556 15596 3836 15652
rect 3892 15596 4732 15652
rect 4788 15596 17836 15652
rect 17892 15596 17902 15652
rect 27570 15596 27580 15652
rect 27636 15596 28476 15652
rect 28532 15596 28542 15652
rect 20514 15484 20524 15540
rect 20580 15484 22540 15540
rect 22596 15484 22606 15540
rect 27458 15484 27468 15540
rect 27524 15484 27972 15540
rect 31602 15484 31612 15540
rect 31668 15484 39788 15540
rect 39844 15484 44156 15540
rect 44212 15484 44222 15540
rect 27916 15428 27972 15484
rect 15260 15372 20860 15428
rect 20916 15372 20926 15428
rect 27906 15372 27916 15428
rect 27972 15372 27982 15428
rect 35634 15372 35644 15428
rect 35700 15372 38668 15428
rect 38724 15372 42812 15428
rect 42868 15372 42878 15428
rect 15260 15316 15316 15372
rect 6066 15260 6076 15316
rect 6132 15260 6142 15316
rect 8866 15260 8876 15316
rect 8932 15260 10332 15316
rect 10388 15260 10398 15316
rect 14914 15260 14924 15316
rect 14980 15260 15260 15316
rect 15316 15260 15326 15316
rect 18834 15260 18844 15316
rect 18900 15260 19516 15316
rect 19572 15260 19582 15316
rect 24098 15260 24108 15316
rect 24164 15260 25340 15316
rect 25396 15260 25406 15316
rect 26674 15260 26684 15316
rect 26740 15260 27636 15316
rect 28018 15260 28028 15316
rect 28084 15260 28364 15316
rect 28420 15260 28430 15316
rect 28690 15260 28700 15316
rect 28756 15260 28766 15316
rect 31266 15260 31276 15316
rect 31332 15260 31342 15316
rect 42690 15260 42700 15316
rect 42756 15260 43372 15316
rect 43428 15260 43708 15316
rect 43764 15260 43774 15316
rect 6076 15092 6132 15260
rect 8978 15148 8988 15204
rect 9044 15148 10220 15204
rect 10276 15148 10286 15204
rect 16258 15148 16268 15204
rect 16324 15148 17500 15204
rect 17556 15148 17566 15204
rect 18386 15148 18396 15204
rect 18452 15148 20300 15204
rect 20356 15148 20366 15204
rect 23762 15148 23772 15204
rect 23828 15148 25228 15204
rect 25284 15148 25294 15204
rect 25554 15148 25564 15204
rect 25620 15148 26796 15204
rect 26852 15148 26862 15204
rect 27580 15092 27636 15260
rect 28700 15092 28756 15260
rect 31276 15204 31332 15260
rect 31276 15148 32172 15204
rect 32228 15148 33628 15204
rect 33684 15148 33694 15204
rect 34738 15148 34748 15204
rect 34804 15148 34814 15204
rect 41122 15148 41132 15204
rect 41188 15148 45948 15204
rect 46004 15148 46014 15204
rect 34748 15092 34804 15148
rect 6076 15036 7084 15092
rect 7140 15036 7150 15092
rect 14130 15036 14140 15092
rect 14196 15036 23436 15092
rect 23492 15036 23502 15092
rect 26226 15036 26236 15092
rect 26292 15036 27356 15092
rect 27412 15036 27422 15092
rect 27580 15036 27692 15092
rect 27748 15036 27758 15092
rect 28354 15036 28364 15092
rect 28420 15036 28756 15092
rect 34514 15036 34524 15092
rect 34580 15036 34804 15092
rect 28578 14924 28588 14980
rect 28644 14924 29260 14980
rect 29316 14924 29820 14980
rect 29876 14924 29886 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 13122 14812 13132 14868
rect 13188 14812 15820 14868
rect 15876 14812 15886 14868
rect 8082 14700 8092 14756
rect 8148 14700 20076 14756
rect 20132 14700 20142 14756
rect 26898 14700 26908 14756
rect 26964 14700 27244 14756
rect 27300 14700 29372 14756
rect 29428 14700 29438 14756
rect 29698 14700 29708 14756
rect 29764 14700 33180 14756
rect 33236 14700 35868 14756
rect 35924 14700 36764 14756
rect 36820 14700 36830 14756
rect 7746 14588 7756 14644
rect 7812 14588 10220 14644
rect 10276 14588 10286 14644
rect 13010 14588 13020 14644
rect 13076 14588 14140 14644
rect 14196 14588 14206 14644
rect 27132 14588 27356 14644
rect 27412 14588 27422 14644
rect 30370 14588 30380 14644
rect 30436 14588 30828 14644
rect 30884 14588 30894 14644
rect 27132 14532 27188 14588
rect 4386 14476 4396 14532
rect 4452 14476 5852 14532
rect 5908 14476 5918 14532
rect 9874 14476 9884 14532
rect 9940 14476 10892 14532
rect 10948 14476 10958 14532
rect 12226 14476 12236 14532
rect 12292 14476 13692 14532
rect 13748 14476 13758 14532
rect 27122 14476 27132 14532
rect 27188 14476 27198 14532
rect 28466 14476 28476 14532
rect 28532 14476 31276 14532
rect 31332 14476 31948 14532
rect 32004 14476 32732 14532
rect 32788 14476 35868 14532
rect 35924 14476 35934 14532
rect 36194 14476 36204 14532
rect 36260 14476 37548 14532
rect 37604 14476 37614 14532
rect 40226 14476 40236 14532
rect 40292 14476 42756 14532
rect 42700 14420 42756 14476
rect 5618 14364 5628 14420
rect 5684 14364 6972 14420
rect 7028 14364 7038 14420
rect 10322 14364 10332 14420
rect 10388 14364 11788 14420
rect 11844 14364 11854 14420
rect 12450 14364 12460 14420
rect 12516 14364 13580 14420
rect 13636 14364 13646 14420
rect 20066 14364 20076 14420
rect 20132 14364 22092 14420
rect 22148 14364 22158 14420
rect 27682 14364 27692 14420
rect 27748 14364 29484 14420
rect 29540 14364 29550 14420
rect 30034 14364 30044 14420
rect 30100 14364 30380 14420
rect 30436 14364 30446 14420
rect 30902 14364 30940 14420
rect 30996 14364 31006 14420
rect 33282 14364 33292 14420
rect 33348 14364 33852 14420
rect 33908 14364 37212 14420
rect 37268 14364 37278 14420
rect 39554 14364 39564 14420
rect 39620 14364 40460 14420
rect 40516 14364 40526 14420
rect 42690 14364 42700 14420
rect 42756 14364 42766 14420
rect 42914 14364 42924 14420
rect 42980 14364 43708 14420
rect 43764 14364 43774 14420
rect 11788 14308 11844 14364
rect 7074 14252 7084 14308
rect 7140 14252 8428 14308
rect 8484 14252 8494 14308
rect 11788 14252 12572 14308
rect 12628 14252 13468 14308
rect 13524 14252 13534 14308
rect 22194 14252 22204 14308
rect 22260 14252 22540 14308
rect 22596 14252 24332 14308
rect 24388 14252 24398 14308
rect 26852 14252 29260 14308
rect 29316 14252 29326 14308
rect 36978 14252 36988 14308
rect 37044 14252 41692 14308
rect 41748 14252 41758 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 26852 14084 26908 14252
rect 33170 14140 33180 14196
rect 33236 14140 33740 14196
rect 33796 14140 33806 14196
rect 6178 14028 6188 14084
rect 6244 14028 14028 14084
rect 14084 14028 14588 14084
rect 14644 14028 14654 14084
rect 26338 14028 26348 14084
rect 26404 14028 26572 14084
rect 26628 14028 26908 14084
rect 28018 14028 28028 14084
rect 28084 14028 28700 14084
rect 28756 14028 28766 14084
rect 30258 14028 30268 14084
rect 30324 14028 30548 14084
rect 6738 13916 6748 13972
rect 6804 13916 8876 13972
rect 8932 13916 8942 13972
rect 9538 13916 9548 13972
rect 9604 13916 10444 13972
rect 10500 13916 11116 13972
rect 11172 13916 11182 13972
rect 11442 13916 11452 13972
rect 11508 13916 12124 13972
rect 12180 13916 12190 13972
rect 23538 13916 23548 13972
rect 23604 13916 30324 13972
rect 9548 13860 9604 13916
rect 30268 13860 30324 13916
rect 8754 13804 8764 13860
rect 8820 13804 9604 13860
rect 11554 13804 11564 13860
rect 11620 13804 13132 13860
rect 13188 13804 13198 13860
rect 21634 13804 21644 13860
rect 21700 13804 23660 13860
rect 23716 13804 23726 13860
rect 26786 13804 26796 13860
rect 26852 13804 28028 13860
rect 28084 13804 28094 13860
rect 30258 13804 30268 13860
rect 30324 13804 30334 13860
rect 30492 13748 30548 14028
rect 32162 13916 32172 13972
rect 32228 13916 40236 13972
rect 40292 13916 40302 13972
rect 41468 13860 41524 14252
rect 41468 13804 41916 13860
rect 41972 13804 41982 13860
rect 41468 13748 41524 13804
rect 3602 13692 3612 13748
rect 3668 13692 5180 13748
rect 5236 13692 5246 13748
rect 11106 13692 11116 13748
rect 11172 13692 14700 13748
rect 14756 13692 14766 13748
rect 19170 13692 19180 13748
rect 19236 13692 22988 13748
rect 23044 13692 23054 13748
rect 24546 13692 24556 13748
rect 24612 13692 26460 13748
rect 26516 13692 26526 13748
rect 30492 13692 31500 13748
rect 31556 13692 33292 13748
rect 33348 13692 33358 13748
rect 41458 13692 41468 13748
rect 41524 13692 41534 13748
rect 41794 13692 41804 13748
rect 41860 13692 42364 13748
rect 42420 13692 42430 13748
rect 41468 13636 41524 13692
rect 2258 13580 2268 13636
rect 2324 13580 6636 13636
rect 6692 13580 6702 13636
rect 12002 13580 12012 13636
rect 12068 13580 13804 13636
rect 13860 13580 13870 13636
rect 25778 13580 25788 13636
rect 25844 13580 26572 13636
rect 26628 13580 26638 13636
rect 31378 13580 31388 13636
rect 31444 13580 32508 13636
rect 32564 13580 35644 13636
rect 35700 13580 35710 13636
rect 41122 13580 41132 13636
rect 41188 13580 41524 13636
rect 41682 13580 41692 13636
rect 41748 13580 43036 13636
rect 43092 13580 43102 13636
rect 6738 13468 6748 13524
rect 6804 13468 7308 13524
rect 7364 13468 9772 13524
rect 9828 13468 9838 13524
rect 22082 13468 22092 13524
rect 22148 13468 22540 13524
rect 22596 13468 22606 13524
rect 24434 13468 24444 13524
rect 24500 13468 25228 13524
rect 25284 13468 26460 13524
rect 26516 13468 26526 13524
rect 27916 13468 29820 13524
rect 29876 13468 29886 13524
rect 34962 13468 34972 13524
rect 35028 13468 36092 13524
rect 36148 13468 37996 13524
rect 38052 13468 38062 13524
rect 38612 13468 42140 13524
rect 42196 13468 42206 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 27916 13300 27972 13468
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 38612 13300 38668 13468
rect 40002 13356 40012 13412
rect 40068 13356 43148 13412
rect 43204 13356 43596 13412
rect 43652 13356 43662 13412
rect 27906 13244 27916 13300
rect 27972 13244 27982 13300
rect 37874 13244 37884 13300
rect 37940 13244 38668 13300
rect 12898 13132 12908 13188
rect 12964 13132 13692 13188
rect 13748 13132 13758 13188
rect 28466 13132 28476 13188
rect 28532 13132 29708 13188
rect 29764 13132 29774 13188
rect 32834 13132 32844 13188
rect 32900 13132 45836 13188
rect 45892 13132 45902 13188
rect 3042 13020 3052 13076
rect 3108 13020 5740 13076
rect 5796 13020 5806 13076
rect 18386 13020 18396 13076
rect 18452 13020 19180 13076
rect 19236 13020 19246 13076
rect 27682 13020 27692 13076
rect 27748 13020 29148 13076
rect 29204 13020 29214 13076
rect 36418 13020 36428 13076
rect 36484 13020 37884 13076
rect 37940 13020 37950 13076
rect 42802 13020 42812 13076
rect 42868 13020 43484 13076
rect 43540 13020 43550 13076
rect 4498 12908 4508 12964
rect 4564 12908 5852 12964
rect 5908 12908 5918 12964
rect 12898 12908 12908 12964
rect 12964 12908 14252 12964
rect 14308 12908 14318 12964
rect 28018 12908 28028 12964
rect 28084 12908 28924 12964
rect 28980 12908 28990 12964
rect 32610 12908 32620 12964
rect 32676 12908 33628 12964
rect 33684 12908 33694 12964
rect 39442 12908 39452 12964
rect 39508 12908 40684 12964
rect 40740 12908 42476 12964
rect 42532 12908 42542 12964
rect 43138 12908 43148 12964
rect 43204 12908 43708 12964
rect 43764 12908 43774 12964
rect 44034 12908 44044 12964
rect 44100 12908 45276 12964
rect 45332 12908 45342 12964
rect 3266 12796 3276 12852
rect 3332 12796 3724 12852
rect 3780 12796 3790 12852
rect 18162 12796 18172 12852
rect 18228 12796 19516 12852
rect 19572 12796 19582 12852
rect 28578 12796 28588 12852
rect 28644 12796 28812 12852
rect 28868 12796 28878 12852
rect 29362 12796 29372 12852
rect 29428 12796 31836 12852
rect 31892 12796 31902 12852
rect 5058 12684 5068 12740
rect 5124 12684 6524 12740
rect 6580 12684 7532 12740
rect 7588 12684 7598 12740
rect 13794 12684 13804 12740
rect 13860 12684 15148 12740
rect 18722 12684 18732 12740
rect 18788 12684 19852 12740
rect 19908 12684 19918 12740
rect 27458 12684 27468 12740
rect 27524 12684 33180 12740
rect 33236 12684 33246 12740
rect 39750 12684 39788 12740
rect 39844 12684 39854 12740
rect 15092 12628 15148 12684
rect 4162 12572 4172 12628
rect 4228 12572 6076 12628
rect 6132 12572 6142 12628
rect 15092 12572 19628 12628
rect 19684 12572 19694 12628
rect 32386 12572 32396 12628
rect 32452 12572 33404 12628
rect 33460 12572 33470 12628
rect 19628 12404 19684 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 20178 12460 20188 12516
rect 20244 12460 21084 12516
rect 21140 12460 22428 12516
rect 22484 12460 22494 12516
rect 29586 12460 29596 12516
rect 29652 12460 30492 12516
rect 30548 12460 30558 12516
rect 31714 12460 31724 12516
rect 31780 12460 46060 12516
rect 46116 12460 46126 12516
rect 9650 12348 9660 12404
rect 9716 12348 10108 12404
rect 10164 12348 10174 12404
rect 11330 12348 11340 12404
rect 11396 12348 12236 12404
rect 12292 12348 12302 12404
rect 16146 12348 16156 12404
rect 16212 12348 16604 12404
rect 16660 12348 16670 12404
rect 17042 12348 17052 12404
rect 17108 12348 17836 12404
rect 17892 12348 17902 12404
rect 19628 12348 24108 12404
rect 24164 12348 24174 12404
rect 25554 12348 25564 12404
rect 25620 12348 27580 12404
rect 27636 12348 27646 12404
rect 29250 12348 29260 12404
rect 29316 12348 30268 12404
rect 30324 12348 30334 12404
rect 33170 12348 33180 12404
rect 33236 12348 33964 12404
rect 34020 12348 35084 12404
rect 35140 12348 37884 12404
rect 37940 12348 37950 12404
rect 44706 12348 44716 12404
rect 44772 12348 45164 12404
rect 45220 12348 45230 12404
rect 5506 12236 5516 12292
rect 5572 12236 7084 12292
rect 7140 12236 7150 12292
rect 16258 12236 16268 12292
rect 16324 12236 19292 12292
rect 19348 12236 19358 12292
rect 22866 12236 22876 12292
rect 22932 12236 23996 12292
rect 24052 12236 24062 12292
rect 26450 12236 26460 12292
rect 26516 12236 27244 12292
rect 27300 12236 27310 12292
rect 29138 12236 29148 12292
rect 29204 12236 30156 12292
rect 30212 12236 30222 12292
rect 36642 12236 36652 12292
rect 36708 12236 37548 12292
rect 37604 12236 37614 12292
rect 46060 12180 46116 12460
rect 47200 12180 48000 12208
rect 5730 12124 5740 12180
rect 5796 12124 5964 12180
rect 6020 12124 6636 12180
rect 6692 12124 6702 12180
rect 19170 12124 19180 12180
rect 19236 12124 20076 12180
rect 20132 12124 20142 12180
rect 23874 12124 23884 12180
rect 23940 12124 25788 12180
rect 25844 12124 26908 12180
rect 26964 12124 26974 12180
rect 28018 12124 28028 12180
rect 28084 12124 30828 12180
rect 30884 12124 30894 12180
rect 32498 12124 32508 12180
rect 32564 12124 33180 12180
rect 33236 12124 33246 12180
rect 33730 12124 33740 12180
rect 33796 12124 35868 12180
rect 35924 12124 36428 12180
rect 36484 12124 36494 12180
rect 43474 12124 43484 12180
rect 43540 12124 44492 12180
rect 44548 12124 44558 12180
rect 46060 12124 48000 12180
rect 47200 12096 48000 12124
rect 23650 12012 23660 12068
rect 23716 12012 26124 12068
rect 26180 12012 26190 12068
rect 28466 12012 28476 12068
rect 28532 12012 29260 12068
rect 29316 12012 29326 12068
rect 32162 12012 32172 12068
rect 32228 12012 34300 12068
rect 34356 12012 34366 12068
rect 35186 12012 35196 12068
rect 35252 12012 35980 12068
rect 36036 12012 36652 12068
rect 36708 12012 36718 12068
rect 24434 11900 24444 11956
rect 24500 11900 26684 11956
rect 26740 11900 27132 11956
rect 27188 11900 27198 11956
rect 28690 11900 28700 11956
rect 28756 11900 31052 11956
rect 31108 11900 31118 11956
rect 36194 11900 36204 11956
rect 36260 11900 36876 11956
rect 36932 11900 36942 11956
rect 6178 11788 6188 11844
rect 6244 11788 6748 11844
rect 6804 11788 6814 11844
rect 18386 11788 18396 11844
rect 18452 11788 20300 11844
rect 20356 11788 21196 11844
rect 21252 11788 21262 11844
rect 21858 11788 21868 11844
rect 21924 11788 22876 11844
rect 22932 11788 28812 11844
rect 28868 11788 28878 11844
rect 29362 11788 29372 11844
rect 29428 11788 32620 11844
rect 32676 11788 32686 11844
rect 36988 11788 37324 11844
rect 37380 11788 37660 11844
rect 37716 11788 37726 11844
rect 41570 11788 41580 11844
rect 41636 11788 41646 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 15810 11732 15820 11788
rect 15876 11732 15886 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 36988 11732 37044 11788
rect 41580 11732 41636 11788
rect 15586 11676 15596 11732
rect 15652 11676 15876 11732
rect 35970 11676 35980 11732
rect 36036 11676 37044 11732
rect 37202 11676 37212 11732
rect 37268 11676 37940 11732
rect 38210 11676 38220 11732
rect 38276 11676 39228 11732
rect 39284 11676 39294 11732
rect 41234 11676 41244 11732
rect 41300 11676 41636 11732
rect 41906 11676 41916 11732
rect 41972 11676 43820 11732
rect 43876 11676 43886 11732
rect 15474 11564 15484 11620
rect 15540 11564 15820 11620
rect 15876 11564 15886 11620
rect 28578 11564 28588 11620
rect 28644 11564 30604 11620
rect 30660 11564 30670 11620
rect 37426 11564 37436 11620
rect 37492 11564 37502 11620
rect 37622 11564 37660 11620
rect 37716 11564 37726 11620
rect 18386 11452 18396 11508
rect 18452 11452 20188 11508
rect 20244 11452 20254 11508
rect 37436 11396 37492 11564
rect 37884 11508 37940 11676
rect 41580 11620 41636 11676
rect 39106 11564 39116 11620
rect 39172 11564 43372 11620
rect 43428 11564 43438 11620
rect 37884 11452 39732 11508
rect 40114 11452 40124 11508
rect 40180 11452 41356 11508
rect 41412 11452 41422 11508
rect 39676 11396 39732 11452
rect 4834 11340 4844 11396
rect 4900 11340 5964 11396
rect 6020 11340 6030 11396
rect 15474 11340 15484 11396
rect 15540 11340 15932 11396
rect 15988 11340 15998 11396
rect 21746 11340 21756 11396
rect 21812 11340 23548 11396
rect 23604 11340 23614 11396
rect 34402 11340 34412 11396
rect 34468 11340 37436 11396
rect 37492 11340 37502 11396
rect 37650 11340 37660 11396
rect 37716 11340 37726 11396
rect 38322 11340 38332 11396
rect 38388 11340 38780 11396
rect 38836 11340 39452 11396
rect 39508 11340 39518 11396
rect 39676 11340 40236 11396
rect 40292 11340 40302 11396
rect 41906 11340 41916 11396
rect 41972 11340 42476 11396
rect 42532 11340 42542 11396
rect 43026 11340 43036 11396
rect 43092 11340 43820 11396
rect 43876 11340 43886 11396
rect 4498 11228 4508 11284
rect 4564 11228 5516 11284
rect 5572 11228 5582 11284
rect 12898 11228 12908 11284
rect 12964 11228 13356 11284
rect 13412 11228 13422 11284
rect 13682 11228 13692 11284
rect 13748 11228 15260 11284
rect 15316 11228 15326 11284
rect 15558 11228 15596 11284
rect 15652 11228 15662 11284
rect 35522 11228 35532 11284
rect 35588 11228 35980 11284
rect 36036 11228 37100 11284
rect 37156 11228 37166 11284
rect 37660 11172 37716 11340
rect 37874 11228 37884 11284
rect 37940 11228 38668 11284
rect 38724 11228 38734 11284
rect 39330 11228 39340 11284
rect 39396 11228 42700 11284
rect 42756 11228 44044 11284
rect 44100 11228 44110 11284
rect 2818 11116 2828 11172
rect 2884 11116 4620 11172
rect 4676 11116 4686 11172
rect 15138 11116 15148 11172
rect 15204 11116 16044 11172
rect 16100 11116 17388 11172
rect 17444 11116 17454 11172
rect 27234 11116 27244 11172
rect 27300 11116 28364 11172
rect 28420 11116 28430 11172
rect 32498 11116 32508 11172
rect 32564 11116 33852 11172
rect 33908 11116 33918 11172
rect 37660 11116 38220 11172
rect 38276 11116 38286 11172
rect 41010 11116 41020 11172
rect 41076 11116 42028 11172
rect 42084 11116 42364 11172
rect 42420 11116 42924 11172
rect 42980 11116 42990 11172
rect 29026 11004 29036 11060
rect 29092 11004 35532 11060
rect 35588 11004 35598 11060
rect 37314 11004 37324 11060
rect 37380 11004 37436 11060
rect 37492 11004 37502 11060
rect 38770 11004 38780 11060
rect 38836 11004 39340 11060
rect 39396 11004 43260 11060
rect 43316 11004 43326 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 27234 10892 27244 10948
rect 27300 10892 31388 10948
rect 31444 10892 31454 10948
rect 31938 10892 31948 10948
rect 32004 10892 33068 10948
rect 33124 10892 33134 10948
rect 36530 10892 36540 10948
rect 36596 10892 36988 10948
rect 37044 10892 37054 10948
rect 37202 10892 37212 10948
rect 37268 10892 39900 10948
rect 39956 10892 39966 10948
rect 2482 10780 2492 10836
rect 2548 10780 5292 10836
rect 5348 10780 5358 10836
rect 32498 10780 32508 10836
rect 32564 10780 35756 10836
rect 35812 10780 36428 10836
rect 36484 10780 36494 10836
rect 39414 10780 39452 10836
rect 39508 10780 39518 10836
rect 40786 10780 40796 10836
rect 40852 10780 42364 10836
rect 42420 10780 42430 10836
rect 7970 10668 7980 10724
rect 8036 10668 8540 10724
rect 8596 10668 20524 10724
rect 20580 10668 20590 10724
rect 27682 10668 27692 10724
rect 27748 10668 28028 10724
rect 28084 10668 28094 10724
rect 28354 10668 28364 10724
rect 28420 10668 28430 10724
rect 36306 10668 36316 10724
rect 36372 10668 45836 10724
rect 45892 10668 45902 10724
rect 28364 10612 28420 10668
rect 36316 10612 36372 10668
rect 10882 10556 10892 10612
rect 10948 10556 11788 10612
rect 11844 10556 12684 10612
rect 12740 10556 12750 10612
rect 15362 10556 15372 10612
rect 15428 10556 15820 10612
rect 15876 10556 15886 10612
rect 16594 10556 16604 10612
rect 16660 10556 18396 10612
rect 18452 10556 21644 10612
rect 21700 10556 21710 10612
rect 28364 10556 29372 10612
rect 29428 10556 29438 10612
rect 31266 10556 31276 10612
rect 31332 10556 33068 10612
rect 33124 10556 33134 10612
rect 35746 10556 35756 10612
rect 35812 10556 36372 10612
rect 36530 10556 36540 10612
rect 36596 10556 37548 10612
rect 37604 10556 37614 10612
rect 38612 10556 39340 10612
rect 39396 10556 39406 10612
rect 39554 10556 39564 10612
rect 39620 10556 40348 10612
rect 40404 10556 40414 10612
rect 42130 10556 42140 10612
rect 42196 10556 42588 10612
rect 42644 10556 42654 10612
rect 9426 10444 9436 10500
rect 9492 10444 11004 10500
rect 11060 10444 11070 10500
rect 12338 10444 12348 10500
rect 12404 10444 12908 10500
rect 12964 10444 12974 10500
rect 30594 10444 30604 10500
rect 30660 10444 32172 10500
rect 32228 10444 32238 10500
rect 37622 10444 37660 10500
rect 37716 10444 37726 10500
rect 38612 10388 38668 10556
rect 28476 10332 38668 10388
rect 28476 10276 28532 10332
rect 27682 10220 27692 10276
rect 27748 10220 28476 10276
rect 28532 10220 28542 10276
rect 38770 10220 38780 10276
rect 38836 10220 42252 10276
rect 42308 10220 42318 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 35634 10108 35644 10164
rect 35700 10108 39004 10164
rect 39060 10108 39070 10164
rect 25330 9996 25340 10052
rect 25396 9996 27132 10052
rect 27188 9996 29260 10052
rect 29316 9996 31276 10052
rect 31332 9996 31342 10052
rect 31490 9996 31500 10052
rect 31556 9996 31612 10052
rect 31668 9996 31678 10052
rect 33282 9996 33292 10052
rect 33348 9996 34748 10052
rect 34804 9996 37436 10052
rect 37492 9996 37502 10052
rect 38882 9996 38892 10052
rect 38948 9996 40012 10052
rect 40068 9996 40078 10052
rect 40338 9996 40348 10052
rect 40404 9996 42812 10052
rect 42868 9996 42878 10052
rect 11442 9884 11452 9940
rect 11508 9884 12012 9940
rect 12068 9884 12078 9940
rect 13010 9884 13020 9940
rect 13076 9884 21308 9940
rect 21364 9884 21374 9940
rect 24210 9884 24220 9940
rect 24276 9884 25004 9940
rect 25060 9884 25070 9940
rect 26562 9884 26572 9940
rect 26628 9884 26908 9940
rect 31154 9884 31164 9940
rect 31220 9884 32508 9940
rect 32564 9884 32956 9940
rect 33012 9884 34412 9940
rect 34468 9884 34478 9940
rect 39442 9884 39452 9940
rect 39508 9884 40908 9940
rect 40964 9884 42028 9940
rect 42084 9884 42094 9940
rect 7074 9772 7084 9828
rect 7140 9772 8428 9828
rect 11890 9772 11900 9828
rect 11956 9772 12236 9828
rect 12292 9772 13468 9828
rect 13524 9772 13534 9828
rect 8372 9716 8428 9772
rect 8372 9660 12348 9716
rect 12404 9660 15596 9716
rect 15652 9660 15662 9716
rect 25218 9660 25228 9716
rect 25284 9660 26348 9716
rect 26404 9660 26414 9716
rect 26852 9604 26908 9884
rect 38882 9772 38892 9828
rect 38948 9772 39900 9828
rect 39956 9772 39966 9828
rect 40114 9772 40124 9828
rect 40180 9772 40460 9828
rect 40516 9772 40526 9828
rect 39666 9660 39676 9716
rect 39732 9660 40012 9716
rect 40068 9660 40796 9716
rect 40852 9660 40862 9716
rect 7522 9548 7532 9604
rect 7588 9548 8428 9604
rect 8484 9548 8494 9604
rect 16594 9548 16604 9604
rect 16660 9548 18172 9604
rect 18228 9548 18238 9604
rect 22754 9548 22764 9604
rect 22820 9548 23436 9604
rect 23492 9548 23502 9604
rect 26852 9548 28140 9604
rect 28196 9548 30940 9604
rect 30996 9548 37100 9604
rect 37156 9548 37436 9604
rect 37492 9548 37502 9604
rect 37846 9548 37884 9604
rect 37940 9548 37950 9604
rect 39554 9548 39564 9604
rect 39620 9548 40684 9604
rect 40740 9548 40750 9604
rect 41906 9548 41916 9604
rect 41972 9548 43596 9604
rect 43652 9548 43662 9604
rect 44790 9548 44828 9604
rect 44884 9548 44894 9604
rect 45826 9548 45836 9604
rect 45892 9548 45902 9604
rect 7746 9436 7756 9492
rect 7812 9436 9436 9492
rect 9492 9436 9502 9492
rect 35522 9436 35532 9492
rect 35588 9436 38668 9492
rect 38994 9436 39004 9492
rect 39060 9436 41132 9492
rect 41188 9436 41198 9492
rect 41346 9436 41356 9492
rect 41412 9436 43932 9492
rect 43988 9436 43998 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 38612 9380 38668 9436
rect 45836 9380 45892 9548
rect 22194 9324 22204 9380
rect 22260 9324 26908 9380
rect 34290 9324 34300 9380
rect 34356 9324 38164 9380
rect 38612 9324 45892 9380
rect 11218 9212 11228 9268
rect 11284 9212 11788 9268
rect 11844 9212 11854 9268
rect 14130 9212 14140 9268
rect 14196 9212 14700 9268
rect 14756 9212 16212 9268
rect 21410 9212 21420 9268
rect 21476 9212 24780 9268
rect 24836 9212 25228 9268
rect 25284 9212 25294 9268
rect 16156 9156 16212 9212
rect 26852 9156 26908 9324
rect 27346 9212 27356 9268
rect 27412 9212 27916 9268
rect 27972 9212 31164 9268
rect 31220 9212 31230 9268
rect 33618 9212 33628 9268
rect 33684 9212 34524 9268
rect 34580 9212 34590 9268
rect 38108 9156 38164 9324
rect 39330 9212 39340 9268
rect 39396 9212 40236 9268
rect 40292 9212 41804 9268
rect 41860 9212 41870 9268
rect 7634 9100 7644 9156
rect 7700 9100 10108 9156
rect 10164 9100 10174 9156
rect 11330 9100 11340 9156
rect 11396 9100 13804 9156
rect 13860 9100 15148 9156
rect 15204 9100 15214 9156
rect 16156 9100 16716 9156
rect 16772 9100 16782 9156
rect 24994 9100 25004 9156
rect 25060 9100 26012 9156
rect 26068 9100 26078 9156
rect 26852 9100 30156 9156
rect 30212 9100 31388 9156
rect 31444 9100 31454 9156
rect 33628 9100 35756 9156
rect 35812 9100 35822 9156
rect 38108 9100 43036 9156
rect 43092 9100 46172 9156
rect 46228 9100 46238 9156
rect 9090 8988 9100 9044
rect 9156 8988 9548 9044
rect 9604 8988 9614 9044
rect 12674 8988 12684 9044
rect 12740 8988 13692 9044
rect 13748 8988 13758 9044
rect 16156 8932 16212 9100
rect 33628 9044 33684 9100
rect 24322 8988 24332 9044
rect 24388 8988 25564 9044
rect 25620 8988 27580 9044
rect 27636 8988 27646 9044
rect 30482 8988 30492 9044
rect 30548 8988 33684 9044
rect 33842 8988 33852 9044
rect 33908 8988 37100 9044
rect 37156 8988 37772 9044
rect 37828 8988 37838 9044
rect 38322 8988 38332 9044
rect 38388 8988 39116 9044
rect 39172 8988 41468 9044
rect 41524 8988 41534 9044
rect 6402 8876 6412 8932
rect 6468 8876 9660 8932
rect 9716 8876 9726 8932
rect 9874 8876 9884 8932
rect 9940 8876 11788 8932
rect 11844 8876 13020 8932
rect 13076 8876 13086 8932
rect 13234 8876 13244 8932
rect 13300 8876 14588 8932
rect 14644 8876 14654 8932
rect 16146 8876 16156 8932
rect 16212 8876 16222 8932
rect 16482 8876 16492 8932
rect 16548 8876 18172 8932
rect 18228 8876 18238 8932
rect 28466 8876 28476 8932
rect 28532 8876 31724 8932
rect 31780 8876 33068 8932
rect 33124 8876 33134 8932
rect 37650 8876 37660 8932
rect 37716 8876 39788 8932
rect 39844 8876 39854 8932
rect 40002 8876 40012 8932
rect 40068 8876 41132 8932
rect 41188 8876 41198 8932
rect 14466 8764 14476 8820
rect 14532 8764 14644 8820
rect 24434 8764 24444 8820
rect 24500 8764 29820 8820
rect 29876 8764 29886 8820
rect 31602 8764 31612 8820
rect 31668 8764 32284 8820
rect 32340 8764 32350 8820
rect 35074 8764 35084 8820
rect 35140 8764 38668 8820
rect 40114 8764 40124 8820
rect 40180 8764 40190 8820
rect 40870 8764 40908 8820
rect 40964 8764 40974 8820
rect 8866 8652 8876 8708
rect 8932 8652 9884 8708
rect 9940 8652 9950 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 8418 8540 8428 8596
rect 8484 8540 9436 8596
rect 9492 8540 9502 8596
rect 14588 8484 14644 8764
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 37846 8540 37884 8596
rect 37940 8540 37950 8596
rect 38612 8484 38668 8764
rect 1810 8428 1820 8484
rect 1876 8428 3612 8484
rect 3668 8428 3678 8484
rect 8978 8428 8988 8484
rect 9044 8428 10108 8484
rect 10164 8428 14644 8484
rect 27458 8428 27468 8484
rect 27524 8428 27534 8484
rect 34290 8428 34300 8484
rect 34356 8428 35532 8484
rect 35588 8428 36092 8484
rect 36148 8428 36158 8484
rect 38612 8428 38892 8484
rect 38948 8428 38958 8484
rect 3266 8316 3276 8372
rect 3332 8316 3500 8372
rect 3556 8316 3566 8372
rect 10658 8316 10668 8372
rect 10724 8316 11676 8372
rect 11732 8316 11742 8372
rect 14588 8260 14644 8428
rect 27468 8372 27524 8428
rect 14802 8316 14812 8372
rect 14868 8316 16380 8372
rect 16436 8316 16446 8372
rect 20738 8316 20748 8372
rect 20804 8316 21980 8372
rect 22036 8316 22046 8372
rect 23650 8316 23660 8372
rect 23716 8316 27524 8372
rect 27794 8316 27804 8372
rect 27860 8316 29596 8372
rect 29652 8316 29932 8372
rect 29988 8316 29998 8372
rect 32610 8316 32620 8372
rect 32676 8316 33404 8372
rect 33460 8316 33470 8372
rect 3602 8204 3612 8260
rect 3668 8204 4508 8260
rect 4564 8204 4574 8260
rect 11442 8204 11452 8260
rect 11508 8204 12124 8260
rect 12180 8204 12190 8260
rect 14588 8204 17948 8260
rect 18004 8204 19740 8260
rect 19796 8204 20860 8260
rect 20916 8204 21420 8260
rect 21476 8204 21486 8260
rect 24098 8204 24108 8260
rect 24164 8204 27692 8260
rect 27748 8204 27758 8260
rect 28354 8204 28364 8260
rect 28420 8204 29036 8260
rect 29092 8204 29102 8260
rect 33170 8204 33180 8260
rect 33236 8204 34076 8260
rect 34132 8204 34142 8260
rect 35074 8204 35084 8260
rect 35140 8204 37212 8260
rect 37268 8204 37278 8260
rect 38770 8204 38780 8260
rect 38836 8204 39676 8260
rect 39732 8204 39742 8260
rect 40124 8148 40180 8764
rect 43250 8428 43260 8484
rect 43316 8428 43932 8484
rect 43988 8428 43998 8484
rect 44258 8316 44268 8372
rect 44324 8316 46060 8372
rect 46116 8316 46126 8372
rect 42914 8204 42924 8260
rect 42980 8204 45052 8260
rect 45108 8204 45118 8260
rect 45378 8204 45388 8260
rect 45444 8204 45948 8260
rect 46004 8204 46014 8260
rect 3042 8092 3052 8148
rect 3108 8092 3948 8148
rect 4004 8092 4284 8148
rect 4340 8092 4350 8148
rect 12898 8092 12908 8148
rect 12964 8092 14140 8148
rect 14196 8092 14206 8148
rect 16818 8092 16828 8148
rect 16884 8092 20748 8148
rect 20804 8092 20814 8148
rect 20962 8092 20972 8148
rect 21028 8092 21756 8148
rect 21812 8092 21822 8148
rect 22866 8092 22876 8148
rect 22932 8092 23660 8148
rect 23716 8092 23726 8148
rect 25330 8092 25340 8148
rect 25396 8092 25788 8148
rect 25844 8092 26124 8148
rect 26180 8092 26190 8148
rect 28466 8092 28476 8148
rect 28532 8092 29260 8148
rect 29316 8092 29326 8148
rect 33506 8092 33516 8148
rect 33572 8092 33964 8148
rect 34020 8092 34030 8148
rect 40124 8092 41244 8148
rect 41300 8092 41310 8148
rect 20972 8036 21028 8092
rect 3490 7980 3500 8036
rect 3556 7980 4620 8036
rect 4676 7980 4686 8036
rect 12674 7980 12684 8036
rect 12740 7980 13804 8036
rect 13860 7980 15148 8036
rect 16370 7980 16380 8036
rect 16436 7980 17388 8036
rect 17444 7980 17454 8036
rect 20178 7980 20188 8036
rect 20244 7980 21028 8036
rect 23202 7980 23212 8036
rect 23268 7980 46284 8036
rect 46340 7980 47348 8036
rect 15092 7924 15148 7980
rect 15092 7868 16604 7924
rect 16660 7868 16670 7924
rect 21522 7868 21532 7924
rect 21588 7868 22316 7924
rect 22372 7868 24444 7924
rect 24500 7868 24510 7924
rect 30146 7868 30156 7924
rect 30212 7868 33292 7924
rect 33348 7868 33358 7924
rect 33516 7868 35084 7924
rect 35140 7868 35150 7924
rect 38546 7868 38556 7924
rect 38612 7868 39452 7924
rect 39508 7868 39788 7924
rect 39844 7868 39854 7924
rect 40002 7868 40012 7924
rect 40068 7868 41132 7924
rect 41188 7868 41198 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 33516 7812 33572 7868
rect 29474 7756 29484 7812
rect 29540 7756 33572 7812
rect 34066 7756 34076 7812
rect 34132 7756 39004 7812
rect 39060 7756 41468 7812
rect 41524 7756 41534 7812
rect 47292 7700 47348 7980
rect 18386 7644 18396 7700
rect 18452 7644 19852 7700
rect 19908 7644 19918 7700
rect 31826 7644 31836 7700
rect 31892 7644 32340 7700
rect 33170 7644 33180 7700
rect 33236 7644 34300 7700
rect 34356 7644 35084 7700
rect 35140 7644 35150 7700
rect 37426 7644 37436 7700
rect 37492 7644 44044 7700
rect 44100 7644 44110 7700
rect 47068 7644 47348 7700
rect 2930 7532 2940 7588
rect 2996 7532 4956 7588
rect 5012 7532 5022 7588
rect 16818 7532 16828 7588
rect 16884 7532 20412 7588
rect 20468 7532 20478 7588
rect 22194 7532 22204 7588
rect 22260 7532 22876 7588
rect 22932 7532 22942 7588
rect 32284 7476 32340 7644
rect 32498 7532 32508 7588
rect 32564 7532 33964 7588
rect 34020 7532 34030 7588
rect 39218 7532 39228 7588
rect 39284 7532 39900 7588
rect 39956 7532 39966 7588
rect 47068 7476 47124 7644
rect 47200 7476 48000 7504
rect 4498 7420 4508 7476
rect 4564 7420 5628 7476
rect 5684 7420 5694 7476
rect 10994 7420 11004 7476
rect 11060 7420 17388 7476
rect 17444 7420 17454 7476
rect 19618 7420 19628 7476
rect 19684 7420 20748 7476
rect 20804 7420 20814 7476
rect 22418 7420 22428 7476
rect 22484 7420 23380 7476
rect 24322 7420 24332 7476
rect 24388 7420 26012 7476
rect 26068 7420 26078 7476
rect 32274 7420 32284 7476
rect 32340 7420 33516 7476
rect 33572 7420 33582 7476
rect 37314 7420 37324 7476
rect 37380 7420 39564 7476
rect 39620 7420 44716 7476
rect 44772 7420 44782 7476
rect 47068 7420 48000 7476
rect 3826 7308 3836 7364
rect 3892 7308 5068 7364
rect 5124 7308 5134 7364
rect 11666 7308 11676 7364
rect 11732 7308 21644 7364
rect 21700 7308 21710 7364
rect 22642 7308 22652 7364
rect 22708 7308 22718 7364
rect 22652 7252 22708 7308
rect 23324 7252 23380 7420
rect 47200 7392 48000 7420
rect 24210 7308 24220 7364
rect 24276 7308 26796 7364
rect 26852 7308 28364 7364
rect 28420 7308 28430 7364
rect 34514 7308 34524 7364
rect 34580 7308 39340 7364
rect 39396 7308 39406 7364
rect 40562 7308 40572 7364
rect 40628 7308 43484 7364
rect 43540 7308 43550 7364
rect 18274 7196 18284 7252
rect 18340 7196 19068 7252
rect 19124 7196 19134 7252
rect 22652 7196 23100 7252
rect 23156 7196 23166 7252
rect 23314 7196 23324 7252
rect 23380 7196 23390 7252
rect 33394 7196 33404 7252
rect 33460 7196 34412 7252
rect 34468 7196 34478 7252
rect 39218 7196 39228 7252
rect 39284 7196 39294 7252
rect 39228 7140 39284 7196
rect 21410 7084 21420 7140
rect 21476 7084 23660 7140
rect 23716 7084 23726 7140
rect 35532 7084 39284 7140
rect 41010 7084 41020 7140
rect 41076 7084 41692 7140
rect 41748 7084 41758 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 12898 6972 12908 7028
rect 12964 6972 15148 7028
rect 15204 6972 15214 7028
rect 35532 6916 35588 7084
rect 37986 6972 37996 7028
rect 38052 6972 38444 7028
rect 38500 6972 38510 7028
rect 38882 6972 38892 7028
rect 38948 6972 39788 7028
rect 39844 6972 42028 7028
rect 42084 6972 42094 7028
rect 43922 6972 43932 7028
rect 43988 6972 45276 7028
rect 45332 6972 45342 7028
rect 2482 6860 2492 6916
rect 2548 6860 5740 6916
rect 5796 6860 5806 6916
rect 12226 6860 12236 6916
rect 12292 6860 15148 6916
rect 33954 6860 33964 6916
rect 34020 6860 35588 6916
rect 36418 6860 36428 6916
rect 36484 6860 41356 6916
rect 41412 6860 41422 6916
rect 42354 6860 42364 6916
rect 42420 6860 42812 6916
rect 42868 6860 43708 6916
rect 43764 6860 43774 6916
rect 44146 6860 44156 6916
rect 44212 6860 45500 6916
rect 45556 6860 45566 6916
rect 15092 6804 15148 6860
rect 2594 6748 2604 6804
rect 2660 6748 3276 6804
rect 3332 6748 4060 6804
rect 4116 6748 4396 6804
rect 4452 6748 4462 6804
rect 4946 6748 4956 6804
rect 5012 6748 5628 6804
rect 5684 6748 5694 6804
rect 10770 6748 10780 6804
rect 10836 6748 12572 6804
rect 12628 6748 12638 6804
rect 13122 6748 13132 6804
rect 13188 6748 14028 6804
rect 14084 6748 14094 6804
rect 15092 6748 15596 6804
rect 15652 6748 15662 6804
rect 16034 6748 16044 6804
rect 16100 6748 20972 6804
rect 21028 6748 21038 6804
rect 23426 6748 23436 6804
rect 23492 6748 23828 6804
rect 25554 6748 25564 6804
rect 25620 6748 26908 6804
rect 26964 6748 28252 6804
rect 28308 6748 30268 6804
rect 30324 6748 30334 6804
rect 33842 6748 33852 6804
rect 33908 6748 36092 6804
rect 36148 6748 36158 6804
rect 40450 6748 40460 6804
rect 40516 6748 45052 6804
rect 45108 6748 45118 6804
rect 23772 6692 23828 6748
rect 1698 6636 1708 6692
rect 1764 6636 2828 6692
rect 2884 6636 3612 6692
rect 3668 6636 3678 6692
rect 4162 6636 4172 6692
rect 4228 6636 5068 6692
rect 5124 6636 5134 6692
rect 8194 6636 8204 6692
rect 8260 6636 8428 6692
rect 12002 6636 12012 6692
rect 12068 6636 13244 6692
rect 13300 6636 14364 6692
rect 14420 6636 14430 6692
rect 21634 6636 21644 6692
rect 21700 6636 23548 6692
rect 23604 6636 23614 6692
rect 23772 6636 24780 6692
rect 24836 6636 24846 6692
rect 28130 6636 28140 6692
rect 28196 6636 29260 6692
rect 29316 6636 29326 6692
rect 30930 6636 30940 6692
rect 30996 6636 31948 6692
rect 32004 6636 32014 6692
rect 33618 6636 33628 6692
rect 33684 6636 33694 6692
rect 36194 6636 36204 6692
rect 36260 6636 39788 6692
rect 39844 6636 40908 6692
rect 40964 6636 40974 6692
rect 41122 6636 41132 6692
rect 41188 6636 41580 6692
rect 41636 6636 42812 6692
rect 42868 6636 42878 6692
rect 6626 6412 6636 6468
rect 6692 6412 7420 6468
rect 7476 6412 8204 6468
rect 8260 6412 8270 6468
rect 8372 6356 8428 6636
rect 12012 6580 12068 6636
rect 9426 6524 9436 6580
rect 9492 6524 12068 6580
rect 13010 6524 13020 6580
rect 13076 6524 14252 6580
rect 14308 6524 15708 6580
rect 15764 6524 15774 6580
rect 21522 6524 21532 6580
rect 21588 6524 26348 6580
rect 26404 6524 26414 6580
rect 28578 6524 28588 6580
rect 28644 6524 30044 6580
rect 30100 6524 30110 6580
rect 33628 6468 33684 6636
rect 36082 6524 36092 6580
rect 36148 6524 37772 6580
rect 37828 6524 37838 6580
rect 41010 6524 41020 6580
rect 41076 6524 42140 6580
rect 42196 6524 42206 6580
rect 42886 6524 42924 6580
rect 42980 6524 42990 6580
rect 10994 6412 11004 6468
rect 11060 6412 12124 6468
rect 12180 6412 12190 6468
rect 13906 6412 13916 6468
rect 13972 6412 14476 6468
rect 14532 6412 14542 6468
rect 14802 6412 14812 6468
rect 14868 6412 15260 6468
rect 15316 6412 15820 6468
rect 15876 6412 16716 6468
rect 16772 6412 16782 6468
rect 16930 6412 16940 6468
rect 16996 6412 19964 6468
rect 20020 6412 20030 6468
rect 20738 6412 20748 6468
rect 20804 6412 21868 6468
rect 21924 6412 21934 6468
rect 33628 6412 37212 6468
rect 37268 6412 37278 6468
rect 40674 6412 40684 6468
rect 40740 6412 42364 6468
rect 42420 6412 42430 6468
rect 44034 6412 44044 6468
rect 44100 6412 45948 6468
rect 46004 6412 46014 6468
rect 14476 6356 14532 6412
rect 8372 6300 8764 6356
rect 8820 6300 9548 6356
rect 9604 6300 9614 6356
rect 14476 6300 15484 6356
rect 15540 6300 16380 6356
rect 16436 6300 16446 6356
rect 39442 6300 39452 6356
rect 39508 6300 46060 6356
rect 46116 6300 46126 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 7074 6188 7084 6244
rect 7140 6188 8316 6244
rect 8372 6188 9100 6244
rect 9156 6188 9166 6244
rect 15092 6188 17724 6244
rect 17780 6188 18620 6244
rect 18676 6188 18686 6244
rect 32162 6188 32172 6244
rect 32228 6188 33740 6244
rect 33796 6188 33806 6244
rect 40450 6188 40460 6244
rect 40516 6188 42252 6244
rect 42308 6188 42318 6244
rect 15092 6132 15148 6188
rect 6178 6076 6188 6132
rect 6244 6076 7196 6132
rect 7252 6076 7262 6132
rect 13570 6076 13580 6132
rect 13636 6076 15148 6132
rect 15362 6076 15372 6132
rect 15428 6076 15438 6132
rect 18050 6076 18060 6132
rect 18116 6076 19628 6132
rect 19684 6076 20524 6132
rect 20580 6076 21308 6132
rect 21364 6076 21374 6132
rect 24770 6076 24780 6132
rect 24836 6076 26236 6132
rect 26292 6076 26302 6132
rect 36306 6076 36316 6132
rect 36372 6076 41020 6132
rect 41076 6076 41916 6132
rect 41972 6076 41982 6132
rect 7858 5964 7868 6020
rect 7924 5964 9100 6020
rect 9156 5964 12796 6020
rect 12852 5964 12862 6020
rect 15372 5908 15428 6076
rect 15810 5964 15820 6020
rect 15876 5964 16940 6020
rect 16996 5964 17006 6020
rect 12898 5852 12908 5908
rect 12964 5852 15428 5908
rect 16594 5852 16604 5908
rect 16660 5852 18396 5908
rect 18452 5852 18462 5908
rect 23202 5852 23212 5908
rect 23268 5852 25228 5908
rect 25284 5852 26012 5908
rect 26068 5852 26078 5908
rect 26236 5796 26292 6076
rect 39442 5964 39452 6020
rect 39508 5964 40348 6020
rect 40404 5964 40908 6020
rect 40964 5964 40974 6020
rect 26562 5852 26572 5908
rect 26628 5852 27580 5908
rect 27636 5852 27646 5908
rect 31826 5852 31836 5908
rect 31892 5852 33180 5908
rect 33236 5852 34300 5908
rect 34356 5852 34366 5908
rect 35298 5852 35308 5908
rect 35364 5852 35644 5908
rect 35700 5852 35710 5908
rect 40114 5852 40124 5908
rect 40180 5852 41692 5908
rect 41748 5852 42140 5908
rect 42196 5852 42206 5908
rect 9650 5740 9660 5796
rect 9716 5740 16492 5796
rect 16548 5740 16558 5796
rect 26236 5740 31948 5796
rect 32004 5740 32014 5796
rect 34626 5740 34636 5796
rect 34692 5740 35420 5796
rect 35476 5740 36204 5796
rect 36260 5740 36270 5796
rect 38612 5740 39228 5796
rect 39284 5740 39294 5796
rect 40786 5740 40796 5796
rect 40852 5740 42812 5796
rect 42868 5740 44940 5796
rect 44996 5740 45006 5796
rect 38612 5684 38668 5740
rect 4834 5628 4844 5684
rect 4900 5628 5516 5684
rect 5572 5628 5964 5684
rect 6020 5628 6030 5684
rect 8372 5628 9100 5684
rect 9156 5628 20748 5684
rect 20804 5628 20814 5684
rect 24210 5628 24220 5684
rect 24276 5628 38668 5684
rect 4946 5516 4956 5572
rect 5012 5516 6636 5572
rect 6692 5516 7084 5572
rect 7140 5516 7150 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 8372 5236 8428 5628
rect 16818 5516 16828 5572
rect 16884 5516 17052 5572
rect 17108 5516 17118 5572
rect 17266 5516 17276 5572
rect 17332 5516 18956 5572
rect 19012 5516 20636 5572
rect 20692 5516 22764 5572
rect 22820 5516 24836 5572
rect 25666 5516 25676 5572
rect 25732 5516 26684 5572
rect 26740 5516 26750 5572
rect 31602 5516 31612 5572
rect 31668 5516 32732 5572
rect 32788 5516 32798 5572
rect 24780 5460 24836 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 12562 5404 12572 5460
rect 12628 5404 14700 5460
rect 14756 5404 16156 5460
rect 16212 5404 16222 5460
rect 18610 5404 18620 5460
rect 18676 5404 23660 5460
rect 23716 5404 24556 5460
rect 24612 5404 24622 5460
rect 24780 5404 27468 5460
rect 27524 5404 27534 5460
rect 37874 5404 37884 5460
rect 37940 5404 38668 5460
rect 38612 5348 38668 5404
rect 17154 5292 17164 5348
rect 17220 5292 18508 5348
rect 18564 5292 18574 5348
rect 18834 5292 18844 5348
rect 18900 5292 20860 5348
rect 20916 5292 26516 5348
rect 27570 5292 27580 5348
rect 27636 5292 29148 5348
rect 29204 5292 29214 5348
rect 30370 5292 30380 5348
rect 30436 5292 31276 5348
rect 31332 5292 31342 5348
rect 34290 5292 34300 5348
rect 34356 5292 35196 5348
rect 35252 5292 35262 5348
rect 35970 5292 35980 5348
rect 36036 5292 37772 5348
rect 37828 5292 37838 5348
rect 38612 5292 40572 5348
rect 40628 5292 44828 5348
rect 44884 5292 44894 5348
rect 26460 5236 26516 5292
rect 4162 5180 4172 5236
rect 4228 5180 6300 5236
rect 6356 5180 7308 5236
rect 7364 5180 7374 5236
rect 8372 5180 8540 5236
rect 8596 5180 8606 5236
rect 9538 5180 9548 5236
rect 9604 5180 14700 5236
rect 14756 5180 14766 5236
rect 22866 5180 22876 5236
rect 22932 5180 24220 5236
rect 24276 5180 24286 5236
rect 26450 5180 26460 5236
rect 26516 5180 26526 5236
rect 34850 5180 34860 5236
rect 34916 5180 36316 5236
rect 36372 5180 36382 5236
rect 43474 5180 43484 5236
rect 43540 5180 44828 5236
rect 44884 5180 44894 5236
rect 5170 5068 5180 5124
rect 5236 5068 6076 5124
rect 6132 5068 6142 5124
rect 8372 5012 8428 5180
rect 10098 5068 10108 5124
rect 10164 5068 13132 5124
rect 13188 5068 13198 5124
rect 18050 5068 18060 5124
rect 18116 5068 19852 5124
rect 19908 5068 21308 5124
rect 21364 5068 21374 5124
rect 21970 5068 21980 5124
rect 22036 5068 23772 5124
rect 23828 5068 23838 5124
rect 25106 5068 25116 5124
rect 25172 5068 26236 5124
rect 26292 5068 26302 5124
rect 27234 5068 27244 5124
rect 27300 5068 27804 5124
rect 27860 5068 27870 5124
rect 30930 5068 30940 5124
rect 30996 5068 33068 5124
rect 33124 5068 34636 5124
rect 34692 5068 34702 5124
rect 36194 5068 36204 5124
rect 36260 5068 36988 5124
rect 37044 5068 37660 5124
rect 37716 5068 37726 5124
rect 43362 5068 43372 5124
rect 43428 5068 44268 5124
rect 44324 5068 44334 5124
rect 7746 4956 7756 5012
rect 7812 4956 8428 5012
rect 31714 4956 31724 5012
rect 31780 4956 32284 5012
rect 32340 4956 32350 5012
rect 33506 4956 33516 5012
rect 33572 4956 34524 5012
rect 34580 4956 35644 5012
rect 35700 4956 35710 5012
rect 35858 4956 35868 5012
rect 35924 4956 38668 5012
rect 42242 4956 42252 5012
rect 42308 4956 44380 5012
rect 44436 4956 44446 5012
rect 38612 4900 38668 4956
rect 8978 4844 8988 4900
rect 9044 4844 10556 4900
rect 10612 4844 10622 4900
rect 26898 4844 26908 4900
rect 26964 4844 29484 4900
rect 29540 4844 29550 4900
rect 35410 4844 35420 4900
rect 35476 4844 35644 4900
rect 35700 4844 35710 4900
rect 38612 4844 38780 4900
rect 38836 4844 39228 4900
rect 39284 4844 39294 4900
rect 41906 4844 41916 4900
rect 41972 4844 45836 4900
rect 45892 4844 45902 4900
rect 38322 4732 38332 4788
rect 38388 4732 38892 4788
rect 38948 4732 38958 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 23986 4620 23996 4676
rect 24052 4620 25228 4676
rect 25284 4620 27356 4676
rect 27412 4620 28588 4676
rect 28644 4620 28654 4676
rect 8642 4508 8652 4564
rect 8708 4508 13916 4564
rect 13972 4508 13982 4564
rect 29810 4508 29820 4564
rect 29876 4508 31836 4564
rect 31892 4508 31902 4564
rect 9650 4396 9660 4452
rect 9716 4396 12124 4452
rect 12180 4396 12190 4452
rect 13570 4396 13580 4452
rect 13636 4396 18732 4452
rect 18788 4396 18798 4452
rect 21522 4396 21532 4452
rect 21588 4396 24444 4452
rect 24500 4396 24510 4452
rect 35746 4396 35756 4452
rect 35812 4396 37100 4452
rect 37156 4396 37166 4452
rect 42466 4396 42476 4452
rect 42532 4396 45052 4452
rect 45108 4396 45118 4452
rect 7074 4284 7084 4340
rect 7140 4284 8764 4340
rect 8820 4284 9772 4340
rect 9828 4284 9838 4340
rect 28802 4284 28812 4340
rect 28868 4284 36260 4340
rect 36204 4228 36260 4284
rect 6290 4172 6300 4228
rect 6356 4172 7532 4228
rect 7588 4172 7598 4228
rect 13346 4172 13356 4228
rect 13412 4172 18732 4228
rect 18788 4172 18798 4228
rect 29250 4172 29260 4228
rect 29316 4172 31612 4228
rect 31668 4172 31678 4228
rect 34738 4172 34748 4228
rect 34804 4172 35980 4228
rect 36036 4172 36046 4228
rect 36194 4172 36204 4228
rect 36260 4172 36270 4228
rect 40002 4172 40012 4228
rect 40068 4172 40796 4228
rect 40852 4172 41580 4228
rect 41636 4172 41646 4228
rect 42690 4172 42700 4228
rect 42756 4172 43260 4228
rect 43316 4172 43326 4228
rect 34066 4060 34076 4116
rect 34132 4060 44604 4116
rect 44660 4060 44670 4116
rect 35970 3948 35980 4004
rect 36036 3948 38892 4004
rect 38948 3948 38958 4004
rect 39218 3948 39228 4004
rect 39284 3948 42812 4004
rect 42868 3948 42878 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 40310 3836 40348 3892
rect 40404 3836 40414 3892
rect 42886 3836 42924 3892
rect 42980 3836 42990 3892
rect 8754 3724 8764 3780
rect 8820 3724 14588 3780
rect 14644 3724 14654 3780
rect 31378 3724 31388 3780
rect 31444 3724 35980 3780
rect 36036 3724 36046 3780
rect 36194 3724 36204 3780
rect 36260 3724 43764 3780
rect 20066 3612 20076 3668
rect 20132 3612 21868 3668
rect 21924 3612 21934 3668
rect 26674 3612 26684 3668
rect 26740 3612 27580 3668
rect 27636 3612 28140 3668
rect 28196 3612 28206 3668
rect 30930 3612 30940 3668
rect 30996 3612 36988 3668
rect 37044 3612 37054 3668
rect 38742 3612 38780 3668
rect 38836 3612 38846 3668
rect 43708 3556 43764 3724
rect 16034 3500 16044 3556
rect 16100 3500 17612 3556
rect 17668 3500 17678 3556
rect 23986 3500 23996 3556
rect 24052 3500 32172 3556
rect 32228 3500 32238 3556
rect 35186 3500 35196 3556
rect 35252 3500 39564 3556
rect 39620 3500 39630 3556
rect 43698 3500 43708 3556
rect 43764 3500 43774 3556
rect 8642 3388 8652 3444
rect 8708 3388 10444 3444
rect 10500 3388 10510 3444
rect 11554 3388 11564 3444
rect 11620 3388 13692 3444
rect 13748 3388 13758 3444
rect 26002 3388 26012 3444
rect 26068 3388 27804 3444
rect 27860 3388 27870 3444
rect 29362 3388 29372 3444
rect 29428 3388 33740 3444
rect 33796 3388 33806 3444
rect 36418 3388 36428 3444
rect 36484 3388 38444 3444
rect 38500 3388 39116 3444
rect 39172 3388 39182 3444
rect 23090 3276 23100 3332
rect 23156 3276 25340 3332
rect 25396 3276 25406 3332
rect 26226 3276 26236 3332
rect 26292 3276 27020 3332
rect 27076 3276 27086 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 47200 2772 48000 2800
rect 43362 2716 43372 2772
rect 43428 2716 48000 2772
rect 47200 2688 48000 2716
<< via3 >>
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 30604 44268 30660 44324
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 43596 43372 43652 43428
rect 30716 43260 30772 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 30716 41020 30772 41076
rect 34188 40908 34244 40964
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 31612 40684 31668 40740
rect 20188 40572 20244 40628
rect 29708 40460 29764 40516
rect 30716 40460 30772 40516
rect 20188 40348 20244 40404
rect 34300 40348 34356 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 33964 39900 34020 39956
rect 31612 39564 31668 39620
rect 29708 39340 29764 39396
rect 34076 39228 34132 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 34636 39116 34692 39172
rect 26908 39004 26964 39060
rect 34076 38780 34132 38836
rect 26908 38668 26964 38724
rect 17164 38444 17220 38500
rect 34636 38444 34692 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 34300 38220 34356 38276
rect 34188 38108 34244 38164
rect 33964 37884 34020 37940
rect 43596 37884 43652 37940
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 17052 36652 17108 36708
rect 34860 36540 34916 36596
rect 17388 36428 17444 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 17164 35980 17220 36036
rect 17388 35980 17444 36036
rect 30604 35980 30660 36036
rect 17052 35868 17108 35924
rect 31164 35756 31220 35812
rect 45836 35308 45892 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 34972 35084 35028 35140
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 26908 34412 26964 34468
rect 17500 34300 17556 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 25676 33740 25732 33796
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 34860 33516 34916 33572
rect 45836 33516 45892 33572
rect 34972 33404 35028 33460
rect 17500 33068 17556 33124
rect 22876 32956 22932 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 26572 32732 26628 32788
rect 38444 32508 38500 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 38444 32284 38500 32340
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 31164 30716 31220 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 22764 30156 22820 30212
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 25452 29596 25508 29652
rect 11676 29484 11732 29540
rect 25452 29260 25508 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 22652 28588 22708 28644
rect 26236 28364 26292 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 11676 28140 11732 28196
rect 32508 28028 32564 28084
rect 41244 27804 41300 27860
rect 41916 27580 41972 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 26908 27356 26964 27412
rect 22652 27244 22708 27300
rect 41244 26796 41300 26852
rect 26572 26684 26628 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 41916 26572 41972 26628
rect 22764 26348 22820 26404
rect 26236 26348 26292 26404
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 43372 25564 43428 25620
rect 32508 25452 32564 25508
rect 25676 25116 25732 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 38108 24892 38164 24948
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 22876 23884 22932 23940
rect 43372 23884 43428 23940
rect 8428 23548 8484 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 22540 23436 22596 23492
rect 31724 23212 31780 23268
rect 30940 22988 30996 23044
rect 38108 22876 38164 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 8428 21420 8484 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 31724 20636 31780 20692
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 31724 20188 31780 20244
rect 33740 19964 33796 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 33740 18172 33796 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 20524 17388 20580 17444
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 34972 17164 35028 17220
rect 31724 16940 31780 16996
rect 20524 16604 20580 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 30044 15932 30100 15988
rect 34972 15932 35028 15988
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 31612 15484 31668 15540
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 30044 14364 30100 14420
rect 30940 14364 30996 14420
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 37884 13244 37940 13300
rect 39788 12684 39844 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 37884 12348 37940 12404
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 15596 11676 15652 11732
rect 37660 11564 37716 11620
rect 37436 11340 37492 11396
rect 15596 11228 15652 11284
rect 39340 11228 39396 11284
rect 37436 11004 37492 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 39452 10780 39508 10836
rect 39340 10556 39396 10612
rect 37660 10444 37716 10500
rect 38780 10220 38836 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 31612 9996 31668 10052
rect 40012 9996 40068 10052
rect 40348 9996 40404 10052
rect 40908 9884 40964 9940
rect 15596 9660 15652 9716
rect 37884 9548 37940 9604
rect 44828 9548 44884 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 41132 8876 41188 8932
rect 40908 8764 40964 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 37884 8540 37940 8596
rect 39452 7868 39508 7924
rect 40012 7868 40068 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 39788 6972 39844 7028
rect 41132 6636 41188 6692
rect 42924 6524 42980 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 35644 5852 35700 5908
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 44828 5180 44884 5236
rect 35644 4844 35700 4900
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 36204 4172 36260 4228
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 40348 3836 40404 3892
rect 42924 3836 42980 3892
rect 36204 3724 36260 3780
rect 38780 3612 38836 3668
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 44716 4768 44748
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 19808 43932 20128 44748
rect 35168 44716 35488 44748
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 30604 44324 30660 44334
rect 20188 40628 20244 40638
rect 20188 40404 20244 40572
rect 20188 40338 20244 40348
rect 29708 40516 29764 40526
rect 29708 39396 29764 40460
rect 29708 39330 29764 39340
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 17164 38500 17220 38510
rect 17052 36708 17108 36718
rect 17052 35924 17108 36652
rect 17164 36036 17220 38444
rect 19808 37660 20128 39172
rect 26908 39060 26964 39070
rect 26908 38724 26964 39004
rect 26908 38658 26964 38668
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 17164 35970 17220 35980
rect 17388 36484 17444 36494
rect 17388 36036 17444 36428
rect 17388 35970 17444 35980
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 17052 35858 17108 35868
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 34524 20128 36036
rect 30604 36036 30660 44268
rect 30716 43316 30772 43326
rect 30716 41076 30772 43260
rect 30716 40516 30772 41020
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 34188 40964 34244 40974
rect 30716 40450 30772 40460
rect 31612 40740 31668 40750
rect 31612 39620 31668 40684
rect 31612 39554 31668 39564
rect 33964 39956 34020 39966
rect 33964 37940 34020 39900
rect 34076 39284 34132 39294
rect 34076 38836 34132 39228
rect 34076 38770 34132 38780
rect 34188 38164 34244 40908
rect 34300 40404 34356 40414
rect 34300 38276 34356 40348
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 34636 39172 34692 39182
rect 34636 38500 34692 39116
rect 34636 38434 34692 38444
rect 35168 38444 35488 39956
rect 34300 38210 34356 38220
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 34188 38098 34244 38108
rect 33964 37874 34020 37884
rect 35168 36876 35488 38388
rect 43596 43428 43652 43438
rect 43596 37940 43652 43372
rect 43596 37874 43652 37884
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 30604 35970 30660 35980
rect 34860 36596 34916 36606
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 31164 35812 31220 35822
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 17500 34356 17556 34366
rect 17500 33124 17556 34300
rect 17500 33058 17556 33068
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 32956 20128 34468
rect 26908 34468 26964 34478
rect 25676 33796 25732 33806
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 22876 33012 22932 33022
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 11676 29540 11732 29550
rect 11676 28196 11732 29484
rect 11676 28130 11732 28140
rect 19808 28252 20128 29764
rect 22764 30212 22820 30222
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19808 26684 20128 28196
rect 22652 28644 22708 28654
rect 22652 27300 22708 28588
rect 22652 26908 22708 27244
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 8428 23604 8484 23614
rect 8428 21476 8484 23548
rect 8428 21410 8484 21420
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 22540 26852 22708 26908
rect 22540 23492 22596 26852
rect 22764 26404 22820 30156
rect 22764 26338 22820 26348
rect 22876 23940 22932 32956
rect 25452 29652 25508 29662
rect 25452 29316 25508 29596
rect 25452 29250 25508 29260
rect 25676 25172 25732 33740
rect 26572 32788 26628 32798
rect 26236 28420 26292 28430
rect 26236 26404 26292 28364
rect 26572 26740 26628 32732
rect 26908 27412 26964 34412
rect 31164 30772 31220 35756
rect 34860 33572 34916 36540
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 34860 33506 34916 33516
rect 34972 35140 35028 35150
rect 34972 33460 35028 35084
rect 34972 33394 35028 33404
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 31164 30706 31220 30716
rect 35168 32172 35488 33684
rect 45836 35364 45892 35374
rect 45836 33572 45892 35308
rect 45836 33506 45892 33516
rect 38444 32564 38500 32574
rect 38444 32340 38500 32508
rect 38444 32274 38500 32284
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 26908 27346 26964 27356
rect 32508 28084 32564 28094
rect 26572 26674 26628 26684
rect 26236 26338 26292 26348
rect 32508 25508 32564 28028
rect 32508 25442 32564 25452
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 41244 27860 41300 27870
rect 41244 26852 41300 27804
rect 41244 26786 41300 26796
rect 41916 27636 41972 27646
rect 41916 26628 41972 27580
rect 41916 26562 41972 26572
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 25676 25106 25732 25116
rect 22876 23874 22932 23884
rect 35168 24332 35488 25844
rect 43372 25620 43428 25630
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 22540 23426 22596 23436
rect 31724 23268 31780 23278
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 30940 23044 30996 23054
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20524 17444 20580 17454
rect 20524 16660 20580 17388
rect 20524 16594 20580 16604
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 30044 15988 30100 15998
rect 30044 14420 30100 15932
rect 30044 14354 30100 14364
rect 30940 14420 30996 22988
rect 31724 20692 31780 23212
rect 31724 20244 31780 20636
rect 31724 16996 31780 20188
rect 35168 22764 35488 24276
rect 38108 24948 38164 24958
rect 38108 22932 38164 24892
rect 43372 23940 43428 25564
rect 43372 23874 43428 23884
rect 38108 22866 38164 22876
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 33740 20020 33796 20030
rect 33740 18228 33796 19964
rect 33740 18162 33796 18172
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 31724 16930 31780 16940
rect 34972 17220 35028 17230
rect 34972 15988 35028 17164
rect 34972 15922 35028 15932
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 30940 14354 30996 14364
rect 31612 15540 31668 15550
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 15596 11732 15652 11742
rect 15596 11284 15652 11676
rect 15596 9716 15652 11228
rect 15596 9650 15652 9660
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 9436 20128 10948
rect 31612 10052 31668 15484
rect 31612 9986 31668 9996
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 37884 13300 37940 13310
rect 37884 12404 37940 13244
rect 37660 11620 37716 11630
rect 37436 11396 37492 11406
rect 37436 11060 37492 11340
rect 37436 10994 37492 11004
rect 37660 10500 37716 11564
rect 37660 10434 37716 10444
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 37884 9604 37940 12348
rect 39788 12740 39844 12750
rect 39340 11284 39396 11294
rect 39340 10612 39396 11228
rect 39340 10546 39396 10556
rect 39452 10836 39508 10846
rect 37884 8596 37940 9548
rect 37884 8530 37940 8540
rect 38780 10276 38836 10286
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35644 5908 35700 5918
rect 35644 4900 35700 5852
rect 35644 4834 35700 4844
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 36204 4228 36260 4238
rect 36204 3780 36260 4172
rect 36204 3714 36260 3724
rect 38780 3668 38836 10220
rect 39452 7924 39508 10780
rect 39452 7858 39508 7868
rect 39788 7028 39844 12684
rect 40012 10052 40068 10062
rect 40012 7924 40068 9996
rect 40012 7858 40068 7868
rect 40348 10052 40404 10062
rect 39788 6962 39844 6972
rect 40348 3892 40404 9996
rect 40908 9940 40964 9950
rect 40908 8820 40964 9884
rect 44828 9604 44884 9614
rect 40908 8754 40964 8764
rect 41132 8932 41188 8942
rect 41132 6692 41188 8876
rect 41132 6626 41188 6636
rect 40348 3826 40404 3836
rect 42924 6580 42980 6590
rect 42924 3892 42980 6524
rect 44828 5236 44884 9548
rect 44828 5170 44884 5180
rect 42924 3826 42980 3836
rect 38780 3602 38836 3612
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1024_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 -1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1025_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19040 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1026_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1027_
timestamp 1698431365
transform 1 0 21728 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1028_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1029_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1030_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26880 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1031_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1032_
timestamp 1698431365
transform -1 0 23856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1033_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1034_
timestamp 1698431365
transform 1 0 17808 0 -1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1035_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1036_
timestamp 1698431365
transform -1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1037_
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1038_
timestamp 1698431365
transform 1 0 17808 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1039_
timestamp 1698431365
transform -1 0 19488 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1040_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1041_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17920 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1043_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1044_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform 1 0 17808 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1046_
timestamp 1698431365
transform 1 0 21728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698431365
transform 1 0 28000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1049_
timestamp 1698431365
transform -1 0 29792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1050_
timestamp 1698431365
transform 1 0 32256 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1051_
timestamp 1698431365
transform -1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1052_
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1053_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1054_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1055_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1056_
timestamp 1698431365
transform -1 0 31024 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1057_
timestamp 1698431365
transform -1 0 21728 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1058_
timestamp 1698431365
transform 1 0 22848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1059_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1060_
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1061_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29344 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1062_
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1063_
timestamp 1698431365
transform -1 0 30688 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1064_
timestamp 1698431365
transform 1 0 29680 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1065_
timestamp 1698431365
transform 1 0 30688 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1066_
timestamp 1698431365
transform -1 0 33152 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1067_
timestamp 1698431365
transform 1 0 29792 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1068_
timestamp 1698431365
transform 1 0 29120 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1069_
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1070_
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1071_
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform -1 0 46144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1073_
timestamp 1698431365
transform 1 0 34160 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1074_
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1075_
timestamp 1698431365
transform -1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1076_
timestamp 1698431365
transform 1 0 25200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1077_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1078_
timestamp 1698431365
transform -1 0 28112 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1079_
timestamp 1698431365
transform 1 0 29344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1080_
timestamp 1698431365
transform 1 0 31024 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1081_
timestamp 1698431365
transform -1 0 20944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1082_
timestamp 1698431365
transform 1 0 21392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1083_
timestamp 1698431365
transform 1 0 31024 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1084_
timestamp 1698431365
transform -1 0 32704 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1085_
timestamp 1698431365
transform -1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1086_
timestamp 1698431365
transform -1 0 33936 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1087_
timestamp 1698431365
transform -1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1088_
timestamp 1698431365
transform -1 0 36064 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1089_
timestamp 1698431365
transform 1 0 35504 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1090_
timestamp 1698431365
transform -1 0 35056 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1091_
timestamp 1698431365
transform -1 0 39536 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1092_
timestamp 1698431365
transform -1 0 26432 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1093_
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698431365
transform 1 0 31920 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1095_
timestamp 1698431365
transform 1 0 22512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1096_
timestamp 1698431365
transform -1 0 24416 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1097_
timestamp 1698431365
transform 1 0 20944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1098_
timestamp 1698431365
transform 1 0 31136 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1099_
timestamp 1698431365
transform -1 0 23856 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1100_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1101_
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1102_
timestamp 1698431365
transform -1 0 23856 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1103_
timestamp 1698431365
transform 1 0 22176 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1104_
timestamp 1698431365
transform -1 0 25536 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1105_
timestamp 1698431365
transform 1 0 34720 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1107_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1108_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1109_
timestamp 1698431365
transform -1 0 15232 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1110_
timestamp 1698431365
transform 1 0 16016 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1698431365
transform 1 0 20608 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1112_
timestamp 1698431365
transform 1 0 34608 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1113_
timestamp 1698431365
transform -1 0 24640 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1114_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1115_
timestamp 1698431365
transform -1 0 23408 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1116_
timestamp 1698431365
transform -1 0 35728 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1117_
timestamp 1698431365
transform -1 0 22848 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1118_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1119_
timestamp 1698431365
transform 1 0 21952 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1120_
timestamp 1698431365
transform 1 0 21392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1121_
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1122_
timestamp 1698431365
transform 1 0 17360 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1123_
timestamp 1698431365
transform -1 0 19600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1124_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698431365
transform 1 0 19824 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1126_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1127_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1128_
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1129_
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 19824 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1131_
timestamp 1698431365
transform -1 0 15568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1132_
timestamp 1698431365
transform -1 0 14336 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1133_
timestamp 1698431365
transform -1 0 18704 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform 1 0 19376 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1135_
timestamp 1698431365
transform -1 0 18928 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1136_
timestamp 1698431365
transform -1 0 18592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1137_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 -1 12544
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1138_
timestamp 1698431365
transform -1 0 16464 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1139_
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1140_
timestamp 1698431365
transform -1 0 18144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1141_
timestamp 1698431365
transform -1 0 17696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1142_
timestamp 1698431365
transform -1 0 15904 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1143_
timestamp 1698431365
transform -1 0 16464 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform 1 0 15344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1145_
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1146_
timestamp 1698431365
transform -1 0 15904 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1147_
timestamp 1698431365
transform -1 0 14000 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1148_
timestamp 1698431365
transform -1 0 15568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform -1 0 13888 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1150_
timestamp 1698431365
transform -1 0 13104 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1151_
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1152_
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1153_
timestamp 1698431365
transform 1 0 10528 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1154_
timestamp 1698431365
transform -1 0 11536 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1155_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11984 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1156_
timestamp 1698431365
transform -1 0 10640 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1157_
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1158_
timestamp 1698431365
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1159_
timestamp 1698431365
transform 1 0 11536 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1160_
timestamp 1698431365
transform 1 0 13552 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1161_
timestamp 1698431365
transform -1 0 29904 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform -1 0 26768 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1163_
timestamp 1698431365
transform -1 0 27776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1164_
timestamp 1698431365
transform -1 0 28448 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1165_
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698431365
transform -1 0 22400 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1167_
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1169_
timestamp 1698431365
transform -1 0 28000 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1170_
timestamp 1698431365
transform -1 0 23856 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1171_
timestamp 1698431365
transform -1 0 26880 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1172_
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1173_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1174_
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1175_
timestamp 1698431365
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1176_
timestamp 1698431365
transform -1 0 14336 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1177_
timestamp 1698431365
transform -1 0 25536 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform 1 0 17584 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1179_
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1180_
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1181_
timestamp 1698431365
transform 1 0 20160 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1182_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1183_
timestamp 1698431365
transform 1 0 19376 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1184_
timestamp 1698431365
transform -1 0 18592 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1185_
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698431365
transform 1 0 13440 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1187_
timestamp 1698431365
transform -1 0 16016 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1188_
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1698431365
transform -1 0 14896 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1190_
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1191_
timestamp 1698431365
transform -1 0 12432 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1192_
timestamp 1698431365
transform 1 0 14112 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1193_
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1194_
timestamp 1698431365
transform 1 0 16016 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1195_
timestamp 1698431365
transform -1 0 9856 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1196_
timestamp 1698431365
transform 1 0 18256 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1197_
timestamp 1698431365
transform -1 0 13776 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1198_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19488 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1199_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1200_
timestamp 1698431365
transform -1 0 16912 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1201_
timestamp 1698431365
transform -1 0 17024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform -1 0 15456 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1204_
timestamp 1698431365
transform -1 0 5712 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1205_
timestamp 1698431365
transform -1 0 6384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1206_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1207_
timestamp 1698431365
transform -1 0 5264 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1208_
timestamp 1698431365
transform 1 0 4368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1209_
timestamp 1698431365
transform -1 0 7840 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1211_
timestamp 1698431365
transform -1 0 5824 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1212_
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1213_
timestamp 1698431365
transform 1 0 4368 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1214_
timestamp 1698431365
transform -1 0 7168 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1215_
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1216_
timestamp 1698431365
transform 1 0 7392 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1217_
timestamp 1698431365
transform -1 0 7952 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1218_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1219_
timestamp 1698431365
transform -1 0 9856 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1220_
timestamp 1698431365
transform 1 0 8176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1221_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1222_
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1698431365
transform -1 0 34160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1224_
timestamp 1698431365
transform 1 0 21728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1698431365
transform -1 0 33488 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1227_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1228_
timestamp 1698431365
transform -1 0 30800 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1229_
timestamp 1698431365
transform -1 0 33936 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1230_
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1231_
timestamp 1698431365
transform -1 0 34944 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1232_
timestamp 1698431365
transform 1 0 34944 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1233_
timestamp 1698431365
transform -1 0 34048 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1234_
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1235_
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1236_
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1237_
timestamp 1698431365
transform -1 0 39088 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1238_
timestamp 1698431365
transform -1 0 40208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1239_
timestamp 1698431365
transform 1 0 42336 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1240_
timestamp 1698431365
transform -1 0 42000 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1242_
timestamp 1698431365
transform 1 0 43232 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1243_
timestamp 1698431365
transform -1 0 43904 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1244_
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1245_
timestamp 1698431365
transform 1 0 42224 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1246_
timestamp 1698431365
transform -1 0 43120 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1247_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1249_
timestamp 1698431365
transform 1 0 30016 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1251_
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1252_
timestamp 1698431365
transform -1 0 33936 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1253_
timestamp 1698431365
transform -1 0 33376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1254_
timestamp 1698431365
transform -1 0 32256 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1255_
timestamp 1698431365
transform -1 0 31472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1256_
timestamp 1698431365
transform -1 0 34944 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1257_
timestamp 1698431365
transform -1 0 35840 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1258_
timestamp 1698431365
transform -1 0 34160 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1260_
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1261_
timestamp 1698431365
transform 1 0 30688 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_
timestamp 1698431365
transform -1 0 33824 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1263_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1264_
timestamp 1698431365
transform -1 0 34272 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1265_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1266_
timestamp 1698431365
transform 1 0 33040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1267_
timestamp 1698431365
transform -1 0 32480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1268_
timestamp 1698431365
transform -1 0 31920 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1269_
timestamp 1698431365
transform -1 0 30912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1270_
timestamp 1698431365
transform -1 0 33152 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1271_
timestamp 1698431365
transform -1 0 32928 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1272_
timestamp 1698431365
transform -1 0 31360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1273_
timestamp 1698431365
transform -1 0 34496 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1274_
timestamp 1698431365
transform -1 0 33936 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1275_
timestamp 1698431365
transform -1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1277_
timestamp 1698431365
transform 1 0 36960 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1278_
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1279_
timestamp 1698431365
transform -1 0 40432 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1280_
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1281_
timestamp 1698431365
transform -1 0 45136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1282_
timestamp 1698431365
transform -1 0 43344 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1283_
timestamp 1698431365
transform -1 0 44352 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1284_
timestamp 1698431365
transform 1 0 40208 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1285_
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1287_
timestamp 1698431365
transform 1 0 24192 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1289_
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1290_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1291_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1292_
timestamp 1698431365
transform 1 0 24864 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1293_
timestamp 1698431365
transform 1 0 25760 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1294_
timestamp 1698431365
transform 1 0 25872 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1295_
timestamp 1698431365
transform 1 0 23968 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform 1 0 29904 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1298_
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1299_
timestamp 1698431365
transform -1 0 28672 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1300_
timestamp 1698431365
transform -1 0 4480 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1301_
timestamp 1698431365
transform 1 0 3696 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1302_
timestamp 1698431365
transform -1 0 3696 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1303_
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1304_
timestamp 1698431365
transform 1 0 3472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1305_
timestamp 1698431365
transform -1 0 3472 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1306_
timestamp 1698431365
transform -1 0 5040 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1307_
timestamp 1698431365
transform 1 0 6160 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698431365
transform 1 0 3248 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1309_
timestamp 1698431365
transform -1 0 3136 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1310_
timestamp 1698431365
transform 1 0 3472 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1311_
timestamp 1698431365
transform -1 0 3248 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform 1 0 4816 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1313_
timestamp 1698431365
transform 1 0 4816 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1314_
timestamp 1698431365
transform 1 0 5712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1315_
timestamp 1698431365
transform -1 0 5264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1316_
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1317_
timestamp 1698431365
transform 1 0 15232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1318_
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1319_
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1320_
timestamp 1698431365
transform -1 0 22400 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1321_
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1322_
timestamp 1698431365
transform 1 0 5824 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1323_
timestamp 1698431365
transform 1 0 7280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1324_
timestamp 1698431365
transform 1 0 6832 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1325_
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1326_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1327_
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform -1 0 22736 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1329_
timestamp 1698431365
transform -1 0 21728 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1330_
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1331_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1332_
timestamp 1698431365
transform -1 0 36400 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1333_
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1334_
timestamp 1698431365
transform 1 0 19712 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1335_
timestamp 1698431365
transform -1 0 23184 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1336_
timestamp 1698431365
transform -1 0 20608 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1337_
timestamp 1698431365
transform 1 0 21504 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1698431365
transform -1 0 19600 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1339_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1340_
timestamp 1698431365
transform -1 0 16016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1341_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1342_
timestamp 1698431365
transform -1 0 15680 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1343_
timestamp 1698431365
transform -1 0 18816 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1344_
timestamp 1698431365
transform -1 0 18256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1345_
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1346_
timestamp 1698431365
transform 1 0 18368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform 1 0 22400 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1349_
timestamp 1698431365
transform 1 0 22736 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1351_
timestamp 1698431365
transform 1 0 25984 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1352_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1353_
timestamp 1698431365
transform 1 0 22400 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1354_
timestamp 1698431365
transform 1 0 23408 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1355_
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1356_
timestamp 1698431365
transform -1 0 20384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1357_
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1358_
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1359_
timestamp 1698431365
transform -1 0 32144 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1698431365
transform -1 0 26656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1361_
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1362_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1363_
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1364_
timestamp 1698431365
transform -1 0 7728 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1366_
timestamp 1698431365
transform -1 0 29904 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1367_
timestamp 1698431365
transform -1 0 26544 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1698431365
transform -1 0 27776 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698431365
transform -1 0 25760 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1370_
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1371_
timestamp 1698431365
transform -1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1372_
timestamp 1698431365
transform 1 0 18144 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1373_
timestamp 1698431365
transform -1 0 17024 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1374_
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1375_
timestamp 1698431365
transform -1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1376_
timestamp 1698431365
transform -1 0 20832 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1377_
timestamp 1698431365
transform -1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1378_
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1379_
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1380_
timestamp 1698431365
transform 1 0 25424 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1381_
timestamp 1698431365
transform -1 0 24752 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1382_
timestamp 1698431365
transform 1 0 29904 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform -1 0 38192 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1385_
timestamp 1698431365
transform 1 0 37744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1386_
timestamp 1698431365
transform 1 0 35392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1387_
timestamp 1698431365
transform -1 0 38864 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1698431365
transform -1 0 37520 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform 1 0 35056 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1390_
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1391_
timestamp 1698431365
transform -1 0 37520 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1698431365
transform 1 0 35168 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1393_
timestamp 1698431365
transform 1 0 35392 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1394_
timestamp 1698431365
transform -1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1698431365
transform 1 0 38192 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1698431365
transform -1 0 35168 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1397_
timestamp 1698431365
transform 1 0 38864 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1398_
timestamp 1698431365
transform -1 0 39536 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1399_
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1400_
timestamp 1698431365
transform 1 0 39648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1401_
timestamp 1698431365
transform -1 0 46368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1402_
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1403_
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1404_
timestamp 1698431365
transform -1 0 45696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1405_
timestamp 1698431365
transform 1 0 44016 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1406_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1407_
timestamp 1698431365
transform -1 0 46144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1408_
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1409_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1410_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1411_
timestamp 1698431365
transform -1 0 15008 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform -1 0 5600 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1413_
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1414_
timestamp 1698431365
transform 1 0 8736 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1415_
timestamp 1698431365
transform -1 0 10752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1416_
timestamp 1698431365
transform -1 0 10304 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1417_
timestamp 1698431365
transform -1 0 7504 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1418_
timestamp 1698431365
transform -1 0 5488 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1419_
timestamp 1698431365
transform 1 0 12432 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1420_
timestamp 1698431365
transform -1 0 10976 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1421_
timestamp 1698431365
transform 1 0 2576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1422_
timestamp 1698431365
transform -1 0 2576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1423_
timestamp 1698431365
transform -1 0 12208 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1424_
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1425_
timestamp 1698431365
transform 1 0 2800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1426_
timestamp 1698431365
transform -1 0 4928 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1427_
timestamp 1698431365
transform -1 0 3472 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform 1 0 3248 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1429_
timestamp 1698431365
transform 1 0 4144 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform -1 0 4480 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform -1 0 3248 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1432_
timestamp 1698431365
transform 1 0 2800 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1433_
timestamp 1698431365
transform 1 0 3472 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1434_
timestamp 1698431365
transform 1 0 3696 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1435_
timestamp 1698431365
transform 1 0 6160 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1436_
timestamp 1698431365
transform -1 0 6160 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1437_
timestamp 1698431365
transform 1 0 33264 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1438_
timestamp 1698431365
transform -1 0 35168 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1439_
timestamp 1698431365
transform -1 0 34384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1440_
timestamp 1698431365
transform 1 0 33824 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1441_
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1442_
timestamp 1698431365
transform -1 0 33376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1443_
timestamp 1698431365
transform -1 0 32592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_
timestamp 1698431365
transform 1 0 29680 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1445_
timestamp 1698431365
transform -1 0 32144 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1446_
timestamp 1698431365
transform 1 0 31584 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 29008 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1448_
timestamp 1698431365
transform 1 0 29120 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1449_
timestamp 1698431365
transform -1 0 30576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1450_
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1451_
timestamp 1698431365
transform -1 0 30464 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1452_
timestamp 1698431365
transform 1 0 27888 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 30016 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1454_
timestamp 1698431365
transform 1 0 24976 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1455_
timestamp 1698431365
transform 1 0 27552 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1456_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1457_
timestamp 1698431365
transform -1 0 31584 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1458_
timestamp 1698431365
transform 1 0 30128 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1459_
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1460_
timestamp 1698431365
transform -1 0 33600 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1461_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32144 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1462_
timestamp 1698431365
transform 1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1463_
timestamp 1698431365
transform -1 0 45472 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1464_
timestamp 1698431365
transform 1 0 43904 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1465_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43120 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1466_
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1467_
timestamp 1698431365
transform -1 0 38528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1468_
timestamp 1698431365
transform -1 0 36624 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1469_
timestamp 1698431365
transform -1 0 43344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1470_
timestamp 1698431365
transform 1 0 38528 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1471_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41664 0 1 36064
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1472_
timestamp 1698431365
transform 1 0 34944 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1473_
timestamp 1698431365
transform -1 0 46256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1474_
timestamp 1698431365
transform -1 0 46368 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1475_
timestamp 1698431365
transform 1 0 44576 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1698431365
transform -1 0 46368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1477_
timestamp 1698431365
transform 1 0 42672 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1478_
timestamp 1698431365
transform 1 0 42896 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1480_
timestamp 1698431365
transform -1 0 43008 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1481_
timestamp 1698431365
transform -1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1482_
timestamp 1698431365
transform 1 0 34832 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1483_
timestamp 1698431365
transform -1 0 39984 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1484_
timestamp 1698431365
transform -1 0 37296 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1485_
timestamp 1698431365
transform 1 0 41664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1486_
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1487_
timestamp 1698431365
transform -1 0 45696 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1488_
timestamp 1698431365
transform 1 0 35728 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1490_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1491_
timestamp 1698431365
transform -1 0 27552 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1492_
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1493_
timestamp 1698431365
transform 1 0 33376 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1494_
timestamp 1698431365
transform 1 0 28336 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1495_
timestamp 1698431365
transform -1 0 34832 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1496_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31472 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1497_
timestamp 1698431365
transform 1 0 30352 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1498_
timestamp 1698431365
transform 1 0 31136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform 1 0 43456 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1500_
timestamp 1698431365
transform -1 0 15120 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1501_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25648 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1502_
timestamp 1698431365
transform 1 0 13552 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1503_
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1504_
timestamp 1698431365
transform -1 0 26880 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1505_
timestamp 1698431365
transform -1 0 34048 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1506_
timestamp 1698431365
transform -1 0 32480 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1507_
timestamp 1698431365
transform -1 0 32816 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1508_
timestamp 1698431365
transform -1 0 10304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1509_
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1511_
timestamp 1698431365
transform 1 0 7616 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1512_
timestamp 1698431365
transform -1 0 9072 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1513_
timestamp 1698431365
transform -1 0 33824 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1514_
timestamp 1698431365
transform -1 0 26432 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1515_
timestamp 1698431365
transform -1 0 24416 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1516_
timestamp 1698431365
transform 1 0 30576 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1517_
timestamp 1698431365
transform 1 0 35392 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1518_
timestamp 1698431365
transform -1 0 32480 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1519_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698431365
transform 1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1521_
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1522_
timestamp 1698431365
transform 1 0 28336 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1523_
timestamp 1698431365
transform 1 0 31024 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1524_
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform -1 0 30128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform 1 0 31696 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1527_
timestamp 1698431365
transform -1 0 29904 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1528_
timestamp 1698431365
transform 1 0 30352 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1529_
timestamp 1698431365
transform 1 0 30800 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1530_
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1531_
timestamp 1698431365
transform 1 0 30352 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1532_
timestamp 1698431365
transform -1 0 32144 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 32032 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1534_
timestamp 1698431365
transform 1 0 29120 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1535_
timestamp 1698431365
transform 1 0 32144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1536_
timestamp 1698431365
transform 1 0 34944 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1538_
timestamp 1698431365
transform 1 0 33040 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1539_
timestamp 1698431365
transform -1 0 33936 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1542_
timestamp 1698431365
transform 1 0 34272 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1543_
timestamp 1698431365
transform 1 0 35168 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1544_
timestamp 1698431365
transform -1 0 37296 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1698431365
transform 1 0 33712 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1546_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1547_
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1548_
timestamp 1698431365
transform -1 0 38192 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1549_
timestamp 1698431365
transform -1 0 37072 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1550_
timestamp 1698431365
transform -1 0 38416 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1551_
timestamp 1698431365
transform -1 0 37520 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1552_
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1554_
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1555_
timestamp 1698431365
transform -1 0 39648 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1556_
timestamp 1698431365
transform 1 0 44128 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1557_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1558_
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1559_
timestamp 1698431365
transform -1 0 42784 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1560_
timestamp 1698431365
transform 1 0 42560 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1561_
timestamp 1698431365
transform 1 0 45696 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1562_
timestamp 1698431365
transform -1 0 44240 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1563_
timestamp 1698431365
transform -1 0 45808 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1564_
timestamp 1698431365
transform -1 0 45584 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1565_
timestamp 1698431365
transform 1 0 44016 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform 1 0 45584 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698431365
transform -1 0 44464 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1568_
timestamp 1698431365
transform 1 0 45360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1569_
timestamp 1698431365
transform -1 0 10640 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1571_
timestamp 1698431365
transform -1 0 9520 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1572_
timestamp 1698431365
transform 1 0 7616 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1573_
timestamp 1698431365
transform 1 0 6720 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1574_
timestamp 1698431365
transform 1 0 5824 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1575_
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1576_
timestamp 1698431365
transform 1 0 7392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 7840 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform -1 0 8848 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1580_
timestamp 1698431365
transform -1 0 6608 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform 1 0 6048 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1584_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1698431365
transform -1 0 10864 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1587_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1588_
timestamp 1698431365
transform 1 0 7616 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698431365
transform 1 0 8176 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1590_
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1591_
timestamp 1698431365
transform -1 0 9072 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1698431365
transform -1 0 5488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1698431365
transform -1 0 7280 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1595_
timestamp 1698431365
transform -1 0 6272 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1596_
timestamp 1698431365
transform -1 0 6944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1698431365
transform 1 0 2576 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1698431365
transform -1 0 4928 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1698431365
transform 1 0 3696 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1600_
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1698431365
transform -1 0 2576 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1602_
timestamp 1698431365
transform -1 0 6048 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1603_
timestamp 1698431365
transform -1 0 2800 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1698431365
transform 1 0 2576 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1698431365
transform -1 0 6048 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1606_
timestamp 1698431365
transform -1 0 4032 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform -1 0 6160 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1698431365
transform -1 0 5712 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform -1 0 6048 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1610_
timestamp 1698431365
transform -1 0 5488 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1611_
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 5152 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1614_
timestamp 1698431365
transform 1 0 3024 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1615_
timestamp 1698431365
transform 1 0 3584 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1698431365
transform 1 0 2912 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1698431365
transform -1 0 4928 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1618_
timestamp 1698431365
transform -1 0 4368 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1698431365
transform -1 0 6048 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1698431365
transform 1 0 2352 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1621_
timestamp 1698431365
transform 1 0 3472 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1622_
timestamp 1698431365
transform -1 0 6160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform 1 0 2912 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform -1 0 2352 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1625_
timestamp 1698431365
transform -1 0 10080 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1626_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1628_
timestamp 1698431365
transform -1 0 7392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 6048 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1630_
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698431365
transform -1 0 8736 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1698431365
transform 1 0 6160 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1633_
timestamp 1698431365
transform 1 0 6720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform 1 0 7168 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform 1 0 7616 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1636_
timestamp 1698431365
transform 1 0 7728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 7504 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1638_
timestamp 1698431365
transform 1 0 6944 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 8064 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1640_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3248 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1641_
timestamp 1698431365
transform 1 0 4368 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1642_
timestamp 1698431365
transform -1 0 7280 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform -1 0 6608 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1644_
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1645_
timestamp 1698431365
transform 1 0 7392 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1646_
timestamp 1698431365
transform -1 0 7504 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1647_
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1648_
timestamp 1698431365
transform -1 0 7616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1649_
timestamp 1698431365
transform -1 0 6944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1651_
timestamp 1698431365
transform -1 0 28784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1698431365
transform -1 0 27440 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1653_
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1654_
timestamp 1698431365
transform 1 0 27216 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform -1 0 27440 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1698431365
transform -1 0 29568 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1698431365
transform -1 0 27104 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1658_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29680 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1659_
timestamp 1698431365
transform -1 0 27888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1660_
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1662_
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1663_
timestamp 1698431365
transform -1 0 23184 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1664_
timestamp 1698431365
transform 1 0 22288 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform 1 0 23408 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1666_
timestamp 1698431365
transform -1 0 26656 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1667_
timestamp 1698431365
transform 1 0 23968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1668_
timestamp 1698431365
transform -1 0 25760 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1669_
timestamp 1698431365
transform -1 0 28112 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1670_
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1671_
timestamp 1698431365
transform -1 0 26880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1672_
timestamp 1698431365
transform -1 0 25984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1673_
timestamp 1698431365
transform -1 0 25984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform -1 0 26768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1675_
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1676_
timestamp 1698431365
transform -1 0 27440 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1677_
timestamp 1698431365
transform -1 0 26880 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1678_
timestamp 1698431365
transform -1 0 24416 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1679_
timestamp 1698431365
transform -1 0 23184 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform -1 0 25984 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1681_
timestamp 1698431365
transform -1 0 15120 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1682_
timestamp 1698431365
transform 1 0 13216 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1683_
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1684_
timestamp 1698431365
transform -1 0 11760 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1685_
timestamp 1698431365
transform -1 0 10752 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1686_
timestamp 1698431365
transform 1 0 11312 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1687_
timestamp 1698431365
transform 1 0 10864 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1688_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1689_
timestamp 1698431365
transform 1 0 11760 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1690_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1691_
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1692_
timestamp 1698431365
transform -1 0 32816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1693_
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1694_
timestamp 1698431365
transform -1 0 40096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1695_
timestamp 1698431365
transform -1 0 39088 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1696_
timestamp 1698431365
transform 1 0 42672 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1697_
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1698_
timestamp 1698431365
transform 1 0 38752 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1699_
timestamp 1698431365
transform 1 0 40768 0 1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform -1 0 39760 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1701_
timestamp 1698431365
transform -1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1702_
timestamp 1698431365
transform -1 0 37296 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1703_
timestamp 1698431365
transform -1 0 44240 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform 1 0 33824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1705_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1706_
timestamp 1698431365
transform -1 0 38528 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform 1 0 37968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1708_
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1709_
timestamp 1698431365
transform -1 0 39424 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1711_
timestamp 1698431365
transform -1 0 39536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1712_
timestamp 1698431365
transform -1 0 38416 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1713_
timestamp 1698431365
transform 1 0 38080 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1714_
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1715_
timestamp 1698431365
transform -1 0 40544 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1716_
timestamp 1698431365
transform -1 0 40992 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1717_
timestamp 1698431365
transform 1 0 38752 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1718_
timestamp 1698431365
transform -1 0 42896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1719_
timestamp 1698431365
transform -1 0 43344 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1720_
timestamp 1698431365
transform 1 0 41104 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1721_
timestamp 1698431365
transform 1 0 37296 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1722_
timestamp 1698431365
transform -1 0 37968 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1723_
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1724_
timestamp 1698431365
transform -1 0 41888 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1725_
timestamp 1698431365
transform -1 0 44128 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1726_
timestamp 1698431365
transform -1 0 42560 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1727_
timestamp 1698431365
transform -1 0 40432 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1728_
timestamp 1698431365
transform -1 0 40432 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1729_
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1730_
timestamp 1698431365
transform 1 0 36960 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 35728 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1732_
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1733_
timestamp 1698431365
transform -1 0 40320 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1734_
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1735_
timestamp 1698431365
transform 1 0 40432 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1736_
timestamp 1698431365
transform -1 0 39760 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1737_
timestamp 1698431365
transform -1 0 40432 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1739_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1740_
timestamp 1698431365
transform -1 0 35056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1741_
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1742_
timestamp 1698431365
transform -1 0 37408 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1743_
timestamp 1698431365
transform -1 0 34720 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1744_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1745_
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1698431365
transform 1 0 34720 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1747_
timestamp 1698431365
transform -1 0 35392 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1749_
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1750_
timestamp 1698431365
transform 1 0 38528 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1751_
timestamp 1698431365
transform 1 0 39088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1752_
timestamp 1698431365
transform 1 0 39872 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1753_
timestamp 1698431365
transform -1 0 38192 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1754_
timestamp 1698431365
transform 1 0 41104 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1755_
timestamp 1698431365
transform 1 0 41552 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1756_
timestamp 1698431365
transform 1 0 42000 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform 1 0 43568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1758_
timestamp 1698431365
transform 1 0 42000 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1759_
timestamp 1698431365
transform 1 0 43344 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1760_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1761_
timestamp 1698431365
transform -1 0 35616 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform -1 0 28784 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1763_
timestamp 1698431365
transform 1 0 40992 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1764_
timestamp 1698431365
transform 1 0 41216 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1765_
timestamp 1698431365
transform 1 0 40880 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1766_
timestamp 1698431365
transform 1 0 42112 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1767_
timestamp 1698431365
transform -1 0 44128 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1768_
timestamp 1698431365
transform 1 0 30240 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1769_
timestamp 1698431365
transform 1 0 42560 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1770_
timestamp 1698431365
transform -1 0 41216 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1771_
timestamp 1698431365
transform 1 0 43344 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1772_
timestamp 1698431365
transform -1 0 46256 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1773_
timestamp 1698431365
transform 1 0 41776 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1774_
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1775_
timestamp 1698431365
transform -1 0 46256 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1776_
timestamp 1698431365
transform -1 0 40768 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1777_
timestamp 1698431365
transform 1 0 41888 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1778_
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1779_
timestamp 1698431365
transform -1 0 45696 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1780_
timestamp 1698431365
transform -1 0 41216 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 41328 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1782_
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1783_
timestamp 1698431365
transform 1 0 34944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform 1 0 41328 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1785_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1786_
timestamp 1698431365
transform -1 0 45360 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1787_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1788_
timestamp 1698431365
transform -1 0 38080 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1789_
timestamp 1698431365
transform -1 0 27104 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1790_
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1791_
timestamp 1698431365
transform -1 0 28000 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1792_
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1793_
timestamp 1698431365
transform 1 0 33936 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1795_
timestamp 1698431365
transform -1 0 40544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1796_
timestamp 1698431365
transform -1 0 40096 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1797_
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1798_
timestamp 1698431365
transform -1 0 44352 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1799_
timestamp 1698431365
transform 1 0 41328 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1800_
timestamp 1698431365
transform 1 0 42000 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1801_
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1802_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1803_
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1804_
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1805_
timestamp 1698431365
transform -1 0 40992 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1806_
timestamp 1698431365
transform -1 0 39088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1807_
timestamp 1698431365
transform 1 0 36624 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1808_
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1809_
timestamp 1698431365
transform 1 0 33264 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1810_
timestamp 1698431365
transform 1 0 34048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1811_
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1812_
timestamp 1698431365
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1813_
timestamp 1698431365
transform 1 0 34160 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_
timestamp 1698431365
transform -1 0 37744 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1815_
timestamp 1698431365
transform 1 0 36960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1816_
timestamp 1698431365
transform -1 0 38528 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1817_
timestamp 1698431365
transform -1 0 40208 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1818_
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1819_
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1820_
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1821_
timestamp 1698431365
transform -1 0 39648 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1822_
timestamp 1698431365
transform 1 0 38528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1823_
timestamp 1698431365
transform -1 0 46368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1824_
timestamp 1698431365
transform -1 0 46368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1825_
timestamp 1698431365
transform -1 0 44464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1826_
timestamp 1698431365
transform 1 0 39312 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1827_
timestamp 1698431365
transform 1 0 40768 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1828_
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1829_
timestamp 1698431365
transform -1 0 41776 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1830_
timestamp 1698431365
transform -1 0 40656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1831_
timestamp 1698431365
transform 1 0 39648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1832_
timestamp 1698431365
transform -1 0 45920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1698431365
transform -1 0 42896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1834_
timestamp 1698431365
transform -1 0 39424 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1835_
timestamp 1698431365
transform 1 0 39088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1836_
timestamp 1698431365
transform 1 0 39424 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1837_
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1838_
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1839_
timestamp 1698431365
transform -1 0 39200 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1840_
timestamp 1698431365
transform -1 0 40096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1841_
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1842_
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 41328 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1844_
timestamp 1698431365
transform 1 0 37856 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1845_
timestamp 1698431365
transform -1 0 40432 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1846_
timestamp 1698431365
transform 1 0 38752 0 -1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1847_
timestamp 1698431365
transform -1 0 40432 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1848_
timestamp 1698431365
transform -1 0 32032 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1849_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1850_
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1851_
timestamp 1698431365
transform -1 0 37520 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1852_
timestamp 1698431365
transform 1 0 37632 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1853_
timestamp 1698431365
transform -1 0 36624 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 35280 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1855_
timestamp 1698431365
transform 1 0 35168 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1856_
timestamp 1698431365
transform 1 0 36400 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1857_
timestamp 1698431365
transform -1 0 38976 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1858_
timestamp 1698431365
transform -1 0 35616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1859_
timestamp 1698431365
transform 1 0 35616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1860_
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1861_
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1862_
timestamp 1698431365
transform 1 0 37968 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1863_
timestamp 1698431365
transform 1 0 41664 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1864_
timestamp 1698431365
transform 1 0 41552 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1866_
timestamp 1698431365
transform -1 0 45472 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1867_
timestamp 1698431365
transform -1 0 44240 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1868_
timestamp 1698431365
transform 1 0 41216 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1869_
timestamp 1698431365
transform 1 0 43008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1870_
timestamp 1698431365
transform 1 0 41776 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1872_
timestamp 1698431365
transform 1 0 42000 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1873_
timestamp 1698431365
transform -1 0 43456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1874_
timestamp 1698431365
transform 1 0 43456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1875_
timestamp 1698431365
transform 1 0 42000 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1876_
timestamp 1698431365
transform -1 0 42560 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1877_
timestamp 1698431365
transform -1 0 45584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1878_
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1879_
timestamp 1698431365
transform -1 0 42000 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1880_
timestamp 1698431365
transform -1 0 45584 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1881_
timestamp 1698431365
transform 1 0 39872 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1882_
timestamp 1698431365
transform 1 0 40544 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1883_
timestamp 1698431365
transform -1 0 45472 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1884_
timestamp 1698431365
transform -1 0 44912 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1885_
timestamp 1698431365
transform -1 0 30800 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1886_
timestamp 1698431365
transform -1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1887_
timestamp 1698431365
transform -1 0 29792 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1888_
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1889_
timestamp 1698431365
transform -1 0 18704 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1890_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1891_
timestamp 1698431365
transform 1 0 22400 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1892_
timestamp 1698431365
transform -1 0 24864 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1893_
timestamp 1698431365
transform -1 0 13104 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1894_
timestamp 1698431365
transform -1 0 20384 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1895_
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1896_
timestamp 1698431365
transform 1 0 16800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1897_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1898_
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1899_
timestamp 1698431365
transform -1 0 17696 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1900_
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1901_
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1902_
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1903_
timestamp 1698431365
transform -1 0 18816 0 1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1905_
timestamp 1698431365
transform -1 0 22736 0 -1 39200
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1906_
timestamp 1698431365
transform -1 0 24864 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1907_
timestamp 1698431365
transform -1 0 17920 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1908_
timestamp 1698431365
transform -1 0 19152 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1909_
timestamp 1698431365
transform -1 0 18144 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1910_
timestamp 1698431365
transform -1 0 20944 0 1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1911_
timestamp 1698431365
transform 1 0 14336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1912_
timestamp 1698431365
transform 1 0 18816 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1914_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform -1 0 17920 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1916_
timestamp 1698431365
transform -1 0 22400 0 -1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1917_
timestamp 1698431365
transform 1 0 12880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1918_
timestamp 1698431365
transform -1 0 20944 0 1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1919_
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1920_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1921_
timestamp 1698431365
transform -1 0 20944 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1922_
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1923_
timestamp 1698431365
transform 1 0 12208 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1924_
timestamp 1698431365
transform 1 0 13328 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1925_
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1926_
timestamp 1698431365
transform -1 0 18816 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform -1 0 19712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1928_
timestamp 1698431365
transform -1 0 16016 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1698431365
transform -1 0 17024 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1930_
timestamp 1698431365
transform -1 0 18704 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1931_
timestamp 1698431365
transform -1 0 16688 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1932_
timestamp 1698431365
transform -1 0 15904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1933_
timestamp 1698431365
transform -1 0 14672 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1934_
timestamp 1698431365
transform -1 0 16016 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1935_
timestamp 1698431365
transform -1 0 14000 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1936_
timestamp 1698431365
transform -1 0 16128 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1937_
timestamp 1698431365
transform 1 0 15344 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1938_
timestamp 1698431365
transform 1 0 16128 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1939_
timestamp 1698431365
transform -1 0 16464 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1940_
timestamp 1698431365
transform -1 0 16352 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1941_
timestamp 1698431365
transform -1 0 15568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1942_
timestamp 1698431365
transform -1 0 15232 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1943_
timestamp 1698431365
transform -1 0 11648 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1944_
timestamp 1698431365
transform -1 0 14448 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform -1 0 14224 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1946_
timestamp 1698431365
transform -1 0 12096 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1947_
timestamp 1698431365
transform 1 0 9632 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1948_
timestamp 1698431365
transform -1 0 10304 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1949_
timestamp 1698431365
transform 1 0 10304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1950_
timestamp 1698431365
transform -1 0 10752 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1951_
timestamp 1698431365
transform 1 0 8960 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1952_
timestamp 1698431365
transform -1 0 10304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1953_
timestamp 1698431365
transform 1 0 9520 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1954_
timestamp 1698431365
transform 1 0 10864 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 9520 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1956_
timestamp 1698431365
transform 1 0 11088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 22960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1958_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 22848 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1960_
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1961_
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1962_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1963_
timestamp 1698431365
transform 1 0 18928 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1964_
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1965_
timestamp 1698431365
transform -1 0 12656 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1966_
timestamp 1698431365
transform 1 0 10080 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1967_
timestamp 1698431365
transform -1 0 14000 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1968_
timestamp 1698431365
transform 1 0 11424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1969_
timestamp 1698431365
transform -1 0 11424 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1970_
timestamp 1698431365
transform 1 0 14448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1971_
timestamp 1698431365
transform -1 0 13776 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1972_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1973_
timestamp 1698431365
transform 1 0 12880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform -1 0 14896 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1975_
timestamp 1698431365
transform 1 0 13664 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform 1 0 14560 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1977_
timestamp 1698431365
transform 1 0 14672 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1978_
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1979_
timestamp 1698431365
transform -1 0 13776 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1980_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1981_
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1982_
timestamp 1698431365
transform -1 0 12432 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1983_
timestamp 1698431365
transform -1 0 14896 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1698431365
transform -1 0 11424 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1985_
timestamp 1698431365
transform 1 0 42224 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1986_
timestamp 1698431365
transform -1 0 28784 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1987_
timestamp 1698431365
transform -1 0 26880 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1988_
timestamp 1698431365
transform -1 0 24416 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1989_
timestamp 1698431365
transform -1 0 23968 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1990_
timestamp 1698431365
transform -1 0 23744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1991_
timestamp 1698431365
transform 1 0 24416 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1992_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1993_
timestamp 1698431365
transform -1 0 25984 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform -1 0 24864 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1995_
timestamp 1698431365
transform -1 0 26544 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1996_
timestamp 1698431365
transform -1 0 27104 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1997_
timestamp 1698431365
transform -1 0 28000 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1998_
timestamp 1698431365
transform -1 0 27664 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 28000 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2000_
timestamp 1698431365
transform 1 0 29120 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2001_
timestamp 1698431365
transform -1 0 31024 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2003_
timestamp 1698431365
transform -1 0 31696 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2004_
timestamp 1698431365
transform 1 0 27776 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2005_
timestamp 1698431365
transform -1 0 26208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2006_
timestamp 1698431365
transform -1 0 30016 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2007_
timestamp 1698431365
transform -1 0 26656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2008_
timestamp 1698431365
transform 1 0 30576 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2009_
timestamp 1698431365
transform -1 0 30464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2010_
timestamp 1698431365
transform 1 0 29344 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2011_
timestamp 1698431365
transform -1 0 35056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2012_
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2013_
timestamp 1698431365
transform -1 0 34608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2014_
timestamp 1698431365
transform 1 0 31584 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2015_
timestamp 1698431365
transform -1 0 34608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2016_
timestamp 1698431365
transform -1 0 33936 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2017_
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2018_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2019_
timestamp 1698431365
transform -1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2020_
timestamp 1698431365
transform -1 0 32704 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2021_
timestamp 1698431365
transform -1 0 34272 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2022_
timestamp 1698431365
transform 1 0 14896 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2023_
timestamp 1698431365
transform -1 0 14672 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform 1 0 15456 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2025_
timestamp 1698431365
transform -1 0 11984 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2026_
timestamp 1698431365
transform -1 0 15232 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2027_
timestamp 1698431365
transform 1 0 12656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2028_
timestamp 1698431365
transform -1 0 11424 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2029_
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2030_
timestamp 1698431365
transform 1 0 9408 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2031_
timestamp 1698431365
transform 1 0 10304 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2032_
timestamp 1698431365
transform -1 0 10304 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2033_
timestamp 1698431365
transform 1 0 9968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2034_
timestamp 1698431365
transform -1 0 9184 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2035_
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2036_
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2037_
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2038_
timestamp 1698431365
transform -1 0 10752 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2039_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2040_
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1698431365
transform -1 0 11760 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2042_
timestamp 1698431365
transform -1 0 11872 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform -1 0 10528 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2044_
timestamp 1698431365
transform 1 0 11760 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2045_
timestamp 1698431365
transform -1 0 14000 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1698431365
transform -1 0 25984 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1698431365
transform -1 0 24528 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2048_
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2049_
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2050_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31584 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2051_
timestamp 1698431365
transform -1 0 32368 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2052_
timestamp 1698431365
transform -1 0 32816 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2053_
timestamp 1698431365
transform -1 0 31584 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2054_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2055_
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2056_
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2057_
timestamp 1698431365
transform 1 0 36176 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2058_
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2059_
timestamp 1698431365
transform 1 0 19600 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2060_
timestamp 1698431365
transform 1 0 21616 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2061_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2062_
timestamp 1698431365
transform -1 0 22288 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2063_
timestamp 1698431365
transform -1 0 23856 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2064_
timestamp 1698431365
transform -1 0 19376 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2065_
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2066_
timestamp 1698431365
transform 1 0 16128 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2067_
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2068_
timestamp 1698431365
transform 1 0 11648 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2069_
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2070_
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2071_
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2072_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2073_
timestamp 1698431365
transform -1 0 23744 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2074_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2075_
timestamp 1698431365
transform 1 0 16128 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2076_
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2077_
timestamp 1698431365
transform 1 0 9856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2078_
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2079_
timestamp 1698431365
transform 1 0 9520 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2080_
timestamp 1698431365
transform 1 0 13776 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_
timestamp 1698431365
transform 1 0 17808 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform 1 0 1904 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform -1 0 9184 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform -1 0 36400 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform -1 0 46368 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform -1 0 46368 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 29792 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform 1 0 29344 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform -1 0 36288 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 37408 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform -1 0 44464 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform 1 0 43120 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform 1 0 40656 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform -1 0 27328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform -1 0 32256 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2115_
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2118_
timestamp 1698431365
transform -1 0 4816 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform 1 0 5488 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2121_
timestamp 1698431365
transform -1 0 7280 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform -1 0 22960 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 13776 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 13776 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform -1 0 20496 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform -1 0 24416 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2130_
timestamp 1698431365
transform -1 0 28112 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2131_
timestamp 1698431365
transform -1 0 24864 0 -1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform 1 0 18144 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform 1 0 21056 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform 1 0 28560 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 5152 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform 1 0 15456 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform 1 0 13776 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform -1 0 29344 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform 1 0 22176 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 35616 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform 1 0 35056 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2146_
timestamp 1698431365
transform 1 0 37296 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698431365
transform 1 0 39088 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698431365
transform 1 0 43120 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698431365
transform 1 0 43120 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698431365
transform 1 0 9408 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2153_
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2155_
timestamp 1698431365
transform -1 0 4816 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2156_
timestamp 1698431365
transform -1 0 8736 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2157_
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2158_
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2159_
timestamp 1698431365
transform -1 0 28336 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2160_
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2161_
timestamp 1698431365
transform 1 0 24752 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2162_
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698431365
transform -1 0 36176 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2164_
timestamp 1698431365
transform -1 0 36176 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698431365
transform 1 0 36176 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2166_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2167_
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2168_
timestamp 1698431365
transform -1 0 42896 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2169_
timestamp 1698431365
transform -1 0 42560 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698431365
transform 1 0 39984 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698431365
transform 1 0 37296 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2173_
timestamp 1698431365
transform -1 0 44464 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2175_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698431365
transform -1 0 11760 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698431365
transform -1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698431365
transform -1 0 4816 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698431365
transform -1 0 4816 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698431365
transform 1 0 3472 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698431365
transform -1 0 10528 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698431365
transform -1 0 10528 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698431365
transform 1 0 5488 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698431365
transform -1 0 23184 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698431365
transform 1 0 23744 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698431365
transform 1 0 22848 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698431365
transform 1 0 21392 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698431365
transform 1 0 5488 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2199_
timestamp 1698431365
transform -1 0 15008 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698431365
transform 1 0 8624 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698431365
transform -1 0 12768 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698431365
transform -1 0 13552 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698431365
transform -1 0 41440 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698431365
transform -1 0 46368 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698431365
transform -1 0 46368 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2208_
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2209_
timestamp 1698431365
transform -1 0 46368 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2210_
timestamp 1698431365
transform -1 0 46368 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2211_
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2212_
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2213_
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2214_
timestamp 1698431365
transform -1 0 37968 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2215_
timestamp 1698431365
transform 1 0 23632 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2216_
timestamp 1698431365
transform 1 0 34384 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2217_
timestamp 1698431365
transform 1 0 30912 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2218_
timestamp 1698431365
transform 1 0 33264 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2219_
timestamp 1698431365
transform -1 0 40096 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2220_
timestamp 1698431365
transform -1 0 46368 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2221_
timestamp 1698431365
transform 1 0 43120 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2222_
timestamp 1698431365
transform -1 0 46368 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2223_
timestamp 1698431365
transform -1 0 46368 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2224_
timestamp 1698431365
transform -1 0 44464 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2225_
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2226_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2227_
timestamp 1698431365
transform 1 0 43120 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2228_
timestamp 1698431365
transform -1 0 29680 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2229_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2230_
timestamp 1698431365
transform -1 0 16800 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2231_
timestamp 1698431365
transform 1 0 13328 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2232_
timestamp 1698431365
transform 1 0 11648 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2233_
timestamp 1698431365
transform 1 0 15568 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2234_
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2235_
timestamp 1698431365
transform 1 0 9856 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2236_
timestamp 1698431365
transform 1 0 10528 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2237_
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2238_
timestamp 1698431365
transform 1 0 5712 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2239_
timestamp 1698431365
transform 1 0 5936 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2240_
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2241_
timestamp 1698431365
transform -1 0 21952 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2242_
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2243_
timestamp 1698431365
transform 1 0 13776 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2244_
timestamp 1698431365
transform 1 0 9184 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2245_
timestamp 1698431365
transform 1 0 10640 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2246_
timestamp 1698431365
transform 1 0 10528 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2247_
timestamp 1698431365
transform 1 0 10864 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2248_
timestamp 1698431365
transform 1 0 9856 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2249_
timestamp 1698431365
transform 1 0 9856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2250_
timestamp 1698431365
transform 1 0 9856 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2251_
timestamp 1698431365
transform 1 0 21616 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2252_
timestamp 1698431365
transform 1 0 21840 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2253_
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2254_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2255_
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2256_
timestamp 1698431365
transform 1 0 24528 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2257_
timestamp 1698431365
transform 1 0 24864 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2258_
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2259_
timestamp 1698431365
transform -1 0 31472 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2260_
timestamp 1698431365
transform -1 0 34160 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2261_
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2262_
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2263_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2264_
timestamp 1698431365
transform -1 0 15680 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2265_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2266_
timestamp 1698431365
transform 1 0 5936 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2267_
timestamp 1698431365
transform 1 0 5824 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2268_
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2269_
timestamp 1698431365
transform 1 0 10976 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2270_
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2271_
timestamp 1698431365
transform 1 0 12544 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2272_
timestamp 1698431365
transform 1 0 20272 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2273_
timestamp 1698431365
transform -1 0 22288 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__B1
timestamp 1698431365
transform 1 0 17584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__B1
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A3
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform 1 0 20272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A3
timestamp 1698431365
transform 1 0 29680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A4
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__I
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__I
timestamp 1698431365
transform -1 0 30912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A1
timestamp 1698431365
transform 1 0 31472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1698431365
transform -1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__I
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A1
timestamp 1698431365
transform 1 0 30128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698431365
transform -1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__I
timestamp 1698431365
transform -1 0 28672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698431365
transform 1 0 19376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698431365
transform 1 0 33376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698431365
transform -1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform -1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698431365
transform -1 0 22176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__I
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__I
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698431365
transform 1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__I
timestamp 1698431365
transform 1 0 37856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A1
timestamp 1698431365
transform 1 0 27104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__I
timestamp 1698431365
transform -1 0 34944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A2
timestamp 1698431365
transform 1 0 21728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__B
timestamp 1698431365
transform -1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform -1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__I
timestamp 1698431365
transform -1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 22512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1698431365
transform -1 0 17248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__I
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A1
timestamp 1698431365
transform 1 0 10640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__A1
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698431365
transform -1 0 21728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__I
timestamp 1698431365
transform 1 0 16240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__I
timestamp 1698431365
transform -1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__I
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__I
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__A1
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__B
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698431365
transform 1 0 8512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__A1
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A1
timestamp 1698431365
transform 1 0 31360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__A1
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A1
timestamp 1698431365
transform 1 0 37520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__I
timestamp 1698431365
transform 1 0 41776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__A1
timestamp 1698431365
transform 1 0 45360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform 1 0 37072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698431365
transform 1 0 38528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A1
timestamp 1698431365
transform -1 0 30800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A1
timestamp 1698431365
transform -1 0 34832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__I
timestamp 1698431365
transform 1 0 29120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A1
timestamp 1698431365
transform -1 0 33824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A1
timestamp 1698431365
transform -1 0 31696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A1
timestamp 1698431365
transform 1 0 33152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__I
timestamp 1698431365
transform -1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__I
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 34160 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A1
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A1
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__C
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__A2
timestamp 1698431365
transform -1 0 3584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__A2
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__B
timestamp 1698431365
transform -1 0 2352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__B
timestamp 1698431365
transform 1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__B
timestamp 1698431365
transform 1 0 3248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__B
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__I
timestamp 1698431365
transform 1 0 22400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1323__A1
timestamp 1698431365
transform 1 0 8512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__A1
timestamp 1698431365
transform -1 0 8288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__A1
timestamp 1698431365
transform -1 0 17808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__A1
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__I
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698431365
transform -1 0 18144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform -1 0 21616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform 1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698431365
transform -1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A1
timestamp 1698431365
transform 1 0 16800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform 1 0 18144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A1
timestamp 1698431365
transform -1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform -1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A1
timestamp 1698431365
transform -1 0 19936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__A1
timestamp 1698431365
transform -1 0 17584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__I
timestamp 1698431365
transform 1 0 19824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__I
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A1
timestamp 1698431365
transform 1 0 29680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__C
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A1
timestamp 1698431365
transform 1 0 7952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A2
timestamp 1698431365
transform -1 0 6832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1698431365
transform 1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform 1 0 18480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1698431365
transform 1 0 19488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A1
timestamp 1698431365
transform -1 0 28784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__A1
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1698431365
transform 1 0 44464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A1
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A1
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A1
timestamp 1698431365
transform 1 0 44912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__I
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A1
timestamp 1698431365
transform -1 0 37296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__A1
timestamp 1698431365
transform 1 0 40880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A1
timestamp 1698431365
transform 1 0 38304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform 1 0 38976 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__I
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1698431365
transform -1 0 9520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1698431365
transform -1 0 11200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A1
timestamp 1698431365
transform 1 0 31696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1698431365
transform 1 0 32144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__B
timestamp 1698431365
transform 1 0 25424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A1
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform 1 0 29792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A3
timestamp 1698431365
transform -1 0 25312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1698431365
transform -1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__B
timestamp 1698431365
transform 1 0 34160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform -1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform -1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A1
timestamp 1698431365
transform 1 0 32816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1698431365
transform 1 0 34272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 26656 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1698431365
transform 1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__I
timestamp 1698431365
transform 1 0 6496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__I
timestamp 1698431365
transform 1 0 6272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__I
timestamp 1698431365
transform -1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__B
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__B
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform -1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform -1 0 22288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1698431365
transform 1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A3
timestamp 1698431365
transform 1 0 28112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A2
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A2
timestamp 1698431365
transform -1 0 15568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform 1 0 11760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform 1 0 12544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform -1 0 14672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1698431365
transform -1 0 12656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A2
timestamp 1698431365
transform -1 0 31472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1698431365
transform 1 0 36064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__B
timestamp 1698431365
transform -1 0 31920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1698431365
transform 1 0 36624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__I
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1698431365
transform 1 0 33152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A4
timestamp 1698431365
transform -1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1698431365
transform 1 0 37856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A1
timestamp 1698431365
transform 1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1698431365
transform 1 0 31024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A2
timestamp 1698431365
transform 1 0 27216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1698431365
transform -1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A2
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__I
timestamp 1698431365
transform 1 0 30016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A1
timestamp 1698431365
transform -1 0 27216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A1
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1698431365
transform -1 0 24192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A1
timestamp 1698431365
transform 1 0 27440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1698431365
transform -1 0 23744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1698431365
transform 1 0 28784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1698431365
transform 1 0 29232 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__C
timestamp 1698431365
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1698431365
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A3
timestamp 1698431365
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__B
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1698431365
transform 1 0 33712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__B
timestamp 1698431365
transform -1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A3
timestamp 1698431365
transform 1 0 36400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1698431365
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A4
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform -1 0 29232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A2
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__B2
timestamp 1698431365
transform 1 0 28112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform -1 0 18032 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__C
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1698431365
transform -1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A3
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A2
timestamp 1698431365
transform -1 0 16576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A4
timestamp 1698431365
transform -1 0 12432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1698431365
transform -1 0 9632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1698431365
transform 1 0 9184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__B
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__B
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1698431365
transform 1 0 11984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1698431365
transform -1 0 11872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A4
timestamp 1698431365
transform -1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1698431365
transform 1 0 27328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__B
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1698431365
transform -1 0 22512 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__B
timestamp 1698431365
transform -1 0 20944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1698431365
transform -1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform 1 0 21616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__B
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__B
timestamp 1698431365
transform -1 0 28896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A1
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform -1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1698431365
transform -1 0 33264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1698431365
transform -1 0 33376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A1
timestamp 1698431365
transform 1 0 34496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1698431365
transform 1 0 33488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__B
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1698431365
transform -1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 23184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 20608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 33488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_wb_clk_i_I
timestamp 1698431365
transform -1 0 9856 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_wb_clk_i_I
timestamp 1698431365
transform 1 0 15904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_wb_clk_i_I
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_wb_clk_i_I
timestamp 1698431365
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_wb_clk_i_I
timestamp 1698431365
transform 1 0 8400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_wb_clk_i_I
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_wb_clk_i_I
timestamp 1698431365
transform 1 0 7392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_wb_clk_i_I
timestamp 1698431365
transform -1 0 15232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_wb_clk_i_I
timestamp 1698431365
transform -1 0 19376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_wb_clk_i_I
timestamp 1698431365
transform 1 0 13664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_wb_clk_i_I
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_wb_clk_i_I
timestamp 1698431365
transform 1 0 20384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_wb_clk_i_I
timestamp 1698431365
transform 1 0 31584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_wb_clk_i_I
timestamp 1698431365
transform 1 0 34720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_wb_clk_i_I
timestamp 1698431365
transform 1 0 31472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_wb_clk_i_I
timestamp 1698431365
transform -1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_wb_clk_i_I
timestamp 1698431365
transform -1 0 33264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_wb_clk_i_I
timestamp 1698431365
transform 1 0 31920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_wb_clk_i_I
timestamp 1698431365
transform 1 0 45360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_wb_clk_i_I
timestamp 1698431365
transform 1 0 44912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_wb_clk_i_I
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_wb_clk_i_I
timestamp 1698431365
transform 1 0 45360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_wb_clk_i_I
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_wb_clk_i_I
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_wb_clk_i_I
timestamp 1698431365
transform 1 0 39648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_wb_clk_i_I
timestamp 1698431365
transform 1 0 46144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_wb_clk_i_I
timestamp 1698431365
transform -1 0 27440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_wb_clk_i_I
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_wb_clk_i_I
timestamp 1698431365
transform 1 0 32928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_wb_clk_i_I
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_wb_clk_i_I
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_wb_clk_i_I
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_wb_clk_i_I
timestamp 1698431365
transform -1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_wb_clk_i_I
timestamp 1698431365
transform 1 0 14448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_wb_clk_i_I
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 46032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 34496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 23296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 31808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 38976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 41888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 45920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 45696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 41552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 15680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1698431365
transform 1 0 46032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 19824 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 33712 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 33936 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1698431365
transform -1 0 8400 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1698431365
transform 1 0 11424 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1698431365
transform 1 0 17584 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1698431365
transform 1 0 6944 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1698431365
transform -1 0 8176 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1698431365
transform -1 0 11088 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1698431365
transform -1 0 15008 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1698431365
transform 1 0 19264 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1698431365
transform 1 0 18928 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1698431365
transform -1 0 30688 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1698431365
transform -1 0 35168 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1698431365
transform -1 0 30800 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1698431365
transform -1 0 42448 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1698431365
transform -1 0 44464 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1698431365
transform -1 0 39984 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1698431365
transform -1 0 36176 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1698431365
transform -1 0 42448 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1698431365
transform -1 0 46368 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1698431365
transform -1 0 39872 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1698431365
transform -1 0 32368 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1698431365
transform -1 0 34608 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1698431365
transform -1 0 38528 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1698431365
transform 1 0 23184 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_wb_clk_i
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_wb_clk_i
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_wb_clk_i
timestamp 1698431365
transform -1 0 19936 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_wb_clk_i
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_wb_clk_i
timestamp 1698431365
transform -1 0 8736 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_12 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_17
timestamp 1698431365
transform 1 0 3248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_25
timestamp 1698431365
transform 1 0 4144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_31
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_40
timestamp 1698431365
transform 1 0 5824 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_45
timestamp 1698431365
transform 1 0 6384 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_53
timestamp 1698431365
transform 1 0 7280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133
timestamp 1698431365
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_208
timestamp 1698431365
transform 1 0 24640 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_217
timestamp 1698431365
transform 1 0 25648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698431365
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_242
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_344
timestamp 1698431365
transform 1 0 39872 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_22
timestamp 1698431365
transform 1 0 3808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_59
timestamp 1698431365
transform 1 0 7952 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698431365
transform 1 0 17472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_26
timestamp 1698431365
transform 1 0 4256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_39
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_52
timestamp 1698431365
transform 1 0 7168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_62
timestamp 1698431365
transform 1 0 8288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_109
timestamp 1698431365
transform 1 0 13552 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_136
timestamp 1698431365
transform 1 0 16576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_261
timestamp 1698431365
transform 1 0 30576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_310
timestamp 1698431365
transform 1 0 36064 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_401
timestamp 1698431365
transform 1 0 46256 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_45
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_144
timestamp 1698431365
transform 1 0 17472 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_218
timestamp 1698431365
transform 1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_291
timestamp 1698431365
transform 1 0 33936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_293
timestamp 1698431365
transform 1 0 34160 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_372
timestamp 1698431365
transform 1 0 43008 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_10
timestamp 1698431365
transform 1 0 2464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_14
timestamp 1698431365
transform 1 0 2912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_16
timestamp 1698431365
transform 1 0 3136 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_88
timestamp 1698431365
transform 1 0 11200 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_170
timestamp 1698431365
transform 1 0 20384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_187
timestamp 1698431365
transform 1 0 22288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_229
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_231
timestamp 1698431365
transform 1 0 27216 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_276
timestamp 1698431365
transform 1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_278
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_343
timestamp 1698431365
transform 1 0 39760 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_397
timestamp 1698431365
transform 1 0 45808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_401
timestamp 1698431365
transform 1 0 46256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_101
timestamp 1698431365
transform 1 0 12656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_103
timestamp 1698431365
transform 1 0 12880 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_177
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_179
timestamp 1698431365
transform 1 0 21392 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_218
timestamp 1698431365
transform 1 0 25760 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_229
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_259
timestamp 1698431365
transform 1 0 30352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_261
timestamp 1698431365
transform 1 0 30576 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_264
timestamp 1698431365
transform 1 0 30912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_327
timestamp 1698431365
transform 1 0 37968 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_6
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_33
timestamp 1698431365
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_76
timestamp 1698431365
transform 1 0 9856 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_95
timestamp 1698431365
transform 1 0 11984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_191
timestamp 1698431365
transform 1 0 22736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_193
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_196
timestamp 1698431365
transform 1 0 23296 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_200
timestamp 1698431365
transform 1 0 23744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_226
timestamp 1698431365
transform 1 0 26656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_230
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_306
timestamp 1698431365
transform 1 0 35616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_308
timestamp 1698431365
transform 1 0 35840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_328
timestamp 1698431365
transform 1 0 38080 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_401
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_6
timestamp 1698431365
transform 1 0 2016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_82
timestamp 1698431365
transform 1 0 10528 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_85
timestamp 1698431365
transform 1 0 10864 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_102
timestamp 1698431365
transform 1 0 12768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_106
timestamp 1698431365
transform 1 0 13216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_108
timestamp 1698431365
transform 1 0 13440 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_121
timestamp 1698431365
transform 1 0 14896 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_130
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_200
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_204
timestamp 1698431365
transform 1 0 24192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_222
timestamp 1698431365
transform 1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_224
timestamp 1698431365
transform 1 0 26432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_227
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_231
timestamp 1698431365
transform 1 0 27216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_235
timestamp 1698431365
transform 1 0 27664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_239
timestamp 1698431365
transform 1 0 28112 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_243
timestamp 1698431365
transform 1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_251
timestamp 1698431365
transform 1 0 29456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_255
timestamp 1698431365
transform 1 0 29904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_263
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_321
timestamp 1698431365
transform 1 0 37296 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_334
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_49
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_59
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_113
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_154
timestamp 1698431365
transform 1 0 18592 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_179
timestamp 1698431365
transform 1 0 21392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_188
timestamp 1698431365
transform 1 0 22400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_201
timestamp 1698431365
transform 1 0 23856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_232
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_276
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_280
timestamp 1698431365
transform 1 0 32704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_321
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_332
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_357
timestamp 1698431365
transform 1 0 41328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1698431365
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_393
timestamp 1698431365
transform 1 0 45360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_4
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_40
timestamp 1698431365
transform 1 0 5824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_52
timestamp 1698431365
transform 1 0 7168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_62
timestamp 1698431365
transform 1 0 8288 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_327
timestamp 1698431365
transform 1 0 37968 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_333
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_354
timestamp 1698431365
transform 1 0 40992 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_371
timestamp 1698431365
transform 1 0 42896 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_112
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_116
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_118
timestamp 1698431365
transform 1 0 14560 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_135
timestamp 1698431365
transform 1 0 16464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_142
timestamp 1698431365
transform 1 0 17248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_150
timestamp 1698431365
transform 1 0 18144 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_187
timestamp 1698431365
transform 1 0 22288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_190
timestamp 1698431365
transform 1 0 22624 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_198
timestamp 1698431365
transform 1 0 23520 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_230
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_297
timestamp 1698431365
transform 1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_299
timestamp 1698431365
transform 1 0 34832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_304
timestamp 1698431365
transform 1 0 35392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_306
timestamp 1698431365
transform 1 0 35616 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_348
timestamp 1698431365
transform 1 0 40320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_374
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_393
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_31
timestamp 1698431365
transform 1 0 4816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_35
timestamp 1698431365
transform 1 0 5264 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_58
timestamp 1698431365
transform 1 0 7840 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_94
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_98
timestamp 1698431365
transform 1 0 12320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_173
timestamp 1698431365
transform 1 0 20720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_233
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_239
timestamp 1698431365
transform 1 0 28112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_263
timestamp 1698431365
transform 1 0 30800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_267
timestamp 1698431365
transform 1 0 31248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_271
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_291
timestamp 1698431365
transform 1 0 33936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_293
timestamp 1698431365
transform 1 0 34160 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_331
timestamp 1698431365
transform 1 0 38416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_333
timestamp 1698431365
transform 1 0 38640 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_364
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_10
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_117
timestamp 1698431365
transform 1 0 14448 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_125
timestamp 1698431365
transform 1 0 15344 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_129
timestamp 1698431365
transform 1 0 15792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_281
timestamp 1698431365
transform 1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_283
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_341
timestamp 1698431365
transform 1 0 39536 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_361
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_45
timestamp 1698431365
transform 1 0 6384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_57
timestamp 1698431365
transform 1 0 7728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_61
timestamp 1698431365
transform 1 0 8176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_63
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_116
timestamp 1698431365
transform 1 0 14336 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_130
timestamp 1698431365
transform 1 0 15904 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698431365
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_154
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_271
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_354
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_10
timestamp 1698431365
transform 1 0 2464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_14
timestamp 1698431365
transform 1 0 2912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_29
timestamp 1698431365
transform 1 0 4592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_33
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_92
timestamp 1698431365
transform 1 0 11648 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_115
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_117
timestamp 1698431365
transform 1 0 14448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_161
timestamp 1698431365
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_163
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_183
timestamp 1698431365
transform 1 0 21840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_233
timestamp 1698431365
transform 1 0 27440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_252
timestamp 1698431365
transform 1 0 29568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_266
timestamp 1698431365
transform 1 0 31136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_358
timestamp 1698431365
transform 1 0 41440 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_364
timestamp 1698431365
transform 1 0 42112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_366
timestamp 1698431365
transform 1 0 42336 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_375
timestamp 1698431365
transform 1 0 43344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_399
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_401
timestamp 1698431365
transform 1 0 46256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_39
timestamp 1698431365
transform 1 0 5712 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_85
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_135
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_153
timestamp 1698431365
transform 1 0 18480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_187
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_191
timestamp 1698431365
transform 1 0 22736 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698431365
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698431365
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_230
timestamp 1698431365
transform 1 0 27104 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_245
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_340
timestamp 1698431365
transform 1 0 39424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_61
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_63
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_86
timestamp 1698431365
transform 1 0 10976 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_140
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_142
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_198
timestamp 1698431365
transform 1 0 23520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_239
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_249
timestamp 1698431365
transform 1 0 29232 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_269
timestamp 1698431365
transform 1 0 31472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_293
timestamp 1698431365
transform 1 0 34160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_295
timestamp 1698431365
transform 1 0 34384 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_395
timestamp 1698431365
transform 1 0 45584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_399
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_401
timestamp 1698431365
transform 1 0 46256 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_39
timestamp 1698431365
transform 1 0 5712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_109
timestamp 1698431365
transform 1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_168
timestamp 1698431365
transform 1 0 20160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_226
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_233
timestamp 1698431365
transform 1 0 27440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_237
timestamp 1698431365
transform 1 0 27888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_325
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_327
timestamp 1698431365
transform 1 0 37968 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_347
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_363
timestamp 1698431365
transform 1 0 42000 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_16
timestamp 1698431365
transform 1 0 3136 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_20
timestamp 1698431365
transform 1 0 3584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_44
timestamp 1698431365
transform 1 0 6272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_48
timestamp 1698431365
transform 1 0 6720 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_64
timestamp 1698431365
transform 1 0 8512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_72
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_169
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_198
timestamp 1698431365
transform 1 0 23520 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_239
timestamp 1698431365
transform 1 0 28112 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_265
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_267
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_380
timestamp 1698431365
transform 1 0 43904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_391
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_395
timestamp 1698431365
transform 1 0 45584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_31
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_33
timestamp 1698431365
transform 1 0 5040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698431365
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_90
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_92
timestamp 1698431365
transform 1 0 11648 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_128
timestamp 1698431365
transform 1 0 15680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_148
timestamp 1698431365
transform 1 0 17920 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_176
timestamp 1698431365
transform 1 0 21056 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_218
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_260
timestamp 1698431365
transform 1 0 30464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_264
timestamp 1698431365
transform 1 0 30912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_266
timestamp 1698431365
transform 1 0 31136 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_339
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_398
timestamp 1698431365
transform 1 0 45920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_31
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_50
timestamp 1698431365
transform 1 0 6944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_67
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_71
timestamp 1698431365
transform 1 0 9296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698431365
transform 1 0 9744 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_129
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_168
timestamp 1698431365
transform 1 0 20160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_190
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_283
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_285
timestamp 1698431365
transform 1 0 33264 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_322
timestamp 1698431365
transform 1 0 37408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_324
timestamp 1698431365
transform 1 0 37632 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_340
timestamp 1698431365
transform 1 0 39424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_401
timestamp 1698431365
transform 1 0 46256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_4
timestamp 1698431365
transform 1 0 1792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_76
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_162
timestamp 1698431365
transform 1 0 19488 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_166
timestamp 1698431365
transform 1 0 19936 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_202
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_238
timestamp 1698431365
transform 1 0 28000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_242
timestamp 1698431365
transform 1 0 28448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_246
timestamp 1698431365
transform 1 0 28896 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_250
timestamp 1698431365
transform 1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_258
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_269
timestamp 1698431365
transform 1 0 31472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_308
timestamp 1698431365
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_312
timestamp 1698431365
transform 1 0 36288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_317
timestamp 1698431365
transform 1 0 36848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_321
timestamp 1698431365
transform 1 0 37296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_74
timestamp 1698431365
transform 1 0 9632 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_82
timestamp 1698431365
transform 1 0 10528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_90
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_94
timestamp 1698431365
transform 1 0 11872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_96
timestamp 1698431365
transform 1 0 12096 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_111
timestamp 1698431365
transform 1 0 13776 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_120
timestamp 1698431365
transform 1 0 14784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_122
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698431365
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_164
timestamp 1698431365
transform 1 0 19712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_167
timestamp 1698431365
transform 1 0 20048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_187
timestamp 1698431365
transform 1 0 22288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_265
timestamp 1698431365
transform 1 0 31024 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_295
timestamp 1698431365
transform 1 0 34384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_299
timestamp 1698431365
transform 1 0 34832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_308
timestamp 1698431365
transform 1 0 35840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_310
timestamp 1698431365
transform 1 0 36064 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_401
timestamp 1698431365
transform 1 0 46256 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_44
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_53
timestamp 1698431365
transform 1 0 7280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_55
timestamp 1698431365
transform 1 0 7504 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_96
timestamp 1698431365
transform 1 0 12096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_127
timestamp 1698431365
transform 1 0 15568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_129
timestamp 1698431365
transform 1 0 15792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_148
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_187
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_218
timestamp 1698431365
transform 1 0 25760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_286
timestamp 1698431365
transform 1 0 33376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_288
timestamp 1698431365
transform 1 0 33600 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_291
timestamp 1698431365
transform 1 0 33936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_354
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_371
timestamp 1698431365
transform 1 0 42896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_10
timestamp 1698431365
transform 1 0 2464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_16
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_42
timestamp 1698431365
transform 1 0 6048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_46
timestamp 1698431365
transform 1 0 6496 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_146
timestamp 1698431365
transform 1 0 17696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_240
timestamp 1698431365
transform 1 0 28224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_254
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_258
timestamp 1698431365
transform 1 0 30240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_260
timestamp 1698431365
transform 1 0 30464 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_333
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_349
timestamp 1698431365
transform 1 0 40432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_351
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_356
timestamp 1698431365
transform 1 0 41216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_393
timestamp 1698431365
transform 1 0 45360 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_42
timestamp 1698431365
transform 1 0 6048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_85
timestamp 1698431365
transform 1 0 10864 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_101
timestamp 1698431365
transform 1 0 12656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_214
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_241
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_249
timestamp 1698431365
transform 1 0 29232 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_284
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_311
timestamp 1698431365
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_319
timestamp 1698431365
transform 1 0 37072 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_323
timestamp 1698431365
transform 1 0 37520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_325
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_361
timestamp 1698431365
transform 1 0 41776 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_61
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_63
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_93
timestamp 1698431365
transform 1 0 11760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_109
timestamp 1698431365
transform 1 0 13552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_124
timestamp 1698431365
transform 1 0 15232 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_155
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_161
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_163
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_182
timestamp 1698431365
transform 1 0 21728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_191
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_333
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_337
timestamp 1698431365
transform 1 0 39088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_351
timestamp 1698431365
transform 1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_355
timestamp 1698431365
transform 1 0 41104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_359
timestamp 1698431365
transform 1 0 41552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_393
timestamp 1698431365
transform 1 0 45360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_395
timestamp 1698431365
transform 1 0 45584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_39
timestamp 1698431365
transform 1 0 5712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_41
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_56
timestamp 1698431365
transform 1 0 7616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_114
timestamp 1698431365
transform 1 0 14112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_116
timestamp 1698431365
transform 1 0 14336 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_125
timestamp 1698431365
transform 1 0 15344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_218
timestamp 1698431365
transform 1 0 25760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_250
timestamp 1698431365
transform 1 0 29344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_310
timestamp 1698431365
transform 1 0 36064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_312
timestamp 1698431365
transform 1 0 36288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_332
timestamp 1698431365
transform 1 0 38528 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_138
timestamp 1698431365
transform 1 0 16800 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_142
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_146
timestamp 1698431365
transform 1 0 17696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_163
timestamp 1698431365
transform 1 0 19600 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_225
timestamp 1698431365
transform 1 0 26544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_233
timestamp 1698431365
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_259
timestamp 1698431365
transform 1 0 30352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_282
timestamp 1698431365
transform 1 0 32928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_286
timestamp 1698431365
transform 1 0 33376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_290
timestamp 1698431365
transform 1 0 33824 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_298
timestamp 1698431365
transform 1 0 34720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_326
timestamp 1698431365
transform 1 0 37856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_340
timestamp 1698431365
transform 1 0 39424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_354
timestamp 1698431365
transform 1 0 40992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_367
timestamp 1698431365
transform 1 0 42448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_393
timestamp 1698431365
transform 1 0 45360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_397
timestamp 1698431365
transform 1 0 45808 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_32
timestamp 1698431365
transform 1 0 4928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_78
timestamp 1698431365
transform 1 0 10080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_201
timestamp 1698431365
transform 1 0 23856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_245
timestamp 1698431365
transform 1 0 28784 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_249
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_284
timestamp 1698431365
transform 1 0 33152 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_319
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_336
timestamp 1698431365
transform 1 0 38976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_342
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_47
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_54
timestamp 1698431365
transform 1 0 7392 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_206
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_268
timestamp 1698431365
transform 1 0 31360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_272
timestamp 1698431365
transform 1 0 31808 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_276
timestamp 1698431365
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_280
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_282
timestamp 1698431365
transform 1 0 32928 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_291
timestamp 1698431365
transform 1 0 33936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_295
timestamp 1698431365
transform 1 0 34384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_297
timestamp 1698431365
transform 1 0 34608 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_306
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_324
timestamp 1698431365
transform 1 0 37632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_328
timestamp 1698431365
transform 1 0 38080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_330
timestamp 1698431365
transform 1 0 38304 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_365
timestamp 1698431365
transform 1 0 42224 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_10
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_47
timestamp 1698431365
transform 1 0 6608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_49
timestamp 1698431365
transform 1 0 6832 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698431365
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_92
timestamp 1698431365
transform 1 0 11648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_160
timestamp 1698431365
transform 1 0 19264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_201
timestamp 1698431365
transform 1 0 23856 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_214
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_268
timestamp 1698431365
transform 1 0 31360 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_337
timestamp 1698431365
transform 1 0 39088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_358
timestamp 1698431365
transform 1 0 41440 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_371
timestamp 1698431365
transform 1 0 42896 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_31
timestamp 1698431365
transform 1 0 4816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_98
timestamp 1698431365
transform 1 0 12320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_113
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_212
timestamp 1698431365
transform 1 0 25088 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_233
timestamp 1698431365
transform 1 0 27440 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_282
timestamp 1698431365
transform 1 0 32928 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_346
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_395
timestamp 1698431365
transform 1 0 45584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_399
timestamp 1698431365
transform 1 0 46032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_48
timestamp 1698431365
transform 1 0 6720 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_112
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_133
timestamp 1698431365
transform 1 0 16240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_151
timestamp 1698431365
transform 1 0 18256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_184
timestamp 1698431365
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_90
timestamp 1698431365
transform 1 0 11424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_92
timestamp 1698431365
transform 1 0 11648 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_97
timestamp 1698431365
transform 1 0 12208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_203
timestamp 1698431365
transform 1 0 24080 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_205
timestamp 1698431365
transform 1 0 24304 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_220
timestamp 1698431365
transform 1 0 25984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_249
timestamp 1698431365
transform 1 0 29232 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_254
timestamp 1698431365
transform 1 0 29792 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_265
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_274
timestamp 1698431365
transform 1 0 32032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_284
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_296
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_10
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_78
timestamp 1698431365
transform 1 0 10080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_109
timestamp 1698431365
transform 1 0 13552 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_171
timestamp 1698431365
transform 1 0 20496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_383
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_387
timestamp 1698431365
transform 1 0 44688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_391
timestamp 1698431365
transform 1 0 45136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_395
timestamp 1698431365
transform 1 0 45584 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_400
timestamp 1698431365
transform 1 0 46144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_31
timestamp 1698431365
transform 1 0 4816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_42
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_94
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_122
timestamp 1698431365
transform 1 0 15008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_124
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_131
timestamp 1698431365
transform 1 0 16016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_135
timestamp 1698431365
transform 1 0 16464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_137
timestamp 1698431365
transform 1 0 16688 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_140
timestamp 1698431365
transform 1 0 17024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_144
timestamp 1698431365
transform 1 0 17472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_148
timestamp 1698431365
transform 1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_156
timestamp 1698431365
transform 1 0 18816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_160
timestamp 1698431365
transform 1 0 19264 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_235
timestamp 1698431365
transform 1 0 27664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_237
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_257
timestamp 1698431365
transform 1 0 30128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_301
timestamp 1698431365
transform 1 0 35056 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_303
timestamp 1698431365
transform 1 0 35280 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_335
timestamp 1698431365
transform 1 0 38864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_400
timestamp 1698431365
transform 1 0 46144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_50
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_122
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_130
timestamp 1698431365
transform 1 0 15904 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_228
timestamp 1698431365
transform 1 0 26880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_238
timestamp 1698431365
transform 1 0 28000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_242
timestamp 1698431365
transform 1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_246
timestamp 1698431365
transform 1 0 28896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_250
timestamp 1698431365
transform 1 0 29344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_262
timestamp 1698431365
transform 1 0 30688 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_269
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_341
timestamp 1698431365
transform 1 0 39536 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_345
timestamp 1698431365
transform 1 0 39984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_31
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_66
timestamp 1698431365
transform 1 0 8736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_70
timestamp 1698431365
transform 1 0 9184 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_83
timestamp 1698431365
transform 1 0 10640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_85
timestamp 1698431365
transform 1 0 10864 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_88
timestamp 1698431365
transform 1 0 11200 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_92
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_95
timestamp 1698431365
transform 1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_99
timestamp 1698431365
transform 1 0 12432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_165
timestamp 1698431365
transform 1 0 19824 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_179
timestamp 1698431365
transform 1 0 21392 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_186
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_249
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_271
timestamp 1698431365
transform 1 0 31696 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_19
timestamp 1698431365
transform 1 0 3472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_21
timestamp 1698431365
transform 1 0 3696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_38
timestamp 1698431365
transform 1 0 5600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_64
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_84
timestamp 1698431365
transform 1 0 10752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_98
timestamp 1698431365
transform 1 0 12320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_102
timestamp 1698431365
transform 1 0 12768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_115
timestamp 1698431365
transform 1 0 14224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_119
timestamp 1698431365
transform 1 0 14672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_123
timestamp 1698431365
transform 1 0 15120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_125
timestamp 1698431365
transform 1 0 15344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_132
timestamp 1698431365
transform 1 0 16128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_146
timestamp 1698431365
transform 1 0 17696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_151
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_153
timestamp 1698431365
transform 1 0 18480 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_161
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_165
timestamp 1698431365
transform 1 0 19824 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_168
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_185
timestamp 1698431365
transform 1 0 22064 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_217
timestamp 1698431365
transform 1 0 25648 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_226
timestamp 1698431365
transform 1 0 26656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_230
timestamp 1698431365
transform 1 0 27104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_234
timestamp 1698431365
transform 1 0 27552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_238
timestamp 1698431365
transform 1 0 28000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_10
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_49
timestamp 1698431365
transform 1 0 6832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_102
timestamp 1698431365
transform 1 0 12768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_302
timestamp 1698431365
transform 1 0 35168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_328
timestamp 1698431365
transform 1 0 38080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_31
timestamp 1698431365
transform 1 0 4816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_122
timestamp 1698431365
transform 1 0 15008 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_131
timestamp 1698431365
transform 1 0 16016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_133
timestamp 1698431365
transform 1 0 16240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_155
timestamp 1698431365
transform 1 0 18704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_270
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_311
timestamp 1698431365
transform 1 0 36176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_357
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_10
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_25
timestamp 1698431365
transform 1 0 4144 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_185
timestamp 1698431365
transform 1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_202
timestamp 1698431365
transform 1 0 23968 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_208
timestamp 1698431365
transform 1 0 24640 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_242
timestamp 1698431365
transform 1 0 28448 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_260
timestamp 1698431365
transform 1 0 30464 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_290
timestamp 1698431365
transform 1 0 33824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_292
timestamp 1698431365
transform 1 0 34048 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_307
timestamp 1698431365
transform 1 0 35728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_368
timestamp 1698431365
transform 1 0 42560 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_86
timestamp 1698431365
transform 1 0 10976 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_88
timestamp 1698431365
transform 1 0 11200 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_105
timestamp 1698431365
transform 1 0 13104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_155
timestamp 1698431365
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_157
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_187
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_194
timestamp 1698431365
transform 1 0 23072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_214
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_217
timestamp 1698431365
transform 1 0 25648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_219
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_265
timestamp 1698431365
transform 1 0 31024 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_274
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_300
timestamp 1698431365
transform 1 0 34944 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_10
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698431365
transform 1 0 24864 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_281
timestamp 1698431365
transform 1 0 32816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_285
timestamp 1698431365
transform 1 0 33264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_289
timestamp 1698431365
transform 1 0 33712 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_10
timestamp 1698431365
transform 1 0 2464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_28
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698431365
transform 1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_63
timestamp 1698431365
transform 1 0 8400 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_119
timestamp 1698431365
transform 1 0 14672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_121
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_200
timestamp 1698431365
transform 1 0 23744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_252
timestamp 1698431365
transform 1 0 29568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_256
timestamp 1698431365
transform 1 0 30016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_258
timestamp 1698431365
transform 1 0 30240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_269
timestamp 1698431365
transform 1 0 31472 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_273
timestamp 1698431365
transform 1 0 31920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_277
timestamp 1698431365
transform 1 0 32368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_303
timestamp 1698431365
transform 1 0 35280 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_305
timestamp 1698431365
transform 1 0 35504 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_385
timestamp 1698431365
transform 1 0 44464 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_31
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_45
timestamp 1698431365
transform 1 0 6384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_49
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_52
timestamp 1698431365
transform 1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_69
timestamp 1698431365
transform 1 0 9072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_84
timestamp 1698431365
transform 1 0 10752 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_97
timestamp 1698431365
transform 1 0 12208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_249
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_274
timestamp 1698431365
transform 1 0 32032 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_393
timestamp 1698431365
transform 1 0 45360 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_38
timestamp 1698431365
transform 1 0 5600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_40
timestamp 1698431365
transform 1 0 5824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_85
timestamp 1698431365
transform 1 0 10864 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_288
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_292
timestamp 1698431365
transform 1 0 34048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_296
timestamp 1698431365
transform 1 0 34496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_310
timestamp 1698431365
transform 1 0 36064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_312
timestamp 1698431365
transform 1 0 36288 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_331
timestamp 1698431365
transform 1 0 38416 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_401
timestamp 1698431365
transform 1 0 46256 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_53
timestamp 1698431365
transform 1 0 7280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_61
timestamp 1698431365
transform 1 0 8176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_65
timestamp 1698431365
transform 1 0 8624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_67
timestamp 1698431365
transform 1 0 8848 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_109
timestamp 1698431365
transform 1 0 13552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_210
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_279
timestamp 1698431365
transform 1 0 32592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_291
timestamp 1698431365
transform 1 0 33936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_295
timestamp 1698431365
transform 1 0 34384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_297
timestamp 1698431365
transform 1 0 34608 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_308
timestamp 1698431365
transform 1 0 35840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_383
timestamp 1698431365
transform 1 0 44240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_401
timestamp 1698431365
transform 1 0 46256 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_38
timestamp 1698431365
transform 1 0 5600 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_122
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_159
timestamp 1698431365
transform 1 0 19152 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_96
timestamp 1698431365
transform 1 0 12096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_98
timestamp 1698431365
transform 1 0 12320 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_117
timestamp 1698431365
transform 1 0 14448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_229
timestamp 1698431365
transform 1 0 26992 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_233
timestamp 1698431365
transform 1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_237
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_267
timestamp 1698431365
transform 1 0 31248 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_271
timestamp 1698431365
transform 1 0 31696 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_289
timestamp 1698431365
transform 1 0 33712 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_293
timestamp 1698431365
transform 1 0 34160 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_401
timestamp 1698431365
transform 1 0 46256 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_34
timestamp 1698431365
transform 1 0 5152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_38
timestamp 1698431365
transform 1 0 5600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_80
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_245
timestamp 1698431365
transform 1 0 28784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_275
timestamp 1698431365
transform 1 0 32144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_370
timestamp 1698431365
transform 1 0 42784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_372
timestamp 1698431365
transform 1 0 43008 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_36
timestamp 1698431365
transform 1 0 5376 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_70
timestamp 1698431365
transform 1 0 9184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_80
timestamp 1698431365
transform 1 0 10304 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_96
timestamp 1698431365
transform 1 0 12096 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_106
timestamp 1698431365
transform 1 0 13216 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_120
timestamp 1698431365
transform 1 0 14784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_124
timestamp 1698431365
transform 1 0 15232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_134
timestamp 1698431365
transform 1 0 16352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_138
timestamp 1698431365
transform 1 0 16800 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_145
timestamp 1698431365
transform 1 0 17584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_157
timestamp 1698431365
transform 1 0 18928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_161
timestamp 1698431365
transform 1 0 19376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_201
timestamp 1698431365
transform 1 0 23856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_203
timestamp 1698431365
transform 1 0 24080 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_206
timestamp 1698431365
transform 1 0 24416 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_208
timestamp 1698431365
transform 1 0 24640 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_240
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_242
timestamp 1698431365
transform 1 0 28448 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_245
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_269
timestamp 1698431365
transform 1 0 31472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_271
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_280
timestamp 1698431365
transform 1 0 32704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_282
timestamp 1698431365
transform 1 0 32928 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_308
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_310
timestamp 1698431365
transform 1 0 36064 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_342
timestamp 1698431365
transform 1 0 39648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_344
timestamp 1698431365
transform 1 0 39872 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_400
timestamp 1698431365
transform 1 0 46144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 46368 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 39872 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 46368 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 46368 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform -1 0 46368 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 46368 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 46368 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform -1 0 46368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 46368 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 46368 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698431365
transform -1 0 46144 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input13
timestamp 1698431365
transform 1 0 18032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 32592 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform -1 0 39760 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform -1 0 16576 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_53 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 46592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_54
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 46592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_55
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 46592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 46592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 46592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 46592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 46592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 46592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 46592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 46592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 46592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 46592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 46592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 46592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 46592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 46592 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 46592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 46592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 46592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 46592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 46592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 46592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 46592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 46592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 46592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 46592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 46592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 46592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 46592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 46592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 46592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 46592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 46592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 46592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 46592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 46592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 46592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 46592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 46592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 46592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 46592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 46592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 46592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 46592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 46592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 46592 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 46592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 46592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 46592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_117
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_118
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_119
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_120
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_121
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_122
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_123
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_124
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_125
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_126
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_128
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_129
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_130
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_131
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_132
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_133
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_134
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_135
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_136
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_137
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_139
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_140
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_141
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_142
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_143
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_144
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_145
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_146
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_147
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_148
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_150
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_151
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_152
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_153
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_154
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_155
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_156
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_157
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_158
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_159
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_161
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_162
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_163
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_164
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_165
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_166
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_167
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_168
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_169
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_170
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_172
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_173
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_174
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_175
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_176
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_177
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_178
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_179
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_180
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_181
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_183
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_184
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_191
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_192
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_194
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_195
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_196
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_197
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_198
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_199
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_200
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_201
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_202
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_203
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_205
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_206
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_207
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_208
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_209
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_210
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_211
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_212
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_213
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_214
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_216
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_217
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_218
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_219
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_220
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_221
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_222
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_223
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_224
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_225
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_227
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_228
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_229
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_230
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_231
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_232
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_233
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_234
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_235
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_236
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_238
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_239
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_240
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_241
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_242
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_243
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_244
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_245
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_246
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_247
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_249
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_250
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_251
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_252
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_253
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_254
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_255
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_256
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_257
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_258
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_260
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_261
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_262
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_263
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_264
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_265
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_266
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_267
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_268
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_269
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_271
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_272
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_273
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_274
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_275
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_276
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_277
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_278
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_279
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_280
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_282
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_283
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_284
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_285
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_286
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_287
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_288
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_289
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_290
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_291
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_293
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_294
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_295
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_296
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_297
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_298
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_299
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_300
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_301
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_302
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_304
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_305
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_306
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_307
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_308
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_309
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_310
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_311
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_312
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_313
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_315
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_316
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_317
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_318
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_319
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_320
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_321
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_322
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_323
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_324
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_326
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_327
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_328
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_329
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_330
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_331
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_332
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_333
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_334
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_335
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_337
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_338
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_339
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_340
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_341
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_342
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_343
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_344
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_345
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_346
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_348
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_349
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_350
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_351
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_352
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_353
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_354
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_355
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_356
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_357
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_359
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_360
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_361
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_362
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_363
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_364
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_365
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_366
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_367
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_368
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_370
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_371
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_372
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_373
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_374
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_375
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_376
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_377
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_378
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_379
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_381
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_382
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_383
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_384
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_385
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_386
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_387
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_388
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_389
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_390
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_392
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_393
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_394
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_395
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_396
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_397
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_398
timestamp 1698431365
transform 1 0 8960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_399
timestamp 1698431365
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_400
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_401
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 24192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 31808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 43232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_23 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_24
timestamp 1698431365
transform -1 0 4816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_25
timestamp 1698431365
transform -1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_26
timestamp 1698431365
transform -1 0 7840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_27
timestamp 1698431365
transform 1 0 7840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_28
timestamp 1698431365
transform 1 0 8736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_29
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_30
timestamp 1698431365
transform 1 0 11312 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_31
timestamp 1698431365
transform -1 0 24752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_32
timestamp 1698431365
transform -1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_33
timestamp 1698431365
transform -1 0 25200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_34
timestamp 1698431365
transform -1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_35
timestamp 1698431365
transform 1 0 25760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_36
timestamp 1698431365
transform -1 0 42672 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_37
timestamp 1698431365
transform -1 0 43120 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_38
timestamp 1698431365
transform -1 0 46032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_39
timestamp 1698431365
transform -1 0 45136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_40
timestamp 1698431365
transform -1 0 45584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_ay8913_41
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 534 870
<< labels >>
flabel metal3 s 47200 40320 48000 40432 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 47200 45024 48000 45136 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 47200 2688 48000 2800 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 47200 7392 48000 7504 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 47200 12096 48000 12208 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 47200 16800 48000 16912 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 47200 21504 48000 21616 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 47200 26208 48000 26320 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 47200 30912 48000 31024 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 47200 35616 48000 35728 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal2 s 29792 47200 29904 48000 0 FreeSans 448 90 0 0 io_in_2[0]
port 10 nsew signal input
flabel metal2 s 41664 47200 41776 48000 0 FreeSans 448 90 0 0 io_in_2[1]
port 11 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 24640 0 24752 800 0 FreeSans 448 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 4256 0 4368 800 0 FreeSans 448 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 io_out[27]
port 31 nsew signal tristate
flabel metal2 s 5824 0 5936 800 0 FreeSans 448 90 0 0 io_out[2]
port 32 nsew signal tristate
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 io_out[3]
port 33 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 io_out[4]
port 34 nsew signal tristate
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 io_out[5]
port 35 nsew signal tristate
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 io_out[6]
port 36 nsew signal tristate
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 io_out[7]
port 37 nsew signal tristate
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 io_out[8]
port 38 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 io_out[9]
port 39 nsew signal tristate
flabel metal2 s 17920 47200 18032 48000 0 FreeSans 448 90 0 0 rst_n
port 40 nsew signal input
flabel metal4 s 4448 3076 4768 44748 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 35168 3076 35488 44748 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 19808 3076 20128 44748 0 FreeSans 1280 90 0 0 vss
port 42 nsew ground bidirectional
flabel metal2 s 6048 47200 6160 48000 0 FreeSans 448 90 0 0 wb_clk_i
port 43 nsew signal input
rlabel metal1 23968 44688 23968 44688 0 vdd
rlabel metal1 23968 43904 23968 43904 0 vss
rlabel metal2 30632 16520 30632 16520 0 _0000_
rlabel metal2 31416 15148 31416 15148 0 _0001_
rlabel metal3 30632 12824 30632 12824 0 _0002_
rlabel metal2 30632 11144 30632 11144 0 _0003_
rlabel metal2 27832 18088 27832 18088 0 _0004_
rlabel metal2 31640 8568 31640 8568 0 _0005_
rlabel metal2 32312 4760 32312 4760 0 _0006_
rlabel metal3 36456 4424 36456 4424 0 _0007_
rlabel metal3 39256 7168 39256 7168 0 _0008_
rlabel metal2 20552 31976 20552 31976 0 _0009_
rlabel metal2 23016 34552 23016 34552 0 _0010_
rlabel metal2 21448 34552 21448 34552 0 _0011_
rlabel metal2 21392 36568 21392 36568 0 _0012_
rlabel metal2 22904 17640 22904 17640 0 _0013_
rlabel metal3 19376 15176 19376 15176 0 _0014_
rlabel metal2 19096 10752 19096 10752 0 _0015_
rlabel metal3 17472 12376 17472 12376 0 _0016_
rlabel metal2 15624 10192 15624 10192 0 _0017_
rlabel metal2 12600 11088 12600 11088 0 _0018_
rlabel metal2 9464 10192 9464 10192 0 _0019_
rlabel metal2 10360 7784 10360 7784 0 _0020_
rlabel metal2 14000 7560 14000 7560 0 _0021_
rlabel metal2 22120 6272 22120 6272 0 _0022_
rlabel metal2 22680 8008 22680 8008 0 _0023_
rlabel metal2 16520 8120 16520 8120 0 _0024_
rlabel metal2 17080 7224 17080 7224 0 _0025_
rlabel metal2 19096 6216 19096 6216 0 _0026_
rlabel metal2 10808 5992 10808 5992 0 _0027_
rlabel metal2 10864 4424 10864 4424 0 _0028_
rlabel metal3 9576 3416 9576 3416 0 _0029_
rlabel metal2 14728 4816 14728 4816 0 _0030_
rlabel metal3 16072 4200 16072 4200 0 _0031_
rlabel metal2 16128 20664 16128 20664 0 _0032_
rlabel metal2 14952 16520 14952 16520 0 _0033_
rlabel metal2 2520 16520 2520 16520 0 _0034_
rlabel metal2 5320 10640 5320 10640 0 _0035_
rlabel metal2 2856 10920 2856 10920 0 _0036_
rlabel metal2 8120 10976 8120 10976 0 _0037_
rlabel metal2 6440 8624 6440 8624 0 _0038_
rlabel metal2 13944 4088 13944 4088 0 _0039_
rlabel metal2 30520 9464 30520 9464 0 _0040_
rlabel metal2 33880 10920 33880 10920 0 _0041_
rlabel metal2 35448 9968 35448 9968 0 _0042_
rlabel metal2 34552 7784 34552 7784 0 _0043_
rlabel metal2 38248 16576 38248 16576 0 _0044_
rlabel metal2 41496 16352 41496 16352 0 _0045_
rlabel metal2 45472 15848 45472 15848 0 _0046_
rlabel metal2 45136 15848 45136 15848 0 _0047_
rlabel metal2 32088 20832 32088 20832 0 _0048_
rlabel metal2 30800 19320 30800 19320 0 _0049_
rlabel metal2 35448 17416 35448 17416 0 _0050_
rlabel metal2 35672 19488 35672 19488 0 _0051_
rlabel metal3 33600 27272 33600 27272 0 _0052_
rlabel metal2 30408 25088 30408 25088 0 _0053_
rlabel metal2 31080 26600 31080 26600 0 _0054_
rlabel metal2 35448 28728 35448 28728 0 _0055_
rlabel metal2 38360 30464 38360 30464 0 _0056_
rlabel metal3 44184 28616 44184 28616 0 _0057_
rlabel metal2 44072 31304 44072 31304 0 _0058_
rlabel metal2 41552 30296 41552 30296 0 _0059_
rlabel metal2 26040 4816 26040 4816 0 _0060_
rlabel metal2 25144 9016 25144 9016 0 _0061_
rlabel metal2 24696 7000 24696 7000 0 _0062_
rlabel metal3 30856 5320 30856 5320 0 _0063_
rlabel metal2 28056 7952 28056 7952 0 _0064_
rlabel metal2 3192 14952 3192 14952 0 _0065_
rlabel metal2 2968 13384 2968 13384 0 _0066_
rlabel metal2 2632 9296 2632 9296 0 _0067_
rlabel metal3 4480 7336 4480 7336 0 _0068_
rlabel metal2 2520 6440 2520 6440 0 _0069_
rlabel metal2 6440 7056 6440 7056 0 _0070_
rlabel metal3 6944 4200 6944 4200 0 _0071_
rlabel metal2 8568 6328 8568 6328 0 _0072_
rlabel metal2 23016 26544 23016 26544 0 _0073_
rlabel metal2 20440 25872 20440 25872 0 _0074_
rlabel metal2 15736 31304 15736 31304 0 _0075_
rlabel metal2 15400 32984 15400 32984 0 _0076_
rlabel metal3 17752 33432 17752 33432 0 _0077_
rlabel metal2 19544 31248 19544 31248 0 _0078_
rlabel metal2 21448 40432 21448 40432 0 _0079_
rlabel metal2 25368 42336 25368 42336 0 _0080_
rlabel metal2 23688 43876 23688 43876 0 _0081_
rlabel metal2 19600 44408 19600 44408 0 _0082_
rlabel metal2 31640 4256 31640 4256 0 _0083_
rlabel metal2 21896 4424 21896 4424 0 _0084_
rlabel metal2 29512 4256 29512 4256 0 _0085_
rlabel metal2 5992 14756 5992 14756 0 _0086_
rlabel metal2 16296 27384 16296 27384 0 _0087_
rlabel metal2 16408 24248 16408 24248 0 _0088_
rlabel metal3 23296 24920 23296 24920 0 _0089_
rlabel metal3 16296 27944 16296 27944 0 _0090_
rlabel metal2 28392 24864 28392 24864 0 _0091_
rlabel metal2 23184 22456 23184 22456 0 _0092_
rlabel metal2 35672 32144 35672 32144 0 _0093_
rlabel metal2 37352 34496 37352 34496 0 _0094_
rlabel metal2 35896 36064 35896 36064 0 _0095_
rlabel metal2 38248 34888 38248 34888 0 _0096_
rlabel metal3 38808 31640 38808 31640 0 _0097_
rlabel metal2 43512 34496 43512 34496 0 _0098_
rlabel metal2 44968 34048 44968 34048 0 _0099_
rlabel metal2 44576 42504 44576 42504 0 _0100_
rlabel metal2 12040 34384 12040 34384 0 _0101_
rlabel metal2 2520 33488 2520 33488 0 _0102_
rlabel metal2 2520 36064 2520 36064 0 _0103_
rlabel metal2 2744 39088 2744 39088 0 _0104_
rlabel metal2 3864 36848 3864 36848 0 _0105_
rlabel metal2 5880 36120 5880 36120 0 _0106_
rlabel metal2 6104 39088 6104 39088 0 _0107_
rlabel metal2 24080 37016 24080 37016 0 _0108_
rlabel metal2 28616 40488 28616 40488 0 _0109_
rlabel metal2 26040 40824 26040 40824 0 _0110_
rlabel metal2 25704 43932 25704 43932 0 _0111_
rlabel metal3 28952 43400 28952 43400 0 _0112_
rlabel metal2 32872 43176 32872 43176 0 _0113_
rlabel metal2 33208 41608 33208 41608 0 _0114_
rlabel metal2 35672 43176 35672 43176 0 _0115_
rlabel metal2 41720 41496 41720 41496 0 _0116_
rlabel metal2 36568 39368 36568 39368 0 _0117_
rlabel metal2 39368 39816 39368 39816 0 _0118_
rlabel metal2 41720 42840 41720 42840 0 _0119_
rlabel metal2 40936 43932 40936 43932 0 _0120_
rlabel metal2 38248 41496 38248 41496 0 _0121_
rlabel metal2 41496 42728 41496 42728 0 _0122_
rlabel metal3 45640 40544 45640 40544 0 _0123_
rlabel metal2 6440 33488 6440 33488 0 _0124_
rlabel metal2 9800 25088 9800 25088 0 _0125_
rlabel metal2 9800 23576 9800 23576 0 _0126_
rlabel metal2 9632 21784 9632 21784 0 _0127_
rlabel metal2 6664 19992 6664 19992 0 _0128_
rlabel metal2 2520 18760 2520 18760 0 _0129_
rlabel metal2 2520 19600 2520 19600 0 _0130_
rlabel metal2 3640 21000 3640 21000 0 _0131_
rlabel metal2 2520 23464 2520 23464 0 _0132_
rlabel metal2 3864 25144 3864 25144 0 _0133_
rlabel metal2 2520 26768 2520 26768 0 _0134_
rlabel metal2 3864 28280 3864 28280 0 _0135_
rlabel metal3 4816 30072 4816 30072 0 _0136_
rlabel metal2 2520 30800 2520 30800 0 _0137_
rlabel metal2 4424 29960 4424 29960 0 _0138_
rlabel metal2 8120 29848 8120 29848 0 _0139_
rlabel metal2 8344 28336 8344 28336 0 _0140_
rlabel metal2 6440 25928 6440 25928 0 _0141_
rlabel metal2 22288 13832 22288 13832 0 _0142_
rlabel metal2 24752 16184 24752 16184 0 _0143_
rlabel metal3 24528 15176 24528 15176 0 _0144_
rlabel metal2 24640 11480 24640 11480 0 _0145_
rlabel metal2 22680 10080 22680 10080 0 _0146_
rlabel metal2 25872 10696 25872 10696 0 _0147_
rlabel metal2 8904 39144 8904 39144 0 _0148_
rlabel metal2 14056 32872 14056 32872 0 _0149_
rlabel metal2 9576 32088 9576 32088 0 _0150_
rlabel metal3 11480 34328 11480 34328 0 _0151_
rlabel metal2 12040 30632 12040 30632 0 _0152_
rlabel metal3 36288 16744 36288 16744 0 _0153_
rlabel metal2 34328 13440 34328 13440 0 _0154_
rlabel metal2 39592 14168 39592 14168 0 _0155_
rlabel metal2 45416 11368 45416 11368 0 _0156_
rlabel metal2 45360 9128 45360 9128 0 _0157_
rlabel metal2 43512 9744 43512 9744 0 _0158_
rlabel metal2 45472 4424 45472 4424 0 _0159_
rlabel metal2 45416 6216 45416 6216 0 _0160_
rlabel metal2 42280 4312 42280 4312 0 _0161_
rlabel metal2 35448 3584 35448 3584 0 _0162_
rlabel metal3 44184 5208 44184 5208 0 _0163_
rlabel metal2 37072 7560 37072 7560 0 _0164_
rlabel metal2 24584 18816 24584 18816 0 _0165_
rlabel metal2 35336 21896 35336 21896 0 _0166_
rlabel metal2 31864 24248 31864 24248 0 _0167_
rlabel metal2 34216 25928 34216 25928 0 _0168_
rlabel metal2 38472 28168 38472 28168 0 _0169_
rlabel metal2 45304 27720 45304 27720 0 _0170_
rlabel metal2 43736 24360 43736 24360 0 _0171_
rlabel metal2 45360 23240 45360 23240 0 _0172_
rlabel metal2 44184 21952 44184 21952 0 _0173_
rlabel metal3 44184 20664 44184 20664 0 _0174_
rlabel metal3 44184 19096 44184 19096 0 _0175_
rlabel metal2 41160 20888 41160 20888 0 _0176_
rlabel metal2 44072 17304 44072 17304 0 _0177_
rlabel metal2 28728 21896 28728 21896 0 _0178_
rlabel metal2 14280 36848 14280 36848 0 _0179_
rlabel metal2 15848 35448 15848 35448 0 _0180_
rlabel metal3 14784 38696 14784 38696 0 _0181_
rlabel metal2 13496 40040 13496 40040 0 _0182_
rlabel metal2 16464 42168 16464 42168 0 _0183_
rlabel metal2 14728 43176 14728 43176 0 _0184_
rlabel metal2 11144 40656 11144 40656 0 _0185_
rlabel metal2 11480 43176 11480 43176 0 _0186_
rlabel metal2 6664 43176 6664 43176 0 _0187_
rlabel metal2 6664 42280 6664 42280 0 _0188_
rlabel metal2 6888 40040 6888 40040 0 _0189_
rlabel metal2 10976 38696 10976 38696 0 _0190_
rlabel metal2 21000 29568 21000 29568 0 _0191_
rlabel metal2 21896 21504 21896 21504 0 _0192_
rlabel metal3 17752 23464 17752 23464 0 _0193_
rlabel metal2 10192 26936 10192 26936 0 _0194_
rlabel metal3 11368 28728 11368 28728 0 _0195_
rlabel metal2 11480 25144 11480 25144 0 _0196_
rlabel metal2 14840 24136 14840 24136 0 _0197_
rlabel metal2 13272 21616 13272 21616 0 _0198_
rlabel metal2 11928 18368 11928 18368 0 _0199_
rlabel metal2 10920 17752 10920 17752 0 _0200_
rlabel metal2 22680 31080 22680 31080 0 _0201_
rlabel metal2 22792 29344 22792 29344 0 _0202_
rlabel metal4 26264 27384 26264 27384 0 _0203_
rlabel metal2 29960 29344 29960 29344 0 _0204_
rlabel metal2 29568 31080 29568 31080 0 _0205_
rlabel metal2 25480 33656 25480 33656 0 _0206_
rlabel metal2 26376 34552 26376 34552 0 _0207_
rlabel metal2 28280 36008 28280 36008 0 _0208_
rlabel metal2 30520 33880 30520 33880 0 _0209_
rlabel metal2 33208 32704 33208 32704 0 _0210_
rlabel metal2 32760 35224 32760 35224 0 _0211_
rlabel metal2 31528 36736 31528 36736 0 _0212_
rlabel metal2 33936 35784 33936 35784 0 _0213_
rlabel metal2 15960 16520 15960 16520 0 _0214_
rlabel metal2 10360 17192 10360 17192 0 _0215_
rlabel metal2 10584 16464 10584 16464 0 _0216_
rlabel metal3 7840 13944 7840 13944 0 _0217_
rlabel metal3 9016 14616 9016 14616 0 _0218_
rlabel metal2 11984 14616 11984 14616 0 _0219_
rlabel metal2 10136 11760 10136 11760 0 _0220_
rlabel metal2 13496 12488 13496 12488 0 _0221_
rlabel metal2 21224 20384 21224 20384 0 _0222_
rlabel metal3 22232 21448 22232 21448 0 _0223_
rlabel metal3 45472 40376 45472 40376 0 _0224_
rlabel metal2 45416 40992 45416 40992 0 _0225_
rlabel metal2 9408 33432 9408 33432 0 _0226_
rlabel metal2 7672 35224 7672 35224 0 _0227_
rlabel metal3 7952 34104 7952 34104 0 _0228_
rlabel metal2 7448 34272 7448 34272 0 _0229_
rlabel metal3 6720 34104 6720 34104 0 _0230_
rlabel metal3 8232 19208 8232 19208 0 _0231_
rlabel metal2 8904 20328 8904 20328 0 _0232_
rlabel metal2 8008 24864 8008 24864 0 _0233_
rlabel metal3 9072 24696 9072 24696 0 _0234_
rlabel metal2 6440 23688 6440 23688 0 _0235_
rlabel metal2 6104 23856 6104 23856 0 _0236_
rlabel metal3 7560 24808 7560 24808 0 _0237_
rlabel metal2 9016 24024 9016 24024 0 _0238_
rlabel metal2 10136 22400 10136 22400 0 _0239_
rlabel metal3 10136 23128 10136 23128 0 _0240_
rlabel metal2 9184 23128 9184 23128 0 _0241_
rlabel metal3 8960 21560 8960 21560 0 _0242_
rlabel metal2 9072 21560 9072 21560 0 _0243_
rlabel metal2 5320 20664 5320 20664 0 _0244_
rlabel metal2 2744 21224 2744 21224 0 _0245_
rlabel metal2 6440 19712 6440 19712 0 _0246_
rlabel metal2 6776 20384 6776 20384 0 _0247_
rlabel metal2 3304 20496 3304 20496 0 _0248_
rlabel metal2 3080 18704 3080 18704 0 _0249_
rlabel metal2 5880 19040 5880 19040 0 _0250_
rlabel metal2 4200 19152 4200 19152 0 _0251_
rlabel metal2 2128 20552 2128 20552 0 _0252_
rlabel metal2 5544 19600 5544 19600 0 _0253_
rlabel metal3 3304 20664 3304 20664 0 _0254_
rlabel metal2 3976 21448 3976 21448 0 _0255_
rlabel metal2 3080 27104 3080 27104 0 _0256_
rlabel metal2 3864 24192 3864 24192 0 _0257_
rlabel metal3 4536 23352 4536 23352 0 _0258_
rlabel metal2 4144 23912 4144 23912 0 _0259_
rlabel metal2 3192 25592 3192 25592 0 _0260_
rlabel metal3 2800 24696 2800 24696 0 _0261_
rlabel metal2 3640 24696 3640 24696 0 _0262_
rlabel metal2 3192 27216 3192 27216 0 _0263_
rlabel metal2 4424 26320 4424 26320 0 _0264_
rlabel metal3 4760 27832 4760 27832 0 _0265_
rlabel metal2 2856 28672 2856 28672 0 _0266_
rlabel metal3 3220 29400 3220 29400 0 _0267_
rlabel metal2 3248 29176 3248 29176 0 _0268_
rlabel metal2 5656 29624 5656 29624 0 _0269_
rlabel metal3 8512 31640 8512 31640 0 _0270_
rlabel metal3 7784 29624 7784 29624 0 _0271_
rlabel metal2 6888 26852 6888 26852 0 _0272_
rlabel metal2 6440 30464 6440 30464 0 _0273_
rlabel metal2 8232 31136 8232 31136 0 _0274_
rlabel metal2 6776 31640 6776 31640 0 _0275_
rlabel metal2 7672 29232 7672 29232 0 _0276_
rlabel metal2 7952 29512 7952 29512 0 _0277_
rlabel metal3 8288 27832 8288 27832 0 _0278_
rlabel metal2 7448 28224 7448 28224 0 _0279_
rlabel metal3 6272 22456 6272 22456 0 _0280_
rlabel metal2 6328 28000 6328 28000 0 _0281_
rlabel metal2 6496 27944 6496 27944 0 _0282_
rlabel metal2 6384 23128 6384 23128 0 _0283_
rlabel metal2 7392 23128 7392 23128 0 _0284_
rlabel metal2 6888 23632 6888 23632 0 _0285_
rlabel metal2 7448 24024 7448 24024 0 _0286_
rlabel metal2 7784 24080 7784 24080 0 _0287_
rlabel metal2 7336 25144 7336 25144 0 _0288_
rlabel metal2 27048 13216 27048 13216 0 _0289_
rlabel metal2 27608 15456 27608 15456 0 _0290_
rlabel metal2 27104 16968 27104 16968 0 _0291_
rlabel metal3 28224 15288 28224 15288 0 _0292_
rlabel metal3 27944 15456 27944 15456 0 _0293_
rlabel metal2 27216 16632 27216 16632 0 _0294_
rlabel metal2 29064 14000 29064 14000 0 _0295_
rlabel metal3 27440 13832 27440 13832 0 _0296_
rlabel metal2 30072 13832 30072 13832 0 _0297_
rlabel metal2 25592 12264 25592 12264 0 _0298_
rlabel metal2 27944 13160 27944 13160 0 _0299_
rlabel metal3 29456 12152 29456 12152 0 _0300_
rlabel metal2 23576 13888 23576 13888 0 _0301_
rlabel metal2 22008 12656 22008 12656 0 _0302_
rlabel metal3 24752 15288 24752 15288 0 _0303_
rlabel metal2 24360 16800 24360 16800 0 _0304_
rlabel metal3 25088 17080 25088 17080 0 _0305_
rlabel metal3 26208 15176 26208 15176 0 _0306_
rlabel metal2 26712 19264 26712 19264 0 _0307_
rlabel metal2 25816 15400 25816 15400 0 _0308_
rlabel metal3 24864 13496 24864 13496 0 _0309_
rlabel metal3 25536 13720 25536 13720 0 _0310_
rlabel metal3 24864 12152 24864 12152 0 _0311_
rlabel metal2 23688 12096 23688 12096 0 _0312_
rlabel metal2 23016 10864 23016 10864 0 _0313_
rlabel metal2 13720 31360 13720 31360 0 _0314_
rlabel metal2 12824 33712 12824 33712 0 _0315_
rlabel metal2 10584 32368 10584 32368 0 _0316_
rlabel metal3 11424 33992 11424 33992 0 _0317_
rlabel metal2 11928 30856 11928 30856 0 _0318_
rlabel metal2 36120 17360 36120 17360 0 _0319_
rlabel metal2 35672 16800 35672 16800 0 _0320_
rlabel metal2 15960 30688 15960 30688 0 _0321_
rlabel metal2 36456 4144 36456 4144 0 _0322_
rlabel metal2 38920 7224 38920 7224 0 _0323_
rlabel metal2 38584 7784 38584 7784 0 _0324_
rlabel metal2 42952 3976 42952 3976 0 _0325_
rlabel metal2 41944 6384 41944 6384 0 _0326_
rlabel metal3 40656 5992 40656 5992 0 _0327_
rlabel metal3 39984 10584 39984 10584 0 _0328_
rlabel metal2 38808 9464 38808 9464 0 _0329_
rlabel metal3 35784 11256 35784 11256 0 _0330_
rlabel metal2 36568 10864 36568 10864 0 _0331_
rlabel metal2 43960 15484 43960 15484 0 _0332_
rlabel metal2 34104 7728 34104 7728 0 _0333_
rlabel metal2 39144 9072 39144 9072 0 _0334_
rlabel metal2 37968 8792 37968 8792 0 _0335_
rlabel metal2 38584 11648 38584 11648 0 _0336_
rlabel metal2 39032 12040 39032 12040 0 _0337_
rlabel metal2 38808 11424 38808 11424 0 _0338_
rlabel metal2 38696 11704 38696 11704 0 _0339_
rlabel metal2 39256 12208 39256 12208 0 _0340_
rlabel metal2 37800 11424 37800 11424 0 _0341_
rlabel metal2 38080 9016 38080 9016 0 _0342_
rlabel metal2 38472 8232 38472 8232 0 _0343_
rlabel metal2 40152 11872 40152 11872 0 _0344_
rlabel metal3 41608 12936 41608 12936 0 _0345_
rlabel metal2 40040 9744 40040 9744 0 _0346_
rlabel metal2 42168 10248 42168 10248 0 _0347_
rlabel metal2 41496 11872 41496 11872 0 _0348_
rlabel metal2 39480 9856 39480 9856 0 _0349_
rlabel metal2 37576 12208 37576 12208 0 _0350_
rlabel metal2 39032 9912 39032 9912 0 _0351_
rlabel metal2 41328 6104 41328 6104 0 _0352_
rlabel metal2 40040 10360 40040 10360 0 _0353_
rlabel metal2 42280 6104 42280 6104 0 _0354_
rlabel metal2 40264 9800 40264 9800 0 _0355_
rlabel metal3 39424 9800 39424 9800 0 _0356_
rlabel metal2 38696 9016 38696 9016 0 _0357_
rlabel metal3 39592 7560 39592 7560 0 _0358_
rlabel metal2 39928 11032 39928 11032 0 _0359_
rlabel metal2 36232 11648 36232 11648 0 _0360_
rlabel metal2 40208 11256 40208 11256 0 _0361_
rlabel metal3 40320 9800 40320 9800 0 _0362_
rlabel metal2 41104 8456 41104 8456 0 _0363_
rlabel metal2 39592 9408 39592 9408 0 _0364_
rlabel metal2 40264 8064 40264 8064 0 _0365_
rlabel metal2 40040 7952 40040 7952 0 _0366_
rlabel metal2 40264 6216 40264 6216 0 _0367_
rlabel metal2 34552 17080 34552 17080 0 _0368_
rlabel metal2 34776 16296 34776 16296 0 _0369_
rlabel metal2 38696 15344 38696 15344 0 _0370_
rlabel metal2 42168 13608 42168 13608 0 _0371_
rlabel metal2 36120 14056 36120 14056 0 _0372_
rlabel metal3 32928 20552 32928 20552 0 _0373_
rlabel metal2 34888 13272 34888 13272 0 _0374_
rlabel metal2 34440 12600 34440 12600 0 _0375_
rlabel metal2 38920 14448 38920 14448 0 _0376_
rlabel metal2 39256 14448 39256 14448 0 _0377_
rlabel metal2 41272 13888 41272 13888 0 _0378_
rlabel metal2 41720 14336 41720 14336 0 _0379_
rlabel metal3 42112 13720 42112 13720 0 _0380_
rlabel metal2 42504 14056 42504 14056 0 _0381_
rlabel metal2 42952 14168 42952 14168 0 _0382_
rlabel metal3 43456 12936 43456 12936 0 _0383_
rlabel metal2 44856 12040 44856 12040 0 _0384_
rlabel metal2 35112 8176 35112 8176 0 _0385_
rlabel metal2 42728 11312 42728 11312 0 _0386_
rlabel metal2 41664 11592 41664 11592 0 _0387_
rlabel metal3 42224 11368 42224 11368 0 _0388_
rlabel metal2 42392 11256 42392 11256 0 _0389_
rlabel metal3 43456 11368 43456 11368 0 _0390_
rlabel metal2 23968 26488 23968 26488 0 _0391_
rlabel metal2 42840 9072 42840 9072 0 _0392_
rlabel metal2 43624 7112 43624 7112 0 _0393_
rlabel metal3 45024 6440 45024 6440 0 _0394_
rlabel metal3 44016 8232 44016 8232 0 _0395_
rlabel metal3 45696 8232 45696 8232 0 _0396_
rlabel metal2 40488 6720 40488 6720 0 _0397_
rlabel metal2 40824 5712 40824 5712 0 _0398_
rlabel metal2 45640 9744 45640 9744 0 _0399_
rlabel metal2 40152 4648 40152 4648 0 _0400_
rlabel metal2 40824 4256 40824 4256 0 _0401_
rlabel metal2 39592 3808 39592 3808 0 _0402_
rlabel metal3 43792 4424 43792 4424 0 _0403_
rlabel metal2 45416 5544 45416 5544 0 _0404_
rlabel metal2 37688 8568 37688 8568 0 _0405_
rlabel metal3 27216 19992 27216 19992 0 _0406_
rlabel metal2 27832 20384 27832 20384 0 _0407_
rlabel metal3 38024 23688 38024 23688 0 _0408_
rlabel metal2 35112 21952 35112 21952 0 _0409_
rlabel metal2 38976 20552 38976 20552 0 _0410_
rlabel metal2 39928 20608 39928 20608 0 _0411_
rlabel metal2 39592 21168 39592 21168 0 _0412_
rlabel metal3 39984 21784 39984 21784 0 _0413_
rlabel metal3 43344 23688 43344 23688 0 _0414_
rlabel metal3 41944 24696 41944 24696 0 _0415_
rlabel metal3 41720 24808 41720 24808 0 _0416_
rlabel metal2 40376 26600 40376 26600 0 _0417_
rlabel metal3 43512 27832 43512 27832 0 _0418_
rlabel metal2 40824 27160 40824 27160 0 _0419_
rlabel metal3 40992 25592 40992 25592 0 _0420_
rlabel metal2 39704 24584 39704 24584 0 _0421_
rlabel metal2 37744 26488 37744 26488 0 _0422_
rlabel metal2 37128 26264 37128 26264 0 _0423_
rlabel metal2 38920 25816 38920 25816 0 _0424_
rlabel metal2 35896 23184 35896 23184 0 _0425_
rlabel metal2 34496 24472 34496 24472 0 _0426_
rlabel metal3 36568 24696 36568 24696 0 _0427_
rlabel metal2 37520 23912 37520 23912 0 _0428_
rlabel metal2 35280 23912 35280 23912 0 _0429_
rlabel metal2 38304 23352 38304 23352 0 _0430_
rlabel metal2 37688 24976 37688 24976 0 _0431_
rlabel metal2 38248 25256 38248 25256 0 _0432_
rlabel metal2 39928 27552 39928 27552 0 _0433_
rlabel metal2 39032 27272 39032 27272 0 _0434_
rlabel metal2 41944 26992 41944 26992 0 _0435_
rlabel metal2 39592 26376 39592 26376 0 _0436_
rlabel metal2 39256 25760 39256 25760 0 _0437_
rlabel metal2 39424 23912 39424 23912 0 _0438_
rlabel metal3 44688 25480 44688 25480 0 _0439_
rlabel metal3 45136 24136 45136 24136 0 _0440_
rlabel metal2 41160 24864 41160 24864 0 _0441_
rlabel metal2 39592 24752 39592 24752 0 _0442_
rlabel metal2 41048 22848 41048 22848 0 _0443_
rlabel metal3 40880 23352 40880 23352 0 _0444_
rlabel metal2 40488 24360 40488 24360 0 _0445_
rlabel metal2 40376 24752 40376 24752 0 _0446_
rlabel metal2 39928 22232 39928 22232 0 _0447_
rlabel metal2 44408 18312 44408 18312 0 _0448_
rlabel metal3 41216 18648 41216 18648 0 _0449_
rlabel metal2 38696 19712 38696 19712 0 _0450_
rlabel metal2 40264 19432 40264 19432 0 _0451_
rlabel metal2 39928 19040 39928 19040 0 _0452_
rlabel metal2 39816 19992 39816 19992 0 _0453_
rlabel metal2 38808 20216 38808 20216 0 _0454_
rlabel metal2 38976 21784 38976 21784 0 _0455_
rlabel metal2 39816 22008 39816 22008 0 _0456_
rlabel metal2 39368 21784 39368 21784 0 _0457_
rlabel metal2 38136 23128 38136 23128 0 _0458_
rlabel metal2 41048 24080 41048 24080 0 _0459_
rlabel metal3 38920 23128 38920 23128 0 _0460_
rlabel metal2 39424 23128 39424 23128 0 _0461_
rlabel metal2 40040 22624 40040 22624 0 _0462_
rlabel metal2 31864 22792 31864 22792 0 _0463_
rlabel metal2 37800 22400 37800 22400 0 _0464_
rlabel metal3 44520 21000 44520 21000 0 _0465_
rlabel metal2 35672 21616 35672 21616 0 _0466_
rlabel metal2 40936 20720 40936 20720 0 _0467_
rlabel metal2 35448 24472 35448 24472 0 _0468_
rlabel metal2 35672 23408 35672 23408 0 _0469_
rlabel metal2 38808 25872 38808 25872 0 _0470_
rlabel metal2 41832 26684 41832 26684 0 _0471_
rlabel metal2 35784 25536 35784 25536 0 _0472_
rlabel metal2 45080 24528 45080 24528 0 _0473_
rlabel metal2 37968 27720 37968 27720 0 _0474_
rlabel metal2 42168 26712 42168 26712 0 _0475_
rlabel metal3 43960 25704 43960 25704 0 _0476_
rlabel metal2 43848 27216 43848 27216 0 _0477_
rlabel metal2 43456 24136 43456 24136 0 _0478_
rlabel metal2 42504 24920 42504 24920 0 _0479_
rlabel metal2 44856 24360 44856 24360 0 _0480_
rlabel metal2 43848 22736 43848 22736 0 _0481_
rlabel metal3 43456 22456 43456 22456 0 _0482_
rlabel metal2 45192 21168 45192 21168 0 _0483_
rlabel metal2 45304 21560 45304 21560 0 _0484_
rlabel metal3 45528 19208 45528 19208 0 _0485_
rlabel metal2 45304 18984 45304 18984 0 _0486_
rlabel metal2 40712 20412 40712 20412 0 _0487_
rlabel metal2 44912 18536 44912 18536 0 _0488_
rlabel metal2 29736 22120 29736 22120 0 _0489_
rlabel metal2 29624 21560 29624 21560 0 _0490_
rlabel metal2 17976 35728 17976 35728 0 _0491_
rlabel metal2 17528 36064 17528 36064 0 _0492_
rlabel metal3 10976 39816 10976 39816 0 _0493_
rlabel metal2 24416 40600 24416 40600 0 _0494_
rlabel metal2 21672 40544 21672 40544 0 _0495_
rlabel metal2 18088 41440 18088 41440 0 _0496_
rlabel metal2 19208 40488 19208 40488 0 _0497_
rlabel metal2 18424 39200 18424 39200 0 _0498_
rlabel metal2 19096 34496 19096 34496 0 _0499_
rlabel metal2 18984 34272 18984 34272 0 _0500_
rlabel metal2 19320 36064 19320 36064 0 _0501_
rlabel metal4 17416 36232 17416 36232 0 _0502_
rlabel metal2 17304 36064 17304 36064 0 _0503_
rlabel metal3 20496 38808 20496 38808 0 _0504_
rlabel metal2 16856 40600 16856 40600 0 _0505_
rlabel metal3 21336 38864 21336 38864 0 _0506_
rlabel metal2 20216 39088 20216 39088 0 _0507_
rlabel metal2 20664 39872 20664 39872 0 _0508_
rlabel metal2 24528 40936 24528 40936 0 _0509_
rlabel metal2 15512 41776 15512 41776 0 _0510_
rlabel metal2 18200 41496 18200 41496 0 _0511_
rlabel metal2 17864 42392 17864 42392 0 _0512_
rlabel metal3 21896 40936 21896 40936 0 _0513_
rlabel metal3 20664 44072 20664 44072 0 _0514_
rlabel metal2 21896 42840 21896 42840 0 _0515_
rlabel metal3 22344 43624 22344 43624 0 _0516_
rlabel metal2 21840 40376 21840 40376 0 _0517_
rlabel metal2 20216 40432 20216 40432 0 _0518_
rlabel metal3 22400 38024 22400 38024 0 _0519_
rlabel metal2 19320 39928 19320 39928 0 _0520_
rlabel metal3 20496 38024 20496 38024 0 _0521_
rlabel metal2 23912 37184 23912 37184 0 _0522_
rlabel metal2 20776 37352 20776 37352 0 _0523_
rlabel metal3 14280 39592 14280 39592 0 _0524_
rlabel metal3 11984 42728 11984 42728 0 _0525_
rlabel metal2 13384 38808 13384 38808 0 _0526_
rlabel metal2 15344 38696 15344 38696 0 _0527_
rlabel metal2 17864 36176 17864 36176 0 _0528_
rlabel metal3 17584 35672 17584 35672 0 _0529_
rlabel metal2 15512 38752 15512 38752 0 _0530_
rlabel metal2 16520 39256 16520 39256 0 _0531_
rlabel metal2 15904 40488 15904 40488 0 _0532_
rlabel metal2 11256 39984 11256 39984 0 _0533_
rlabel metal2 14728 39480 14728 39480 0 _0534_
rlabel metal2 16408 41944 16408 41944 0 _0535_
rlabel metal2 16184 43932 16184 43932 0 _0536_
rlabel metal2 14280 44296 14280 44296 0 _0537_
rlabel metal2 15848 44044 15848 44044 0 _0538_
rlabel metal2 11480 40656 11480 40656 0 _0539_
rlabel metal2 9800 43932 9800 43932 0 _0540_
rlabel metal3 12880 44072 12880 44072 0 _0541_
rlabel metal2 10416 44408 10416 44408 0 _0542_
rlabel metal2 9352 41720 9352 41720 0 _0543_
rlabel metal2 10248 40936 10248 40936 0 _0544_
rlabel metal2 9744 41384 9744 41384 0 _0545_
rlabel metal2 11032 40040 11032 40040 0 _0546_
rlabel metal2 11144 38136 11144 38136 0 _0547_
rlabel metal2 23240 28448 23240 28448 0 _0548_
rlabel metal2 22512 22904 22512 22904 0 _0549_
rlabel metal2 23128 22848 23128 22848 0 _0550_
rlabel metal2 21112 21000 21112 21000 0 _0551_
rlabel metal2 19320 23912 19320 23912 0 _0552_
rlabel metal2 14840 24752 14840 24752 0 _0553_
rlabel metal2 13384 27776 13384 27776 0 _0554_
rlabel metal3 11256 28616 11256 28616 0 _0555_
rlabel metal2 12712 24360 12712 24360 0 _0556_
rlabel metal3 13384 23912 13384 23912 0 _0557_
rlabel metal2 13608 23520 13608 23520 0 _0558_
rlabel metal2 13944 16576 13944 16576 0 _0559_
rlabel metal2 14336 24024 14336 24024 0 _0560_
rlabel metal2 15400 21056 15400 21056 0 _0561_
rlabel metal2 13832 21336 13832 21336 0 _0562_
rlabel metal2 12040 19600 12040 19600 0 _0563_
rlabel metal2 12264 18816 12264 18816 0 _0564_
rlabel metal2 13608 19320 13608 19320 0 _0565_
rlabel metal2 42616 31360 42616 31360 0 _0566_
rlabel metal2 24584 31080 24584 31080 0 _0567_
rlabel metal3 24864 32648 24864 32648 0 _0568_
rlabel metal2 23800 31304 23800 31304 0 _0569_
rlabel metal2 23632 29176 23632 29176 0 _0570_
rlabel metal2 25928 30128 25928 30128 0 _0571_
rlabel metal3 24920 29624 24920 29624 0 _0572_
rlabel metal2 24584 28280 24584 28280 0 _0573_
rlabel metal2 27272 30240 27272 30240 0 _0574_
rlabel metal2 27384 32200 27384 32200 0 _0575_
rlabel metal2 30128 32312 30128 32312 0 _0576_
rlabel metal2 29288 36064 29288 36064 0 _0577_
rlabel metal2 31528 33488 31528 33488 0 _0578_
rlabel metal3 28952 33208 28952 33208 0 _0579_
rlabel metal2 26040 33712 26040 33712 0 _0580_
rlabel metal2 26488 34832 26488 34832 0 _0581_
rlabel metal2 31080 36120 31080 36120 0 _0582_
rlabel metal3 32144 33432 32144 33432 0 _0583_
rlabel metal2 31864 34888 31864 34888 0 _0584_
rlabel metal2 32312 33432 32312 33432 0 _0585_
rlabel metal2 32312 32480 32312 32480 0 _0586_
rlabel metal2 33432 34944 33432 34944 0 _0587_
rlabel metal2 32200 36400 32200 36400 0 _0588_
rlabel metal2 32200 34944 32200 34944 0 _0589_
rlabel metal2 15624 17976 15624 17976 0 _0590_
rlabel metal2 14392 16856 14392 16856 0 _0591_
rlabel metal2 11312 16296 11312 16296 0 _0592_
rlabel metal3 12936 13720 12936 13720 0 _0593_
rlabel metal3 12096 16744 12096 16744 0 _0594_
rlabel metal2 9968 13720 9968 13720 0 _0595_
rlabel metal3 10080 15960 10080 15960 0 _0596_
rlabel metal3 10808 13944 10808 13944 0 _0597_
rlabel metal3 9632 15176 9632 15176 0 _0598_
rlabel metal2 11592 14056 11592 14056 0 _0599_
rlabel metal2 11816 14448 11816 14448 0 _0600_
rlabel metal2 10584 14168 10584 14168 0 _0601_
rlabel metal3 13048 14392 13048 14392 0 _0602_
rlabel metal2 11480 12768 11480 12768 0 _0603_
rlabel metal2 10528 12040 10528 12040 0 _0604_
rlabel metal2 13720 13048 13720 13048 0 _0605_
rlabel metal2 24360 21952 24360 21952 0 _0606_
rlabel metal2 24024 22344 24024 22344 0 _0607_
rlabel metal2 17640 26544 17640 26544 0 _0608_
rlabel metal2 19096 21056 19096 21056 0 _0609_
rlabel metal2 23688 20776 23688 20776 0 _0610_
rlabel metal2 22568 21784 22568 21784 0 _0611_
rlabel metal2 23800 22176 23800 22176 0 _0612_
rlabel metal2 25032 20888 25032 20888 0 _0613_
rlabel metal2 18984 20608 18984 20608 0 _0614_
rlabel metal2 17640 19208 17640 19208 0 _0615_
rlabel metal3 22680 26264 22680 26264 0 _0616_
rlabel metal2 19656 26600 19656 26600 0 _0617_
rlabel metal3 19320 19320 19320 19320 0 _0618_
rlabel metal2 16408 22232 16408 22232 0 _0619_
rlabel metal2 21784 23072 21784 23072 0 _0620_
rlabel metal2 19656 22848 19656 22848 0 _0621_
rlabel metal2 19320 20160 19320 20160 0 _0622_
rlabel metal2 18200 16632 18200 16632 0 _0623_
rlabel metal2 20552 18592 20552 18592 0 _0624_
rlabel metal2 15288 18648 15288 18648 0 _0625_
rlabel metal2 17752 16520 17752 16520 0 _0626_
rlabel metal3 19096 16184 19096 16184 0 _0627_
rlabel metal2 18088 15680 18088 15680 0 _0628_
rlabel metal3 23464 29400 23464 29400 0 _0629_
rlabel metal2 30408 20216 30408 20216 0 _0630_
rlabel metal2 30968 28224 30968 28224 0 _0631_
rlabel metal2 29792 23912 29792 23912 0 _0632_
rlabel metal2 26152 27888 26152 27888 0 _0633_
rlabel metal2 24696 31976 24696 31976 0 _0634_
rlabel metal2 26600 29960 26600 29960 0 _0635_
rlabel metal2 25704 23184 25704 23184 0 _0636_
rlabel metal2 29176 18536 29176 18536 0 _0637_
rlabel metal3 30072 16184 30072 16184 0 _0638_
rlabel metal2 22008 19096 22008 19096 0 _0639_
rlabel metal2 23464 22344 23464 22344 0 _0640_
rlabel metal2 29848 18032 29848 18032 0 _0641_
rlabel metal2 29736 16744 29736 16744 0 _0642_
rlabel metal2 30296 16184 30296 16184 0 _0643_
rlabel metal2 30184 7952 30184 7952 0 _0644_
rlabel metal3 30632 14616 30632 14616 0 _0645_
rlabel metal3 31976 17640 31976 17640 0 _0646_
rlabel metal3 29792 12376 29792 12376 0 _0647_
rlabel metal2 33544 17248 33544 17248 0 _0648_
rlabel metal3 28896 12040 28896 12040 0 _0649_
rlabel metal2 39816 32984 39816 32984 0 _0650_
rlabel metal2 38696 23128 38696 23128 0 _0651_
rlabel metal2 27944 18032 27944 18032 0 _0652_
rlabel metal2 25480 29456 25480 29456 0 _0653_
rlabel metal2 28280 28448 28280 28448 0 _0654_
rlabel metal2 22568 23408 22568 23408 0 _0655_
rlabel metal3 30072 16520 30072 16520 0 _0656_
rlabel metal2 34328 5208 34328 5208 0 _0657_
rlabel metal3 10696 38696 10696 38696 0 _0658_
rlabel metal2 44184 16464 44184 16464 0 _0659_
rlabel metal3 32312 7560 32312 7560 0 _0660_
rlabel metal2 32312 7672 32312 7672 0 _0661_
rlabel metal2 32424 4872 32424 4872 0 _0662_
rlabel metal2 35560 5208 35560 5208 0 _0663_
rlabel metal2 34552 6272 34552 6272 0 _0664_
rlabel metal2 26152 21952 26152 21952 0 _0665_
rlabel metal3 20832 20776 20832 20776 0 _0666_
rlabel metal2 22904 29456 22904 29456 0 _0667_
rlabel metal2 24248 32088 24248 32088 0 _0668_
rlabel metal2 23968 32760 23968 32760 0 _0669_
rlabel metal2 20664 36792 20664 36792 0 _0670_
rlabel metal2 22792 18816 22792 18816 0 _0671_
rlabel metal2 23016 33712 23016 33712 0 _0672_
rlabel metal2 20216 32032 20216 32032 0 _0673_
rlabel metal2 23408 24808 23408 24808 0 _0674_
rlabel metal2 23800 34216 23800 34216 0 _0675_
rlabel metal2 23688 40264 23688 40264 0 _0676_
rlabel metal2 24752 26488 24752 26488 0 _0677_
rlabel metal3 24640 33880 24640 33880 0 _0678_
rlabel metal3 18088 15400 18088 15400 0 _0679_
rlabel metal2 14952 14000 14952 14000 0 _0680_
rlabel metal2 16912 15512 16912 15512 0 _0681_
rlabel metal2 21224 34104 21224 34104 0 _0682_
rlabel metal2 26712 30464 26712 30464 0 _0683_
rlabel metal3 23072 34104 23072 34104 0 _0684_
rlabel metal3 22120 36232 22120 36232 0 _0685_
rlabel metal2 22568 36008 22568 36008 0 _0686_
rlabel metal2 21896 36512 21896 36512 0 _0687_
rlabel metal2 22176 17752 22176 17752 0 _0688_
rlabel metal2 8008 10640 8008 10640 0 _0689_
rlabel metal2 18760 15512 18760 15512 0 _0690_
rlabel metal2 19544 17752 19544 17752 0 _0691_
rlabel metal2 19208 17640 19208 17640 0 _0692_
rlabel metal2 19992 15400 19992 15400 0 _0693_
rlabel metal2 18928 16632 18928 16632 0 _0694_
rlabel metal2 18984 15484 18984 15484 0 _0695_
rlabel metal2 19264 11144 19264 11144 0 _0696_
rlabel metal2 18424 11424 18424 11424 0 _0697_
rlabel metal2 6216 14000 6216 14000 0 _0698_
rlabel metal2 13832 13272 13832 13272 0 _0699_
rlabel metal2 18200 12600 18200 12600 0 _0700_
rlabel metal2 18760 12152 18760 12152 0 _0701_
rlabel metal2 17752 12824 17752 12824 0 _0702_
rlabel metal3 17808 12264 17808 12264 0 _0703_
rlabel metal2 16072 12376 16072 12376 0 _0704_
rlabel metal2 17192 12152 17192 12152 0 _0705_
rlabel metal2 15848 9576 15848 9576 0 _0706_
rlabel metal2 7112 9968 7112 9968 0 _0707_
rlabel metal2 16128 10696 16128 10696 0 _0708_
rlabel metal2 15064 10976 15064 10976 0 _0709_
rlabel metal2 13832 9408 13832 9408 0 _0710_
rlabel metal2 11872 9800 11872 9800 0 _0711_
rlabel metal3 14504 11256 14504 11256 0 _0712_
rlabel metal3 13160 11256 13160 11256 0 _0713_
rlabel metal3 11760 9912 11760 9912 0 _0714_
rlabel metal3 11200 8344 11200 8344 0 _0715_
rlabel metal2 11144 8372 11144 8372 0 _0716_
rlabel metal2 10640 8120 10640 8120 0 _0717_
rlabel metal2 21672 13104 21672 13104 0 _0718_
rlabel metal2 8288 5208 8288 5208 0 _0719_
rlabel metal3 13216 9016 13216 9016 0 _0720_
rlabel metal2 27608 5488 27608 5488 0 _0721_
rlabel metal2 23464 7168 23464 7168 0 _0722_
rlabel metal2 27048 5040 27048 5040 0 _0723_
rlabel metal2 20664 5320 20664 5320 0 _0724_
rlabel metal3 22568 7560 22568 7560 0 _0725_
rlabel metal2 22008 8288 22008 8288 0 _0726_
rlabel metal2 21000 7784 21000 7784 0 _0727_
rlabel metal2 24360 8960 24360 8960 0 _0728_
rlabel metal2 22512 8456 22512 8456 0 _0729_
rlabel metal3 25704 5096 25704 5096 0 _0730_
rlabel metal2 23464 6440 23464 6440 0 _0731_
rlabel metal2 17752 22064 17752 22064 0 _0732_
rlabel metal3 13552 8120 13552 8120 0 _0733_
rlabel metal3 13272 8008 13272 8008 0 _0734_
rlabel metal2 13608 6272 13608 6272 0 _0735_
rlabel metal2 19712 6440 19712 6440 0 _0736_
rlabel metal3 18648 7560 18648 7560 0 _0737_
rlabel metal2 20720 7672 20720 7672 0 _0738_
rlabel metal2 19880 7224 19880 7224 0 _0739_
rlabel metal2 16744 5712 16744 5712 0 _0740_
rlabel metal3 14224 6440 14224 6440 0 _0741_
rlabel metal2 12936 6944 12936 6944 0 _0742_
rlabel metal2 12040 6608 12040 6608 0 _0743_
rlabel metal3 13692 6888 13692 6888 0 _0744_
rlabel metal3 11704 3752 11704 3752 0 _0745_
rlabel metal2 9688 5544 9688 5544 0 _0746_
rlabel metal2 18760 5096 18760 5096 0 _0747_
rlabel metal2 16520 19992 16520 19992 0 _0748_
rlabel metal2 16744 19544 16744 19544 0 _0749_
rlabel metal2 16184 17416 16184 17416 0 _0750_
rlabel metal3 15848 15960 15848 15960 0 _0751_
rlabel metal2 4816 13160 4816 13160 0 _0752_
rlabel metal2 6104 13384 6104 13384 0 _0753_
rlabel metal2 5768 15680 5768 15680 0 _0754_
rlabel metal2 7560 12432 7560 12432 0 _0755_
rlabel metal2 7112 12208 7112 12208 0 _0756_
rlabel metal2 5656 10920 5656 10920 0 _0757_
rlabel metal2 5096 11928 5096 11928 0 _0758_
rlabel metal2 7784 10920 7784 10920 0 _0759_
rlabel metal2 7784 9520 7784 9520 0 _0760_
rlabel metal2 7672 9352 7672 9352 0 _0761_
rlabel metal2 8456 4200 8456 4200 0 _0762_
rlabel metal2 26096 26824 26096 26824 0 _0763_
rlabel metal2 30800 23688 30800 23688 0 _0764_
rlabel metal2 33712 15848 33712 15848 0 _0765_
rlabel metal2 22456 20552 22456 20552 0 _0766_
rlabel metal2 33208 16240 33208 16240 0 _0767_
rlabel metal2 32984 15484 32984 15484 0 _0768_
rlabel metal2 30632 9800 30632 9800 0 _0769_
rlabel metal2 32424 12096 32424 12096 0 _0770_
rlabel metal2 34440 8960 34440 8960 0 _0771_
rlabel metal2 34328 7448 34328 7448 0 _0772_
rlabel metal2 41160 16968 41160 16968 0 _0773_
rlabel metal2 38696 17136 38696 17136 0 _0774_
rlabel metal3 39312 16856 39312 16856 0 _0775_
rlabel metal2 26600 42448 26600 42448 0 _0776_
rlabel metal3 40880 16744 40880 16744 0 _0777_
rlabel metal3 21448 43960 21448 43960 0 _0778_
rlabel metal3 44492 16184 44492 16184 0 _0779_
rlabel metal2 22008 43960 22008 43960 0 _0780_
rlabel metal2 44856 16464 44856 16464 0 _0781_
rlabel metal2 29456 25704 29456 25704 0 _0782_
rlabel metal2 31528 22456 31528 22456 0 _0783_
rlabel metal2 33096 20048 33096 20048 0 _0784_
rlabel metal2 31864 20048 31864 20048 0 _0785_
rlabel metal2 33432 20832 33432 20832 0 _0786_
rlabel metal2 31752 19264 31752 19264 0 _0787_
rlabel metal3 35056 19880 35056 19880 0 _0788_
rlabel metal2 33432 18200 33432 18200 0 _0789_
rlabel metal2 16408 29904 16408 29904 0 _0790_
rlabel metal2 33488 30968 33488 30968 0 _0791_
rlabel metal2 32032 25480 32032 25480 0 _0792_
rlabel metal2 34104 32256 34104 32256 0 _0793_
rlabel metal2 33544 29960 33544 29960 0 _0794_
rlabel metal2 33152 27160 33152 27160 0 _0795_
rlabel metal2 18760 25648 18760 25648 0 _0796_
rlabel metal3 30968 25592 30968 25592 0 _0797_
rlabel metal3 25032 25368 25032 25368 0 _0798_
rlabel metal2 32200 25816 32200 25816 0 _0799_
rlabel metal2 20216 28336 20216 28336 0 _0800_
rlabel metal3 34608 29624 34608 29624 0 _0801_
rlabel metal2 41048 28784 41048 28784 0 _0802_
rlabel metal2 40600 28280 40600 28280 0 _0803_
rlabel metal2 40040 29568 40040 29568 0 _0804_
rlabel metal3 43344 28728 43344 28728 0 _0805_
rlabel metal2 42616 28616 42616 28616 0 _0806_
rlabel metal2 40936 29792 40936 29792 0 _0807_
rlabel metal2 25592 5544 25592 5544 0 _0808_
rlabel metal2 24640 7448 24640 7448 0 _0809_
rlabel metal2 26824 5936 26824 5936 0 _0810_
rlabel metal2 20776 20384 20776 20384 0 _0811_
rlabel metal2 25648 8232 25648 8232 0 _0812_
rlabel metal3 25200 7448 25200 7448 0 _0813_
rlabel metal2 28392 7448 28392 7448 0 _0814_
rlabel metal2 30072 5936 30072 5936 0 _0815_
rlabel metal3 28896 8120 28896 8120 0 _0816_
rlabel metal2 3304 14560 3304 14560 0 _0817_
rlabel metal2 3976 14168 3976 14168 0 _0818_
rlabel metal2 3472 8008 3472 8008 0 _0819_
rlabel metal3 3528 12824 3528 12824 0 _0820_
rlabel metal3 3696 8120 3696 8120 0 _0821_
rlabel metal3 3864 6776 3864 6776 0 _0822_
rlabel metal3 3416 8344 3416 8344 0 _0823_
rlabel metal2 5152 6664 5152 6664 0 _0824_
rlabel metal3 3976 7560 3976 7560 0 _0825_
rlabel metal3 5208 5656 5208 5656 0 _0826_
rlabel metal2 7224 6328 7224 6328 0 _0827_
rlabel metal3 5320 6776 5320 6776 0 _0828_
rlabel metal2 7896 6328 7896 6328 0 _0829_
rlabel metal2 7112 6664 7112 6664 0 _0830_
rlabel metal2 7784 4648 7784 4648 0 _0831_
rlabel metal3 5656 5096 5656 5096 0 _0832_
rlabel metal2 7448 4704 7448 4704 0 _0833_
rlabel metal2 8120 5880 8120 5880 0 _0834_
rlabel metal2 28168 28672 28168 28672 0 _0835_
rlabel metal2 25816 22624 25816 22624 0 _0836_
rlabel metal2 22232 24528 22232 24528 0 _0837_
rlabel metal2 20104 25536 20104 25536 0 _0838_
rlabel metal2 21448 25872 21448 25872 0 _0839_
rlabel metal3 21616 25480 21616 25480 0 _0840_
rlabel metal2 19656 25480 19656 25480 0 _0841_
rlabel metal2 21728 33544 21728 33544 0 _0842_
rlabel metal2 17976 32480 17976 32480 0 _0843_
rlabel metal3 22624 33544 22624 33544 0 _0844_
rlabel metal3 17528 32536 17528 32536 0 _0845_
rlabel metal3 16800 29624 16800 29624 0 _0846_
rlabel metal2 15568 32536 15568 32536 0 _0847_
rlabel metal2 18312 33376 18312 33376 0 _0848_
rlabel metal2 19432 30520 19432 30520 0 _0849_
rlabel metal3 22624 44072 22624 44072 0 _0850_
rlabel metal3 22288 44296 22288 44296 0 _0851_
rlabel metal2 23240 39256 23240 39256 0 _0852_
rlabel metal2 26488 42896 26488 42896 0 _0853_
rlabel metal2 23352 44408 23352 44408 0 _0854_
rlabel metal3 21056 44184 21056 44184 0 _0855_
rlabel metal2 14168 14784 14168 14784 0 _0856_
rlabel metal2 23912 18256 23912 18256 0 _0857_
rlabel metal2 26376 5936 26376 5936 0 _0858_
rlabel metal2 23800 4368 23800 4368 0 _0859_
rlabel metal2 7000 14168 7000 14168 0 _0860_
rlabel metal2 26208 25480 26208 25480 0 _0861_
rlabel metal2 18984 25592 18984 25592 0 _0862_
rlabel metal2 25816 24024 25816 24024 0 _0863_
rlabel metal2 25256 25200 25256 25200 0 _0864_
rlabel metal3 18144 27720 18144 27720 0 _0865_
rlabel metal2 16856 25032 16856 25032 0 _0866_
rlabel metal2 24136 25032 24136 25032 0 _0867_
rlabel metal2 17976 28336 17976 28336 0 _0868_
rlabel metal2 27384 23688 27384 23688 0 _0869_
rlabel metal3 25256 23352 25256 23352 0 _0870_
rlabel metal2 38360 31472 38360 31472 0 _0871_
rlabel metal3 36456 31752 36456 31752 0 _0872_
rlabel metal2 41832 32704 41832 32704 0 _0873_
rlabel metal2 36120 32088 36120 32088 0 _0874_
rlabel metal3 39032 37464 39032 37464 0 _0875_
rlabel metal2 40936 35896 40936 35896 0 _0876_
rlabel metal2 35560 34552 35560 34552 0 _0877_
rlabel metal2 39592 37520 39592 37520 0 _0878_
rlabel metal2 35616 35112 35616 35112 0 _0879_
rlabel metal2 39368 37800 39368 37800 0 _0880_
rlabel metal2 39816 33824 39816 33824 0 _0881_
rlabel metal2 38976 34216 38976 34216 0 _0882_
rlabel metal2 37912 32032 37912 32032 0 _0883_
rlabel via2 40936 24584 40936 24584 0 _0884_
rlabel metal3 44296 34328 44296 34328 0 _0885_
rlabel metal3 42224 35112 42224 35112 0 _0886_
rlabel metal2 45640 34328 45640 34328 0 _0887_
rlabel metal2 44744 33544 44744 33544 0 _0888_
rlabel metal2 45416 34552 45416 34552 0 _0889_
rlabel metal2 42168 33768 42168 33768 0 _0890_
rlabel metal3 17808 29176 17808 29176 0 _0891_
rlabel metal2 2968 34440 2968 34440 0 _0892_
rlabel metal3 7112 37464 7112 37464 0 _0893_
rlabel metal2 7000 36064 7000 36064 0 _0894_
rlabel metal2 8792 35000 8792 35000 0 _0895_
rlabel metal2 10024 34552 10024 34552 0 _0896_
rlabel metal2 6552 35392 6552 35392 0 _0897_
rlabel metal2 2632 34104 2632 34104 0 _0898_
rlabel metal2 32760 40936 32760 40936 0 _0899_
rlabel metal2 4536 39032 4536 39032 0 _0900_
rlabel metal2 1960 34216 1960 34216 0 _0901_
rlabel metal3 8232 37016 8232 37016 0 _0902_
rlabel metal3 2856 36400 2856 36400 0 _0903_
rlabel metal2 3080 35728 3080 35728 0 _0904_
rlabel metal2 3192 35504 3192 35504 0 _0905_
rlabel metal3 3192 38920 3192 38920 0 _0906_
rlabel metal2 4368 38248 4368 38248 0 _0907_
rlabel metal2 3976 38752 3976 38752 0 _0908_
rlabel metal2 3640 37016 3640 37016 0 _0909_
rlabel metal2 6328 35168 6328 35168 0 _0910_
rlabel metal3 6440 35560 6440 35560 0 _0911_
rlabel metal2 35224 39424 35224 39424 0 _0912_
rlabel metal2 33432 42672 33432 42672 0 _0913_
rlabel metal4 33992 38920 33992 38920 0 _0914_
rlabel metal3 34832 38808 34832 38808 0 _0915_
rlabel metal2 35112 39088 35112 39088 0 _0916_
rlabel metal3 33264 39704 33264 39704 0 _0917_
rlabel metal2 32256 40600 32256 40600 0 _0918_
rlabel metal4 30744 40768 30744 40768 0 _0919_
rlabel metal2 31864 40656 31864 40656 0 _0920_
rlabel metal2 32536 39648 32536 39648 0 _0921_
rlabel metal2 29512 43904 29512 43904 0 _0922_
rlabel metal2 29456 35112 29456 35112 0 _0923_
rlabel metal2 29904 38024 29904 38024 0 _0924_
rlabel metal2 30296 39872 30296 39872 0 _0925_
rlabel metal2 29680 39704 29680 39704 0 _0926_
rlabel metal2 30296 37576 30296 37576 0 _0927_
rlabel metal2 30632 39060 30632 39060 0 _0928_
rlabel metal2 25928 38724 25928 38724 0 _0929_
rlabel metal3 28728 37912 28728 37912 0 _0930_
rlabel metal2 29400 39368 29400 39368 0 _0931_
rlabel metal2 31136 40376 31136 40376 0 _0932_
rlabel metal2 30632 40656 30632 40656 0 _0933_
rlabel metal2 32312 39536 32312 39536 0 _0934_
rlabel metal2 32760 39536 32760 39536 0 _0935_
rlabel metal3 34440 39592 34440 39592 0 _0936_
rlabel metal2 36120 38696 36120 38696 0 _0937_
rlabel metal2 44968 43960 44968 43960 0 _0938_
rlabel metal2 42952 36736 42952 36736 0 _0939_
rlabel metal3 40880 35448 40880 35448 0 _0940_
rlabel metal2 39032 35336 39032 35336 0 _0941_
rlabel metal2 40264 38864 40264 38864 0 _0942_
rlabel metal2 39648 38696 39648 38696 0 _0943_
rlabel metal2 39984 38696 39984 38696 0 _0944_
rlabel metal2 39480 36792 39480 36792 0 _0945_
rlabel metal2 40264 35728 40264 35728 0 _0946_
rlabel metal2 45864 40600 45864 40600 0 _0947_
rlabel metal2 44744 40712 44744 40712 0 _0948_
rlabel metal2 45080 39312 45080 39312 0 _0949_
rlabel metal3 45136 36232 45136 36232 0 _0950_
rlabel metal2 46032 33544 46032 33544 0 _0951_
rlabel metal2 43960 39480 43960 39480 0 _0952_
rlabel metal2 43176 39592 43176 39592 0 _0953_
rlabel metal2 42728 36008 42728 36008 0 _0954_
rlabel metal2 39592 36008 39592 36008 0 _0955_
rlabel metal2 34328 39144 34328 39144 0 _0956_
rlabel metal2 35728 37912 35728 37912 0 _0957_
rlabel metal2 39256 37912 39256 37912 0 _0958_
rlabel metal2 41832 36064 41832 36064 0 _0959_
rlabel metal3 43400 36344 43400 36344 0 _0960_
rlabel metal2 45192 36736 45192 36736 0 _0961_
rlabel metal3 41804 38136 41804 38136 0 _0962_
rlabel metal3 33936 38024 33936 38024 0 _0963_
rlabel metal2 30744 39088 30744 39088 0 _0964_
rlabel metal2 27608 39984 27608 39984 0 _0965_
rlabel metal2 27272 38528 27272 38528 0 _0966_
rlabel metal2 27384 39144 27384 39144 0 _0967_
rlabel metal3 34272 38808 34272 38808 0 _0968_
rlabel metal3 31584 38808 31584 38808 0 _0969_
rlabel metal3 32424 39032 32424 39032 0 _0970_
rlabel metal2 30968 39312 30968 39312 0 _0971_
rlabel metal2 31416 37240 31416 37240 0 _0972_
rlabel metal2 31416 37744 31416 37744 0 _0973_
rlabel metal2 43736 43960 43736 43960 0 _0974_
rlabel metal2 25480 37072 25480 37072 0 _0975_
rlabel metal2 26096 37240 26096 37240 0 _0976_
rlabel metal2 25368 36232 25368 36232 0 _0977_
rlabel metal2 26712 36512 26712 36512 0 _0978_
rlabel metal2 25816 35560 25816 35560 0 _0979_
rlabel metal3 32928 16856 32928 16856 0 _0980_
rlabel metal2 31696 26936 31696 26936 0 _0981_
rlabel metal2 7784 39088 7784 39088 0 _0982_
rlabel metal2 8680 39200 8680 39200 0 _0983_
rlabel metal3 6888 38808 6888 38808 0 _0984_
rlabel metal2 8232 39592 8232 39592 0 _0985_
rlabel metal2 36120 22064 36120 22064 0 _0986_
rlabel metal3 24808 38696 24808 38696 0 _0987_
rlabel metal2 36344 41216 36344 41216 0 _0988_
rlabel metal2 38920 40656 38920 40656 0 _0989_
rlabel metal3 34328 14504 34328 14504 0 _0990_
rlabel metal3 26544 39032 26544 39032 0 _0991_
rlabel metal2 24360 39592 24360 39592 0 _0992_
rlabel metal2 28560 40152 28560 40152 0 _0993_
rlabel metal2 29736 40600 29736 40600 0 _0994_
rlabel metal2 30072 43288 30072 43288 0 _0995_
rlabel metal2 32200 41720 32200 41720 0 _0996_
rlabel metal3 30576 41944 30576 41944 0 _0997_
rlabel metal2 30744 43848 30744 43848 0 _0998_
rlabel metal2 31752 44016 31752 44016 0 _0999_
rlabel metal2 31864 43848 31864 43848 0 _1000_
rlabel metal2 32536 43680 32536 43680 0 _1001_
rlabel metal2 33208 42448 33208 42448 0 _1002_
rlabel metal2 41160 43120 41160 43120 0 _1003_
rlabel metal2 39480 43288 39480 43288 0 _1004_
rlabel metal2 33600 41384 33600 41384 0 _1005_
rlabel metal2 44968 41776 44968 41776 0 _1006_
rlabel metal2 37184 39368 37184 39368 0 _1007_
rlabel metal2 35448 42952 35448 42952 0 _1008_
rlabel metal2 38696 39872 38696 39872 0 _1009_
rlabel metal3 38724 39480 38724 39480 0 _1010_
rlabel metal2 40376 39592 40376 39592 0 _1011_
rlabel metal2 38024 43064 38024 43064 0 _1012_
rlabel metal2 40712 40040 40712 40040 0 _1013_
rlabel metal2 37296 39816 37296 39816 0 _1014_
rlabel metal2 39144 41552 39144 41552 0 _1015_
rlabel metal2 39984 39032 39984 39032 0 _1016_
rlabel metal2 44184 40712 44184 40712 0 _1017_
rlabel metal3 43400 44072 43400 44072 0 _1018_
rlabel metal2 39144 43232 39144 43232 0 _1019_
rlabel metal2 43960 41048 43960 41048 0 _1020_
rlabel metal3 45472 42280 45472 42280 0 _1021_
rlabel metal2 43960 41328 43960 41328 0 _1022_
rlabel metal2 45192 41160 45192 41160 0 _1023_
rlabel metal3 18312 17080 18312 17080 0 clknet_0_wb_clk_i
rlabel metal3 13608 12936 13608 12936 0 clknet_2_0__leaf_wb_clk_i
rlabel metal3 17248 43736 17248 43736 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 44968 18032 44968 18032 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 39928 26544 39928 26544 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 7112 14392 7112 14392 0 clknet_leaf_0_wb_clk_i
rlabel metal2 14168 43512 14168 43512 0 clknet_leaf_10_wb_clk_i
rlabel metal2 21952 39592 21952 39592 0 clknet_leaf_11_wb_clk_i
rlabel metal3 18648 34888 18648 34888 0 clknet_leaf_12_wb_clk_i
rlabel metal2 16856 33040 16856 33040 0 clknet_leaf_13_wb_clk_i
rlabel metal3 22288 26824 22288 26824 0 clknet_leaf_14_wb_clk_i
rlabel metal2 25144 35112 25144 35112 0 clknet_leaf_15_wb_clk_i
rlabel metal2 25032 43988 25032 43988 0 clknet_leaf_16_wb_clk_i
rlabel metal2 36008 40376 36008 40376 0 clknet_leaf_17_wb_clk_i
rlabel metal2 40152 44072 40152 44072 0 clknet_leaf_18_wb_clk_i
rlabel metal2 44072 38808 44072 38808 0 clknet_leaf_19_wb_clk_i
rlabel metal2 1848 22344 1848 22344 0 clknet_leaf_1_wb_clk_i
rlabel metal2 40488 33768 40488 33768 0 clknet_leaf_20_wb_clk_i
rlabel metal2 43848 30016 43848 30016 0 clknet_leaf_21_wb_clk_i
rlabel metal2 42056 23576 42056 23576 0 clknet_leaf_22_wb_clk_i
rlabel metal2 33320 27832 33320 27832 0 clknet_leaf_23_wb_clk_i
rlabel metal3 34216 22232 34216 22232 0 clknet_leaf_24_wb_clk_i
rlabel metal2 37464 16464 37464 16464 0 clknet_leaf_25_wb_clk_i
rlabel metal2 44296 21168 44296 21168 0 clknet_leaf_26_wb_clk_i
rlabel metal2 40880 16072 40880 16072 0 clknet_leaf_27_wb_clk_i
rlabel metal2 46088 9800 46088 9800 0 clknet_leaf_28_wb_clk_i
rlabel metal3 31472 6664 31472 6664 0 clknet_leaf_29_wb_clk_i
rlabel metal2 15288 20440 15288 20440 0 clknet_leaf_2_wb_clk_i
rlabel metal2 25256 4480 25256 4480 0 clknet_leaf_30_wb_clk_i
rlabel metal2 25368 10304 25368 10304 0 clknet_leaf_31_wb_clk_i
rlabel metal2 32200 15232 32200 15232 0 clknet_leaf_32_wb_clk_i
rlabel metal2 20552 20048 20552 20048 0 clknet_leaf_33_wb_clk_i
rlabel metal2 23016 13608 23016 13608 0 clknet_leaf_34_wb_clk_i
rlabel metal2 21672 6328 21672 6328 0 clknet_leaf_35_wb_clk_i
rlabel metal2 13160 7112 13160 7112 0 clknet_leaf_36_wb_clk_i
rlabel metal3 8316 6664 8316 6664 0 clknet_leaf_37_wb_clk_i
rlabel metal2 4536 7840 4536 7840 0 clknet_leaf_38_wb_clk_i
rlabel metal2 22344 23464 22344 23464 0 clknet_leaf_3_wb_clk_i
rlabel metal2 15512 27440 15512 27440 0 clknet_leaf_4_wb_clk_i
rlabel metal2 11032 25032 11032 25032 0 clknet_leaf_5_wb_clk_i
rlabel metal2 1848 28168 1848 28168 0 clknet_leaf_6_wb_clk_i
rlabel metal3 9352 35560 9352 35560 0 clknet_leaf_7_wb_clk_i
rlabel metal2 1848 37632 1848 37632 0 clknet_leaf_8_wb_clk_i
rlabel metal2 6104 40768 6104 40768 0 clknet_leaf_9_wb_clk_i
rlabel metal2 45976 21448 45976 21448 0 custom_settings[0]
rlabel metal3 45122 45080 45122 45080 0 custom_settings[1]
rlabel metal3 45346 2744 45346 2744 0 io_in_1[0]
rlabel metal3 47194 7448 47194 7448 0 io_in_1[1]
rlabel metal2 46088 12712 46088 12712 0 io_in_1[2]
rlabel metal2 46256 17528 46256 17528 0 io_in_1[3]
rlabel metal2 46256 22232 46256 22232 0 io_in_1[4]
rlabel metal2 45920 24024 45920 24024 0 io_in_1[5]
rlabel metal2 45808 25928 45808 25928 0 io_in_1[6]
rlabel metal2 41552 24024 41552 24024 0 io_in_1[7]
rlabel metal2 29960 44296 29960 44296 0 io_in_2[0]
rlabel metal2 45976 43848 45976 43848 0 io_in_2[1]
rlabel metal2 18424 2058 18424 2058 0 io_out[10]
rlabel metal2 20216 3136 20216 3136 0 io_out[11]
rlabel metal3 31584 3416 31584 3416 0 io_out[17]
rlabel metal3 33992 3640 33992 3640 0 io_out[18]
rlabel metal2 32368 4200 32368 4200 0 io_out[19]
rlabel metal2 44632 3920 44632 3920 0 io_out[20]
rlabel metal2 35672 854 35672 854 0 io_out[21]
rlabel metal2 15288 2058 15288 2058 0 io_out[8]
rlabel metal2 16856 854 16856 854 0 io_out[9]
rlabel metal2 45640 39312 45640 39312 0 net1
rlabel metal2 42504 33040 42504 33040 0 net10
rlabel metal2 24304 33208 24304 33208 0 net11
rlabel metal3 45640 44016 45640 44016 0 net12
rlabel metal2 18760 43988 18760 43988 0 net13
rlabel metal2 16072 3584 16072 3584 0 net14
rlabel metal2 16072 7056 16072 7056 0 net15
rlabel metal2 24136 3864 24136 3864 0 net16
rlabel metal2 31416 3976 31416 3976 0 net17
rlabel metal2 31584 3640 31584 3640 0 net18
rlabel metal2 22064 17416 22064 17416 0 net19
rlabel metal3 41104 44072 41104 44072 0 net2
rlabel metal2 22568 16072 22568 16072 0 net20
rlabel metal2 15568 11704 15568 11704 0 net21
rlabel metal2 11032 7112 11032 7112 0 net22
rlabel metal2 2744 2030 2744 2030 0 net23
rlabel metal2 4312 2030 4312 2030 0 net24
rlabel metal2 5880 2030 5880 2030 0 net25
rlabel metal2 7448 2030 7448 2030 0 net26
rlabel metal2 9016 854 9016 854 0 net27
rlabel metal2 10584 2814 10584 2814 0 net28
rlabel metal2 12152 2590 12152 2590 0 net29
rlabel metal3 45864 9464 45864 9464 0 net3
rlabel metal2 13720 2086 13720 2086 0 net30
rlabel metal3 23016 4424 23016 4424 0 net31
rlabel metal2 23128 2030 23128 2030 0 net32
rlabel metal2 24696 2030 24696 2030 0 net33
rlabel metal2 26264 2030 26264 2030 0 net34
rlabel metal2 26040 3360 26040 3360 0 net35
rlabel metal2 42336 12264 42336 12264 0 net36
rlabel metal2 40376 2310 40376 2310 0 net37
rlabel metal3 43904 4872 43904 4872 0 net38
rlabel metal2 43512 1582 43512 1582 0 net39
rlabel metal2 45864 10920 45864 10920 0 net4
rlabel metal2 45080 854 45080 854 0 net40
rlabel metal3 35448 6440 35448 6440 0 net41
rlabel metal2 45864 12992 45864 12992 0 net5
rlabel metal3 42252 17416 42252 17416 0 net6
rlabel metal2 46144 23800 46144 23800 0 net7
rlabel metal2 45080 23016 45080 23016 0 net8
rlabel metal2 43064 30744 43064 30744 0 net9
rlabel metal2 18200 44744 18200 44744 0 rst_n
rlabel metal2 24696 30968 24696 30968 0 tt_um_rejunity_ay8913.active
rlabel metal2 21336 26208 21336 26208 0 tt_um_rejunity_ay8913.amplitude_A\[0\]
rlabel metal2 20440 22288 20440 22288 0 tt_um_rejunity_ay8913.amplitude_B\[0\]
rlabel metal2 23352 19936 23352 19936 0 tt_um_rejunity_ay8913.amplitude_C\[0\]
rlabel metal2 13608 27440 13608 27440 0 tt_um_rejunity_ay8913.clk_counter\[0\]
rlabel metal2 13832 27832 13832 27832 0 tt_um_rejunity_ay8913.clk_counter\[1\]
rlabel metal2 13720 26152 13720 26152 0 tt_um_rejunity_ay8913.clk_counter\[2\]
rlabel metal2 14056 23520 14056 23520 0 tt_um_rejunity_ay8913.clk_counter\[3\]
rlabel metal2 13720 22400 13720 22400 0 tt_um_rejunity_ay8913.clk_counter\[4\]
rlabel metal2 15736 21672 15736 21672 0 tt_um_rejunity_ay8913.clk_counter\[5\]
rlabel metal2 14504 19488 14504 19488 0 tt_um_rejunity_ay8913.clk_counter\[6\]
rlabel metal2 19320 26152 19320 26152 0 tt_um_rejunity_ay8913.envelope_A
rlabel metal2 19096 23464 19096 23464 0 tt_um_rejunity_ay8913.envelope_B
rlabel metal2 19208 21952 19208 21952 0 tt_um_rejunity_ay8913.envelope_C
rlabel metal2 11592 32480 11592 32480 0 tt_um_rejunity_ay8913.envelope_alternate
rlabel metal2 9688 34608 9688 34608 0 tt_um_rejunity_ay8913.envelope_attack
rlabel metal2 10360 30856 10360 30856 0 tt_um_rejunity_ay8913.envelope_continue
rlabel metal2 5320 33880 5320 33880 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[0\]
rlabel metal2 4312 34720 4312 34720 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[1\]
rlabel metal2 4648 39424 4648 39424 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[2\]
rlabel metal2 3976 36008 3976 36008 0 tt_um_rejunity_ay8913.envelope_generator.envelope_counter\[3\]
rlabel metal2 11928 33264 11928 33264 0 tt_um_rejunity_ay8913.envelope_generator.hold
rlabel metal2 8568 32928 8568 32928 0 tt_um_rejunity_ay8913.envelope_generator.invert_output
rlabel metal3 28392 38696 28392 38696 0 tt_um_rejunity_ay8913.envelope_generator.period\[0\]
rlabel metal2 38136 37296 38136 37296 0 tt_um_rejunity_ay8913.envelope_generator.period\[10\]
rlabel metal2 40376 34888 40376 34888 0 tt_um_rejunity_ay8913.envelope_generator.period\[11\]
rlabel metal2 42168 35728 42168 35728 0 tt_um_rejunity_ay8913.envelope_generator.period\[12\]
rlabel metal2 43848 34552 43848 34552 0 tt_um_rejunity_ay8913.envelope_generator.period\[13\]
rlabel metal2 45864 38920 45864 38920 0 tt_um_rejunity_ay8913.envelope_generator.period\[14\]
rlabel metal3 45864 38808 45864 38808 0 tt_um_rejunity_ay8913.envelope_generator.period\[15\]
rlabel metal2 28728 41048 28728 41048 0 tt_um_rejunity_ay8913.envelope_generator.period\[1\]
rlabel metal2 30408 36344 30408 36344 0 tt_um_rejunity_ay8913.envelope_generator.period\[2\]
rlabel metal2 29288 34048 29288 34048 0 tt_um_rejunity_ay8913.envelope_generator.period\[3\]
rlabel metal2 31080 32592 31080 32592 0 tt_um_rejunity_ay8913.envelope_generator.period\[4\]
rlabel metal2 33320 40376 33320 40376 0 tt_um_rejunity_ay8913.envelope_generator.period\[5\]
rlabel metal2 33208 38668 33208 38668 0 tt_um_rejunity_ay8913.envelope_generator.period\[6\]
rlabel metal3 34832 39144 34832 39144 0 tt_um_rejunity_ay8913.envelope_generator.period\[7\]
rlabel metal2 37912 33936 37912 33936 0 tt_um_rejunity_ay8913.envelope_generator.period\[8\]
rlabel metal2 38696 34384 38696 34384 0 tt_um_rejunity_ay8913.envelope_generator.period\[9\]
rlabel metal2 8680 36680 8680 36680 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.previous_signal_state_0
rlabel metal2 7896 39032 7896 39032 0 tt_um_rejunity_ay8913.envelope_generator.signal_edge.signal
rlabel metal3 8120 35672 8120 35672 0 tt_um_rejunity_ay8913.envelope_generator.stop
rlabel metal2 24640 39704 24640 39704 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[0\]
rlabel metal2 39816 38192 39816 38192 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[10\]
rlabel metal2 44520 43736 44520 43736 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[11\]
rlabel metal2 45192 44352 45192 44352 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[12\]
rlabel metal3 44968 41944 44968 41944 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[13\]
rlabel metal2 44184 43988 44184 43988 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[14\]
rlabel metal2 41384 39648 41384 39648 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[15\]
rlabel metal2 24696 39032 24696 39032 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[1\]
rlabel metal3 29232 41272 29232 41272 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[2\]
rlabel metal2 29176 43680 29176 43680 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[3\]
rlabel metal2 29512 42952 29512 42952 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[4\]
rlabel metal2 33040 43400 33040 43400 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[5\]
rlabel metal2 35056 41272 35056 41272 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[6\]
rlabel metal3 39592 43960 39592 43960 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[7\]
rlabel metal2 43848 39984 43848 39984 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[8\]
rlabel metal2 38696 38668 38696 38668 0 tt_um_rejunity_ay8913.envelope_generator.tone.counter\[9\]
rlabel metal2 24864 28728 24864 28728 0 tt_um_rejunity_ay8913.latched_register\[0\]
rlabel metal2 28448 26488 28448 26488 0 tt_um_rejunity_ay8913.latched_register\[1\]
rlabel metal2 29624 29400 29624 29400 0 tt_um_rejunity_ay8913.latched_register\[2\]
rlabel metal2 32480 30968 32480 30968 0 tt_um_rejunity_ay8913.latched_register\[3\]
rlabel metal2 20664 28112 20664 28112 0 tt_um_rejunity_ay8913.noise_disable_A
rlabel metal2 26712 23352 26712 23352 0 tt_um_rejunity_ay8913.noise_disable_B
rlabel metal3 24640 23128 24640 23128 0 tt_um_rejunity_ay8913.noise_disable_C
rlabel metal2 21168 26376 21168 26376 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[0\]
rlabel metal2 3248 27944 3248 27944 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[10\]
rlabel metal2 2016 29512 2016 29512 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[11\]
rlabel metal2 3192 29960 3192 29960 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[12\]
rlabel metal2 6552 30408 6552 30408 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[13\]
rlabel metal3 7112 30296 7112 30296 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[14\]
rlabel metal2 7448 29120 7448 29120 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[15\]
rlabel metal2 8568 25704 8568 25704 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[16\]
rlabel metal3 7672 24024 7672 24024 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[1\]
rlabel metal2 8456 22512 8456 22512 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[2\]
rlabel metal2 8120 23296 8120 23296 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[3\]
rlabel metal2 5992 22344 5992 22344 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[4\]
rlabel metal2 2856 18424 2856 18424 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[5\]
rlabel metal2 4088 21448 4088 21448 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[6\]
rlabel metal2 2856 21504 2856 21504 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[7\]
rlabel metal3 2520 24920 2520 24920 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[8\]
rlabel metal3 3920 26488 3920 26488 0 tt_um_rejunity_ay8913.noise_generator.lfsr\[9\]
rlabel metal2 28560 16184 28560 16184 0 tt_um_rejunity_ay8913.noise_generator.period\[0\]
rlabel metal2 29288 15064 29288 15064 0 tt_um_rejunity_ay8913.noise_generator.period\[1\]
rlabel metal2 29736 13104 29736 13104 0 tt_um_rejunity_ay8913.noise_generator.period\[2\]
rlabel metal2 28056 13216 28056 13216 0 tt_um_rejunity_ay8913.noise_generator.period\[3\]
rlabel metal2 27720 12600 27720 12600 0 tt_um_rejunity_ay8913.noise_generator.period\[4\]
rlabel metal2 8400 18312 8400 18312 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.previous_signal_state_0
rlabel metal2 8064 13944 8064 13944 0 tt_um_rejunity_ay8913.noise_generator.signal_edge.signal
rlabel metal2 26152 16520 26152 16520 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[0\]
rlabel metal2 26264 15204 26264 15204 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[1\]
rlabel metal2 26600 12600 26600 12600 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[2\]
rlabel metal2 24472 11200 24472 11200 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[3\]
rlabel metal2 28056 10472 28056 10472 0 tt_um_rejunity_ay8913.noise_generator.tone.counter\[4\]
rlabel metal3 14672 17640 14672 17640 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[2\]
rlabel metal2 12488 16464 12488 16464 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[3\]
rlabel metal2 8680 16240 8680 16240 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[4\]
rlabel metal2 10248 14840 10248 14840 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[5\]
rlabel metal3 10416 14504 10416 14504 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[6\]
rlabel metal3 12992 14504 12992 14504 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[7\]
rlabel metal2 12264 12600 12264 12600 0 tt_um_rejunity_ay8913.pwm_A.accumulator\[8\]
rlabel metal2 4480 15064 4480 15064 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[2\]
rlabel metal2 4648 13552 4648 13552 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[3\]
rlabel metal2 3696 8008 3696 8008 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[4\]
rlabel metal2 2856 7336 2856 7336 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[5\]
rlabel metal2 4984 6160 4984 6160 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[6\]
rlabel metal2 7224 5712 7224 5712 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[7\]
rlabel metal2 6328 5152 6328 5152 0 tt_um_rejunity_ay8913.pwm_B.accumulator\[8\]
rlabel metal2 18200 20832 18200 20832 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[2\]
rlabel metal2 16856 17528 16856 17528 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[3\]
rlabel metal2 5544 16576 5544 16576 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[4\]
rlabel metal3 5208 12936 5208 12936 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[5\]
rlabel metal3 6216 12152 6216 12152 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[6\]
rlabel metal2 6104 11424 6104 11424 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[7\]
rlabel metal2 8568 8372 8568 8372 0 tt_um_rejunity_ay8913.pwm_C.accumulator\[8\]
rlabel metal3 20384 16744 20384 16744 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[2\]
rlabel metal3 16912 15176 16912 15176 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[3\]
rlabel metal2 20328 11592 20328 11592 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[4\]
rlabel metal2 19208 12600 19208 12600 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[5\]
rlabel metal2 17752 10248 17752 10248 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[6\]
rlabel metal2 14896 10472 14896 10472 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[7\]
rlabel metal2 11592 10360 11592 10360 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[8\]
rlabel metal3 11816 8232 11816 8232 0 tt_um_rejunity_ay8913.pwm_master.accumulator\[9\]
rlabel metal2 12488 36792 12488 36792 0 tt_um_rejunity_ay8913.restart_envelope
rlabel metal2 26712 3584 26712 3584 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[0\]
rlabel metal2 25032 9072 25032 9072 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[1\]
rlabel metal2 26376 7896 26376 7896 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[2\]
rlabel metal2 29232 6776 29232 6776 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[3\]
rlabel metal2 29624 8288 29624 8288 0 tt_um_rejunity_ay8913.spi_dac_i_2.counter\[4\]
rlabel metal3 17528 5880 17528 5880 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 20888 4760 20888 4760 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 22904 5880 22904 5880 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 20664 9296 20664 9296 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 20328 8568 20328 8568 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 19656 7056 19656 7056 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 16968 5824 16968 5824 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal2 12936 5544 12936 5544 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal3 13664 6552 13664 6552 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 14728 5936 14728 5936 0 tt_um_rejunity_ay8913.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 18928 29288 18928 29288 0 tt_um_rejunity_ay8913.tone_A
rlabel metal2 16408 36288 16408 36288 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[0\]
rlabel metal3 10864 39368 10864 39368 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[10\]
rlabel metal2 12712 38752 12712 38752 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[11\]
rlabel metal2 16968 34944 16968 34944 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[1\]
rlabel metal2 16184 38808 16184 38808 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[2\]
rlabel metal2 15792 41048 15792 41048 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[3\]
rlabel metal2 18704 38696 18704 38696 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[4\]
rlabel metal3 16912 42056 16912 42056 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[5\]
rlabel metal2 12936 41944 12936 41944 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[6\]
rlabel metal2 13608 44576 13608 44576 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[7\]
rlabel metal2 24808 42672 24808 42672 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[8\]
rlabel metal4 20216 40488 20216 40488 0 tt_um_rejunity_ay8913.tone_A_generator.counter\[9\]
rlabel metal2 16968 30856 16968 30856 0 tt_um_rejunity_ay8913.tone_A_generator.period\[0\]
rlabel metal2 18760 39984 18760 39984 0 tt_um_rejunity_ay8913.tone_A_generator.period\[10\]
rlabel metal2 19040 39592 19040 39592 0 tt_um_rejunity_ay8913.tone_A_generator.period\[11\]
rlabel metal2 16744 32984 16744 32984 0 tt_um_rejunity_ay8913.tone_A_generator.period\[1\]
rlabel metal2 20328 38136 20328 38136 0 tt_um_rejunity_ay8913.tone_A_generator.period\[2\]
rlabel metal2 17416 31472 17416 31472 0 tt_um_rejunity_ay8913.tone_A_generator.period\[3\]
rlabel metal2 22904 38976 22904 38976 0 tt_um_rejunity_ay8913.tone_A_generator.period\[4\]
rlabel metal2 24696 41944 24696 41944 0 tt_um_rejunity_ay8913.tone_A_generator.period\[5\]
rlabel metal3 22120 43400 22120 43400 0 tt_um_rejunity_ay8913.tone_A_generator.period\[6\]
rlabel metal2 21560 43932 21560 43932 0 tt_um_rejunity_ay8913.tone_A_generator.period\[7\]
rlabel metal2 22512 40264 22512 40264 0 tt_um_rejunity_ay8913.tone_A_generator.period\[8\]
rlabel metal2 24696 35336 24696 35336 0 tt_um_rejunity_ay8913.tone_A_generator.period\[9\]
rlabel metal2 26600 21392 26600 21392 0 tt_um_rejunity_ay8913.tone_B
rlabel metal2 37240 23968 37240 23968 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[0\]
rlabel metal2 43848 18368 43848 18368 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[10\]
rlabel metal2 46200 16520 46200 16520 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[11\]
rlabel metal2 33992 23800 33992 23800 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[1\]
rlabel metal3 36568 26152 36568 26152 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[2\]
rlabel metal2 39256 27440 39256 27440 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[3\]
rlabel metal2 41048 27776 41048 27776 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[4\]
rlabel metal2 44296 25368 44296 25368 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[5\]
rlabel metal2 41496 24920 41496 24920 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[6\]
rlabel metal2 44184 23576 44184 23576 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[7\]
rlabel metal3 40880 20888 40880 20888 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[8\]
rlabel metal2 45976 19208 45976 19208 0 tt_um_rejunity_ay8913.tone_B_generator.counter\[9\]
rlabel metal2 36008 27776 36008 27776 0 tt_um_rejunity_ay8913.tone_B_generator.period\[0\]
rlabel metal2 39592 18872 39592 18872 0 tt_um_rejunity_ay8913.tone_B_generator.period\[10\]
rlabel metal2 38696 18480 38696 18480 0 tt_um_rejunity_ay8913.tone_B_generator.period\[11\]
rlabel metal3 32144 24584 32144 24584 0 tt_um_rejunity_ay8913.tone_B_generator.period\[1\]
rlabel metal2 37408 25704 37408 25704 0 tt_um_rejunity_ay8913.tone_B_generator.period\[2\]
rlabel metal2 38808 27216 38808 27216 0 tt_um_rejunity_ay8913.tone_B_generator.period\[3\]
rlabel metal3 40544 27048 40544 27048 0 tt_um_rejunity_ay8913.tone_B_generator.period\[4\]
rlabel metal2 46256 24024 46256 24024 0 tt_um_rejunity_ay8913.tone_B_generator.period\[5\]
rlabel metal2 46200 26040 46200 26040 0 tt_um_rejunity_ay8913.tone_B_generator.period\[6\]
rlabel metal2 42840 24360 42840 24360 0 tt_um_rejunity_ay8913.tone_B_generator.period\[7\]
rlabel metal2 39704 21168 39704 21168 0 tt_um_rejunity_ay8913.tone_B_generator.period\[8\]
rlabel metal2 38808 19656 38808 19656 0 tt_um_rejunity_ay8913.tone_B_generator.period\[9\]
rlabel metal2 26488 18872 26488 18872 0 tt_um_rejunity_ay8913.tone_C
rlabel metal2 36288 17640 36288 17640 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[0\]
rlabel metal2 39872 9240 39872 9240 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[10\]
rlabel metal3 35616 5208 35616 5208 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[11\]
rlabel metal2 37912 13664 37912 13664 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[1\]
rlabel metal2 38360 13832 38360 13832 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[2\]
rlabel metal2 38808 11088 38808 11088 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[3\]
rlabel metal2 41608 12264 41608 12264 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[4\]
rlabel metal2 40376 12488 40376 12488 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[5\]
rlabel metal2 42672 9800 42672 9800 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[6\]
rlabel metal2 43960 9016 43960 9016 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[7\]
rlabel metal2 40040 6328 40040 6328 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[8\]
rlabel metal2 39872 5208 39872 5208 0 tt_um_rejunity_ay8913.tone_C_generator.counter\[9\]
rlabel metal3 36120 10808 36120 10808 0 tt_um_rejunity_ay8913.tone_C_generator.period\[0\]
rlabel metal2 39256 4088 39256 4088 0 tt_um_rejunity_ay8913.tone_C_generator.period\[10\]
rlabel metal2 34776 4648 34776 4648 0 tt_um_rejunity_ay8913.tone_C_generator.period\[11\]
rlabel metal3 35112 12152 35112 12152 0 tt_um_rejunity_ay8913.tone_C_generator.period\[1\]
rlabel metal2 37464 10920 37464 10920 0 tt_um_rejunity_ay8913.tone_C_generator.period\[2\]
rlabel metal2 38136 11900 38136 11900 0 tt_um_rejunity_ay8913.tone_C_generator.period\[3\]
rlabel metal2 40376 16240 40376 16240 0 tt_um_rejunity_ay8913.tone_C_generator.period\[4\]
rlabel metal2 41832 16464 41832 16464 0 tt_um_rejunity_ay8913.tone_C_generator.period\[5\]
rlabel metal2 43736 16408 43736 16408 0 tt_um_rejunity_ay8913.tone_C_generator.period\[6\]
rlabel metal2 42952 16184 42952 16184 0 tt_um_rejunity_ay8913.tone_C_generator.period\[7\]
rlabel metal3 33264 7560 33264 7560 0 tt_um_rejunity_ay8913.tone_C_generator.period\[8\]
rlabel metal2 33824 5992 33824 5992 0 tt_um_rejunity_ay8913.tone_C_generator.period\[9\]
rlabel metal2 18424 27104 18424 27104 0 tt_um_rejunity_ay8913.tone_disable_A
rlabel metal2 18592 24024 18592 24024 0 tt_um_rejunity_ay8913.tone_disable_B
rlabel metal2 25144 23576 25144 23576 0 tt_um_rejunity_ay8913.tone_disable_C
rlabel metal2 6104 45486 6104 45486 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 48000 48000
<< end >>
