magic
tech gf180mcuD
magscale 1 5
timestamp 1699958466
<< obsm1 >>
rect 672 1538 29288 33417
<< metal2 >>
rect 1344 34600 1400 35000
rect 2352 34600 2408 35000
rect 3360 34600 3416 35000
rect 4368 34600 4424 35000
rect 5376 34600 5432 35000
rect 6384 34600 6440 35000
rect 7392 34600 7448 35000
rect 8400 34600 8456 35000
rect 9408 34600 9464 35000
rect 10416 34600 10472 35000
rect 11424 34600 11480 35000
rect 12432 34600 12488 35000
rect 13440 34600 13496 35000
rect 14448 34600 14504 35000
rect 15456 34600 15512 35000
rect 16464 34600 16520 35000
rect 17472 34600 17528 35000
rect 18480 34600 18536 35000
rect 19488 34600 19544 35000
rect 20496 34600 20552 35000
rect 21504 34600 21560 35000
rect 22512 34600 22568 35000
rect 23520 34600 23576 35000
rect 24528 34600 24584 35000
rect 25536 34600 25592 35000
rect 26544 34600 26600 35000
rect 27552 34600 27608 35000
rect 28560 34600 28616 35000
<< obsm2 >>
rect 854 34570 1314 34600
rect 1430 34570 2322 34600
rect 2438 34570 3330 34600
rect 3446 34570 4338 34600
rect 4454 34570 5346 34600
rect 5462 34570 6354 34600
rect 6470 34570 7362 34600
rect 7478 34570 8370 34600
rect 8486 34570 9378 34600
rect 9494 34570 10386 34600
rect 10502 34570 11394 34600
rect 11510 34570 12402 34600
rect 12518 34570 13410 34600
rect 13526 34570 14418 34600
rect 14534 34570 15426 34600
rect 15542 34570 16434 34600
rect 16550 34570 17442 34600
rect 17558 34570 18450 34600
rect 18566 34570 19458 34600
rect 19574 34570 20466 34600
rect 20582 34570 21474 34600
rect 21590 34570 22482 34600
rect 22598 34570 23490 34600
rect 23606 34570 24498 34600
rect 24614 34570 25506 34600
rect 25622 34570 26514 34600
rect 26630 34570 27522 34600
rect 27638 34570 28530 34600
rect 28646 34570 29162 34600
rect 854 1549 29162 34570
<< metal3 >>
rect 29600 33040 30000 33096
rect 29600 29568 30000 29624
rect 0 29120 400 29176
rect 29600 26096 30000 26152
rect 29600 22624 30000 22680
rect 29600 19152 30000 19208
rect 0 17472 400 17528
rect 29600 15680 30000 15736
rect 29600 12208 30000 12264
rect 29600 8736 30000 8792
rect 0 5824 400 5880
rect 29600 5264 30000 5320
rect 29600 1792 30000 1848
<< obsm3 >>
rect 400 33126 29600 33418
rect 400 33010 29570 33126
rect 400 29654 29600 33010
rect 400 29538 29570 29654
rect 400 29206 29600 29538
rect 430 29090 29600 29206
rect 400 26182 29600 29090
rect 400 26066 29570 26182
rect 400 22710 29600 26066
rect 400 22594 29570 22710
rect 400 19238 29600 22594
rect 400 19122 29570 19238
rect 400 17558 29600 19122
rect 430 17442 29600 17558
rect 400 15766 29600 17442
rect 400 15650 29570 15766
rect 400 12294 29600 15650
rect 400 12178 29570 12294
rect 400 8822 29600 12178
rect 400 8706 29570 8822
rect 400 5910 29600 8706
rect 430 5794 29600 5910
rect 400 5350 29600 5794
rect 400 5234 29570 5350
rect 400 1878 29600 5234
rect 400 1762 29570 1878
rect 400 1554 29600 1762
<< metal4 >>
rect 2224 1538 2384 33350
rect 9904 1538 10064 33350
rect 17584 1538 17744 33350
rect 25264 1538 25424 33350
<< obsm4 >>
rect 2142 2921 2194 31575
rect 2414 2921 9874 31575
rect 10094 2921 17554 31575
rect 17774 2921 25234 31575
rect 25454 2921 25746 31575
<< labels >>
rlabel metal3 s 29600 29568 30000 29624 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 29600 33040 30000 33096 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 29600 1792 30000 1848 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 29600 5264 30000 5320 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 29600 8736 30000 8792 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 29600 12208 30000 12264 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 29600 15680 30000 15736 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 29600 19152 30000 19208 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 29600 22624 30000 22680 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 29600 26096 30000 26152 6 io_in_1[7]
port 10 nsew signal input
rlabel metal3 s 0 29120 400 29176 6 io_in_2
port 11 nsew signal input
rlabel metal2 s 1344 34600 1400 35000 6 io_out[0]
port 12 nsew signal output
rlabel metal2 s 11424 34600 11480 35000 6 io_out[10]
port 13 nsew signal output
rlabel metal2 s 12432 34600 12488 35000 6 io_out[11]
port 14 nsew signal output
rlabel metal2 s 13440 34600 13496 35000 6 io_out[12]
port 15 nsew signal output
rlabel metal2 s 14448 34600 14504 35000 6 io_out[13]
port 16 nsew signal output
rlabel metal2 s 15456 34600 15512 35000 6 io_out[14]
port 17 nsew signal output
rlabel metal2 s 16464 34600 16520 35000 6 io_out[15]
port 18 nsew signal output
rlabel metal2 s 17472 34600 17528 35000 6 io_out[16]
port 19 nsew signal output
rlabel metal2 s 18480 34600 18536 35000 6 io_out[17]
port 20 nsew signal output
rlabel metal2 s 19488 34600 19544 35000 6 io_out[18]
port 21 nsew signal output
rlabel metal2 s 20496 34600 20552 35000 6 io_out[19]
port 22 nsew signal output
rlabel metal2 s 2352 34600 2408 35000 6 io_out[1]
port 23 nsew signal output
rlabel metal2 s 21504 34600 21560 35000 6 io_out[20]
port 24 nsew signal output
rlabel metal2 s 22512 34600 22568 35000 6 io_out[21]
port 25 nsew signal output
rlabel metal2 s 23520 34600 23576 35000 6 io_out[22]
port 26 nsew signal output
rlabel metal2 s 24528 34600 24584 35000 6 io_out[23]
port 27 nsew signal output
rlabel metal2 s 25536 34600 25592 35000 6 io_out[24]
port 28 nsew signal output
rlabel metal2 s 26544 34600 26600 35000 6 io_out[25]
port 29 nsew signal output
rlabel metal2 s 27552 34600 27608 35000 6 io_out[26]
port 30 nsew signal output
rlabel metal2 s 28560 34600 28616 35000 6 io_out[27]
port 31 nsew signal output
rlabel metal2 s 3360 34600 3416 35000 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 4368 34600 4424 35000 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 5376 34600 5432 35000 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 6384 34600 6440 35000 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 7392 34600 7448 35000 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 8400 34600 8456 35000 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 9408 34600 9464 35000 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 10416 34600 10472 35000 6 io_out[9]
port 39 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 rst_n
port 40 nsew signal input
rlabel metal4 s 2224 1538 2384 33350 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 33350 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 33350 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 33350 6 vss
port 42 nsew ground bidirectional
rlabel metal3 s 0 5824 400 5880 6 wb_clk_i
port 43 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 35000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2874506
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_sn76489/runs/23_11_14_11_37/results/signoff/wrapped_sn76489.magic.gds
string GDS_START 391704
<< end >>

