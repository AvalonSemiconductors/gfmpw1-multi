* NGSPICE file created from wrapped_sn76489.ext - technology: gf180mcuD

.subckt wrapped_sn76489 custom_settings[0] custom_settings[1] io_in_1[0] io_in_1[1]
+ io_in_1[2] io_in_1[3] io_in_1[4] io_in_1[5] io_in_1[6] io_in_1[7] io_in_2 io_out[0]
+ io_out[10] io_out[11] io_out[12] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] rst_n vdd vss wb_clk_i io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[4] io_out[3] io_out[2]
.ends

