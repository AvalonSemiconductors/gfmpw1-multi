VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_avalonsemi_tbb1143
  CLASS BLOCK ;
  FOREIGN tholin_avalonsemi_tbb1143 ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 230.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 13.440 230.000 14.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 47.040 230.000 47.600 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 63.840 230.000 64.400 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 80.640 230.000 81.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 97.440 230.000 98.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    ANTENNADIFFAREA 0.877000 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 114.240 230.000 114.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 131.040 230.000 131.600 ;
    END
  END io_in[5]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 147.840 230.000 148.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 164.640 230.000 165.200 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 181.440 230.000 182.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 198.240 230.000 198.800 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 215.040 230.000 215.600 ;
    END
  END io_out[4]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 226.000 30.240 230.000 30.800 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 209.910 223.310 212.110 ;
      LAYER Nwell ;
        RECT 6.290 205.610 223.310 209.910 ;
      LAYER Pwell ;
        RECT 6.290 202.070 223.310 205.610 ;
      LAYER Nwell ;
        RECT 6.290 197.770 223.310 202.070 ;
      LAYER Pwell ;
        RECT 6.290 194.230 223.310 197.770 ;
      LAYER Nwell ;
        RECT 6.290 189.930 223.310 194.230 ;
      LAYER Pwell ;
        RECT 6.290 186.390 223.310 189.930 ;
      LAYER Nwell ;
        RECT 6.290 182.090 223.310 186.390 ;
      LAYER Pwell ;
        RECT 6.290 178.550 223.310 182.090 ;
      LAYER Nwell ;
        RECT 6.290 174.250 223.310 178.550 ;
      LAYER Pwell ;
        RECT 6.290 170.710 223.310 174.250 ;
      LAYER Nwell ;
        RECT 6.290 166.410 223.310 170.710 ;
      LAYER Pwell ;
        RECT 6.290 162.870 223.310 166.410 ;
      LAYER Nwell ;
        RECT 6.290 158.570 223.310 162.870 ;
      LAYER Pwell ;
        RECT 6.290 155.030 223.310 158.570 ;
      LAYER Nwell ;
        RECT 6.290 150.730 223.310 155.030 ;
      LAYER Pwell ;
        RECT 6.290 147.190 223.310 150.730 ;
      LAYER Nwell ;
        RECT 6.290 142.890 223.310 147.190 ;
      LAYER Pwell ;
        RECT 6.290 139.350 223.310 142.890 ;
      LAYER Nwell ;
        RECT 6.290 135.050 223.310 139.350 ;
      LAYER Pwell ;
        RECT 6.290 131.510 223.310 135.050 ;
      LAYER Nwell ;
        RECT 6.290 127.210 223.310 131.510 ;
      LAYER Pwell ;
        RECT 6.290 123.670 223.310 127.210 ;
      LAYER Nwell ;
        RECT 6.290 119.370 223.310 123.670 ;
      LAYER Pwell ;
        RECT 6.290 115.830 223.310 119.370 ;
      LAYER Nwell ;
        RECT 6.290 111.530 223.310 115.830 ;
      LAYER Pwell ;
        RECT 6.290 107.990 223.310 111.530 ;
      LAYER Nwell ;
        RECT 6.290 103.690 223.310 107.990 ;
      LAYER Pwell ;
        RECT 6.290 100.150 223.310 103.690 ;
      LAYER Nwell ;
        RECT 6.290 95.850 223.310 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 223.310 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 223.310 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 223.310 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 223.310 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 223.310 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 223.310 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 223.310 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 223.310 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 223.310 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 223.310 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 223.310 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 223.310 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 223.310 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 223.310 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 223.310 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 223.310 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 223.310 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 223.310 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 223.310 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 223.310 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 223.310 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 222.880 211.980 ;
      LAYER Metal2 ;
        RECT 22.380 13.530 222.740 215.510 ;
      LAYER Metal3 ;
        RECT 22.330 214.740 225.700 215.460 ;
        RECT 22.330 199.100 226.000 214.740 ;
        RECT 22.330 197.940 225.700 199.100 ;
        RECT 22.330 182.300 226.000 197.940 ;
        RECT 22.330 181.140 225.700 182.300 ;
        RECT 22.330 165.500 226.000 181.140 ;
        RECT 22.330 164.340 225.700 165.500 ;
        RECT 22.330 148.700 226.000 164.340 ;
        RECT 22.330 147.540 225.700 148.700 ;
        RECT 22.330 131.900 226.000 147.540 ;
        RECT 22.330 130.740 225.700 131.900 ;
        RECT 22.330 115.100 226.000 130.740 ;
        RECT 22.330 113.940 225.700 115.100 ;
        RECT 22.330 98.300 226.000 113.940 ;
        RECT 22.330 97.140 225.700 98.300 ;
        RECT 22.330 81.500 226.000 97.140 ;
        RECT 22.330 80.340 225.700 81.500 ;
        RECT 22.330 64.700 226.000 80.340 ;
        RECT 22.330 63.540 225.700 64.700 ;
        RECT 22.330 47.900 226.000 63.540 ;
        RECT 22.330 46.740 225.700 47.900 ;
        RECT 22.330 31.100 226.000 46.740 ;
        RECT 22.330 29.940 225.700 31.100 ;
        RECT 22.330 14.300 226.000 29.940 ;
        RECT 22.330 13.580 225.700 14.300 ;
      LAYER Metal4 ;
        RECT 84.140 21.370 98.740 188.070 ;
        RECT 100.940 21.370 175.540 188.070 ;
        RECT 177.740 21.370 219.940 188.070 ;
  END
END tholin_avalonsemi_tbb1143
END LIBRARY

