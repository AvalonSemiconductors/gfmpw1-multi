VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO diceroll
  CLASS BLOCK ;
  FOREIGN diceroll ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 230.000 ;
  PIN io_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 226.000 47.600 230.000 ;
    END
  END io_in
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 226.000 66.640 230.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 226.000 85.680 230.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 226.000 104.720 230.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 226.000 123.760 230.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 226.000 142.800 230.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 226.000 161.840 230.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 226.000 180.880 230.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 226.000 199.920 230.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 226.000 218.960 230.000 ;
    END
  END io_out[8]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 226.000 28.560 230.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 226.000 9.520 230.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 209.910 223.310 212.110 ;
      LAYER Nwell ;
        RECT 6.290 205.610 223.310 209.910 ;
      LAYER Pwell ;
        RECT 6.290 202.070 223.310 205.610 ;
      LAYER Nwell ;
        RECT 6.290 197.770 223.310 202.070 ;
      LAYER Pwell ;
        RECT 6.290 194.230 223.310 197.770 ;
      LAYER Nwell ;
        RECT 6.290 189.930 223.310 194.230 ;
      LAYER Pwell ;
        RECT 6.290 186.390 223.310 189.930 ;
      LAYER Nwell ;
        RECT 6.290 182.090 223.310 186.390 ;
      LAYER Pwell ;
        RECT 6.290 178.550 223.310 182.090 ;
      LAYER Nwell ;
        RECT 6.290 174.250 223.310 178.550 ;
      LAYER Pwell ;
        RECT 6.290 170.710 223.310 174.250 ;
      LAYER Nwell ;
        RECT 6.290 166.410 223.310 170.710 ;
      LAYER Pwell ;
        RECT 6.290 162.870 223.310 166.410 ;
      LAYER Nwell ;
        RECT 6.290 158.570 223.310 162.870 ;
      LAYER Pwell ;
        RECT 6.290 155.030 223.310 158.570 ;
      LAYER Nwell ;
        RECT 6.290 150.730 223.310 155.030 ;
      LAYER Pwell ;
        RECT 6.290 147.190 223.310 150.730 ;
      LAYER Nwell ;
        RECT 6.290 142.890 223.310 147.190 ;
      LAYER Pwell ;
        RECT 6.290 139.350 223.310 142.890 ;
      LAYER Nwell ;
        RECT 6.290 135.050 223.310 139.350 ;
      LAYER Pwell ;
        RECT 6.290 131.510 223.310 135.050 ;
      LAYER Nwell ;
        RECT 6.290 127.210 223.310 131.510 ;
      LAYER Pwell ;
        RECT 6.290 123.670 223.310 127.210 ;
      LAYER Nwell ;
        RECT 6.290 119.370 223.310 123.670 ;
      LAYER Pwell ;
        RECT 6.290 115.830 223.310 119.370 ;
      LAYER Nwell ;
        RECT 6.290 111.530 223.310 115.830 ;
      LAYER Pwell ;
        RECT 6.290 107.990 223.310 111.530 ;
      LAYER Nwell ;
        RECT 6.290 103.690 223.310 107.990 ;
      LAYER Pwell ;
        RECT 6.290 100.150 223.310 103.690 ;
      LAYER Nwell ;
        RECT 6.290 95.850 223.310 100.150 ;
      LAYER Pwell ;
        RECT 6.290 92.310 223.310 95.850 ;
      LAYER Nwell ;
        RECT 6.290 88.010 223.310 92.310 ;
      LAYER Pwell ;
        RECT 6.290 84.470 223.310 88.010 ;
      LAYER Nwell ;
        RECT 6.290 80.170 223.310 84.470 ;
      LAYER Pwell ;
        RECT 6.290 76.630 223.310 80.170 ;
      LAYER Nwell ;
        RECT 6.290 72.330 223.310 76.630 ;
      LAYER Pwell ;
        RECT 6.290 68.790 223.310 72.330 ;
      LAYER Nwell ;
        RECT 6.290 64.490 223.310 68.790 ;
      LAYER Pwell ;
        RECT 6.290 60.950 223.310 64.490 ;
      LAYER Nwell ;
        RECT 6.290 56.650 223.310 60.950 ;
      LAYER Pwell ;
        RECT 6.290 53.110 223.310 56.650 ;
      LAYER Nwell ;
        RECT 6.290 48.810 223.310 53.110 ;
      LAYER Pwell ;
        RECT 6.290 45.270 223.310 48.810 ;
      LAYER Nwell ;
        RECT 6.290 40.970 223.310 45.270 ;
      LAYER Pwell ;
        RECT 6.290 37.430 223.310 40.970 ;
      LAYER Nwell ;
        RECT 6.290 33.130 223.310 37.430 ;
      LAYER Pwell ;
        RECT 6.290 29.590 223.310 33.130 ;
      LAYER Nwell ;
        RECT 6.290 25.290 223.310 29.590 ;
      LAYER Pwell ;
        RECT 6.290 21.750 223.310 25.290 ;
      LAYER Nwell ;
        RECT 6.290 17.450 223.310 21.750 ;
      LAYER Pwell ;
        RECT 6.290 15.250 223.310 17.450 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 222.880 211.980 ;
      LAYER Metal2 ;
        RECT 8.540 225.700 8.660 226.000 ;
        RECT 9.820 225.700 27.700 226.000 ;
        RECT 28.860 225.700 46.740 226.000 ;
        RECT 47.900 225.700 65.780 226.000 ;
        RECT 66.940 225.700 84.820 226.000 ;
        RECT 85.980 225.700 103.860 226.000 ;
        RECT 105.020 225.700 122.900 226.000 ;
        RECT 124.060 225.700 141.940 226.000 ;
        RECT 143.100 225.700 160.980 226.000 ;
        RECT 162.140 225.700 180.020 226.000 ;
        RECT 181.180 225.700 199.060 226.000 ;
        RECT 200.220 225.700 218.100 226.000 ;
        RECT 219.260 225.700 219.380 226.000 ;
        RECT 8.540 15.490 219.380 225.700 ;
      LAYER Metal3 ;
        RECT 8.490 15.540 219.430 211.820 ;
      LAYER Metal4 ;
        RECT 74.620 122.730 98.740 171.830 ;
        RECT 100.940 122.730 175.540 171.830 ;
        RECT 177.740 122.730 199.220 171.830 ;
  END
END diceroll
END LIBRARY

