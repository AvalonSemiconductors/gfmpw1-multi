* NGSPICE file created from ue1.ext - technology: gf180mcuD

.subckt ue1 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb io_out[0] io_out[1]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ rst_n vdd vss
.ends

