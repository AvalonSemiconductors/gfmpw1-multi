VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO blinker
  CLASS BLOCK ;
  FOREIGN blinker ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 180.000 ;
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END io_out[2]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 26.710 15.380 28.310 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 68.290 15.380 69.890 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 109.870 15.380 111.470 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 151.450 15.380 153.050 161.020 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 47.500 15.380 49.100 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 89.080 15.380 90.680 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 130.660 15.380 132.260 161.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.240 15.380 173.840 161.020 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 158.560 173.470 161.150 ;
      LAYER Pwell ;
        RECT 6.290 155.040 173.470 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 173.470 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 173.470 150.720 ;
      LAYER Nwell ;
        RECT 6.290 143.005 173.470 147.200 ;
        RECT 6.290 142.880 45.745 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 173.470 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 55.265 139.360 ;
        RECT 6.290 135.165 173.470 139.235 ;
        RECT 6.290 135.040 12.705 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 173.470 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 12.705 131.520 ;
        RECT 6.290 127.325 173.470 131.395 ;
        RECT 6.290 127.200 39.025 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 173.470 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 103.580 123.680 ;
        RECT 6.290 119.485 173.470 123.555 ;
        RECT 6.290 119.360 39.585 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 173.470 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 14.385 115.840 ;
        RECT 6.290 111.645 173.470 115.715 ;
        RECT 6.290 111.520 12.705 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 173.470 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 142.280 108.000 ;
        RECT 6.290 103.805 173.470 107.875 ;
        RECT 6.290 103.680 119.105 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 173.470 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 13.265 100.160 ;
        RECT 6.290 95.965 173.470 100.035 ;
        RECT 6.290 95.840 12.705 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 173.470 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 73.745 92.320 ;
        RECT 6.290 88.125 173.470 92.195 ;
        RECT 6.290 88.000 12.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 173.470 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 19.985 84.480 ;
        RECT 6.290 80.285 173.470 84.355 ;
        RECT 6.290 80.160 14.945 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 173.470 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 32.305 76.640 ;
        RECT 6.290 72.445 173.470 76.515 ;
        RECT 6.290 72.320 12.705 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 173.470 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 148.440 68.800 ;
        RECT 6.290 64.605 173.470 68.675 ;
        RECT 6.290 64.480 43.505 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 173.470 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 91.105 60.960 ;
        RECT 6.290 56.765 173.470 60.835 ;
        RECT 6.290 56.640 71.505 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 173.470 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 65.345 53.120 ;
        RECT 6.290 48.925 173.470 52.995 ;
        RECT 6.290 48.800 160.545 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 173.470 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 64.760 45.280 ;
        RECT 6.290 41.085 173.470 45.155 ;
        RECT 6.290 40.960 61.555 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 173.470 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 97.825 37.440 ;
        RECT 6.290 33.245 173.470 37.315 ;
        RECT 6.290 33.120 80.465 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 173.470 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 118.590 29.600 ;
        RECT 6.290 25.405 173.470 29.475 ;
        RECT 6.290 25.280 129.960 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 173.470 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 12.705 21.760 ;
        RECT 6.290 17.565 173.470 21.635 ;
        RECT 6.290 17.440 51.345 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 173.470 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 173.840 161.020 ;
      LAYER Metal2 ;
        RECT 7.980 4.300 173.700 160.910 ;
        RECT 7.980 4.000 17.620 4.300 ;
        RECT 18.780 4.000 53.460 4.300 ;
        RECT 54.620 4.000 89.300 4.300 ;
        RECT 90.460 4.000 125.140 4.300 ;
        RECT 126.300 4.000 160.980 4.300 ;
        RECT 162.140 4.000 173.700 4.300 ;
      LAYER Metal3 ;
        RECT 7.930 15.540 173.750 160.860 ;
      LAYER Metal4 ;
        RECT 23.100 22.490 26.410 126.470 ;
        RECT 28.610 22.490 47.200 126.470 ;
        RECT 49.400 22.490 67.990 126.470 ;
        RECT 70.190 22.490 88.780 126.470 ;
        RECT 90.980 22.490 109.570 126.470 ;
        RECT 111.770 22.490 130.360 126.470 ;
        RECT 132.560 22.490 134.260 126.470 ;
  END
END blinker
END LIBRARY

