magic
tech gf180mcuD
magscale 1 5
timestamp 1754049408
<< nwell >>
rect 629 1525 121843 120779
<< obsm1 >>
rect 672 407 121800 120945
<< metal2 >>
rect 2016 122100 2072 122500
rect 5712 122100 5768 122500
rect 9408 122100 9464 122500
rect 13104 122100 13160 122500
rect 16800 122100 16856 122500
rect 20496 122100 20552 122500
rect 24192 122100 24248 122500
rect 27888 122100 27944 122500
rect 31584 122100 31640 122500
rect 35280 122100 35336 122500
rect 38976 122100 39032 122500
rect 42672 122100 42728 122500
rect 46368 122100 46424 122500
rect 50064 122100 50120 122500
rect 53760 122100 53816 122500
rect 57456 122100 57512 122500
rect 61152 122100 61208 122500
rect 64848 122100 64904 122500
rect 68544 122100 68600 122500
rect 72240 122100 72296 122500
rect 75936 122100 75992 122500
rect 79632 122100 79688 122500
rect 83328 122100 83384 122500
rect 87024 122100 87080 122500
rect 90720 122100 90776 122500
rect 94416 122100 94472 122500
rect 98112 122100 98168 122500
rect 101808 122100 101864 122500
rect 105504 122100 105560 122500
rect 109200 122100 109256 122500
rect 112896 122100 112952 122500
rect 116592 122100 116648 122500
rect 120288 122100 120344 122500
rect 2016 0 2072 400
rect 5712 0 5768 400
rect 9408 0 9464 400
rect 13104 0 13160 400
rect 16800 0 16856 400
rect 20496 0 20552 400
rect 24192 0 24248 400
rect 27888 0 27944 400
rect 31584 0 31640 400
rect 35280 0 35336 400
rect 38976 0 39032 400
rect 42672 0 42728 400
rect 46368 0 46424 400
rect 50064 0 50120 400
rect 53760 0 53816 400
rect 57456 0 57512 400
rect 61152 0 61208 400
rect 64848 0 64904 400
rect 68544 0 68600 400
rect 72240 0 72296 400
rect 75936 0 75992 400
rect 79632 0 79688 400
rect 83328 0 83384 400
rect 87024 0 87080 400
rect 90720 0 90776 400
rect 94416 0 94472 400
rect 98112 0 98168 400
rect 101808 0 101864 400
rect 105504 0 105560 400
rect 109200 0 109256 400
rect 112896 0 112952 400
rect 116592 0 116648 400
rect 120288 0 120344 400
<< obsm2 >>
rect 574 122070 1986 122100
rect 2102 122070 5682 122100
rect 5798 122070 9378 122100
rect 9494 122070 13074 122100
rect 13190 122070 16770 122100
rect 16886 122070 20466 122100
rect 20582 122070 24162 122100
rect 24278 122070 27858 122100
rect 27974 122070 31554 122100
rect 31670 122070 35250 122100
rect 35366 122070 38946 122100
rect 39062 122070 42642 122100
rect 42758 122070 46338 122100
rect 46454 122070 50034 122100
rect 50150 122070 53730 122100
rect 53846 122070 57426 122100
rect 57542 122070 61122 122100
rect 61238 122070 64818 122100
rect 64934 122070 68514 122100
rect 68630 122070 72210 122100
rect 72326 122070 75906 122100
rect 76022 122070 79602 122100
rect 79718 122070 83298 122100
rect 83414 122070 86994 122100
rect 87110 122070 90690 122100
rect 90806 122070 94386 122100
rect 94502 122070 98082 122100
rect 98198 122070 101778 122100
rect 101894 122070 105474 122100
rect 105590 122070 109170 122100
rect 109286 122070 112866 122100
rect 112982 122070 116562 122100
rect 116678 122070 120258 122100
rect 120374 122070 121730 122100
rect 574 430 121730 122070
rect 574 400 1986 430
rect 2102 400 5682 430
rect 5798 400 9378 430
rect 9494 400 13074 430
rect 13190 400 16770 430
rect 16886 400 20466 430
rect 20582 400 24162 430
rect 24278 400 27858 430
rect 27974 400 31554 430
rect 31670 400 35250 430
rect 35366 400 38946 430
rect 39062 400 42642 430
rect 42758 400 46338 430
rect 46454 400 50034 430
rect 50150 400 53730 430
rect 53846 400 57426 430
rect 57542 400 61122 430
rect 61238 400 64818 430
rect 64934 400 68514 430
rect 68630 400 72210 430
rect 72326 400 75906 430
rect 76022 400 79602 430
rect 79718 400 83298 430
rect 83414 400 86994 430
rect 87110 400 90690 430
rect 90806 400 94386 430
rect 94502 400 98082 430
rect 98198 400 101778 430
rect 101894 400 105474 430
rect 105590 400 109170 430
rect 109286 400 112866 430
rect 112982 400 116562 430
rect 116678 400 120258 430
rect 120374 400 121730 430
<< metal3 >>
rect 0 119616 400 119672
rect 0 116368 400 116424
rect 0 113120 400 113176
rect 0 109872 400 109928
rect 0 106624 400 106680
rect 0 103376 400 103432
rect 0 100128 400 100184
rect 0 96880 400 96936
rect 0 93632 400 93688
rect 0 90384 400 90440
rect 0 87136 400 87192
rect 0 83888 400 83944
rect 0 80640 400 80696
rect 0 77392 400 77448
rect 0 74144 400 74200
rect 0 70896 400 70952
rect 0 67648 400 67704
rect 0 64400 400 64456
rect 0 61152 400 61208
rect 0 57904 400 57960
rect 0 54656 400 54712
rect 0 51408 400 51464
rect 0 48160 400 48216
rect 0 44912 400 44968
rect 0 41664 400 41720
rect 0 38416 400 38472
rect 0 35168 400 35224
rect 0 31920 400 31976
rect 0 28672 400 28728
rect 0 25424 400 25480
rect 0 22176 400 22232
rect 0 18928 400 18984
rect 0 15680 400 15736
rect 0 12432 400 12488
rect 0 9184 400 9240
rect 0 5936 400 5992
rect 0 2688 400 2744
<< obsm3 >>
rect 400 119702 121735 121058
rect 430 119586 121735 119702
rect 400 116454 121735 119586
rect 430 116338 121735 116454
rect 400 113206 121735 116338
rect 430 113090 121735 113206
rect 400 109958 121735 113090
rect 430 109842 121735 109958
rect 400 106710 121735 109842
rect 430 106594 121735 106710
rect 400 103462 121735 106594
rect 430 103346 121735 103462
rect 400 100214 121735 103346
rect 430 100098 121735 100214
rect 400 96966 121735 100098
rect 430 96850 121735 96966
rect 400 93718 121735 96850
rect 430 93602 121735 93718
rect 400 90470 121735 93602
rect 430 90354 121735 90470
rect 400 87222 121735 90354
rect 430 87106 121735 87222
rect 400 83974 121735 87106
rect 430 83858 121735 83974
rect 400 80726 121735 83858
rect 430 80610 121735 80726
rect 400 77478 121735 80610
rect 430 77362 121735 77478
rect 400 74230 121735 77362
rect 430 74114 121735 74230
rect 400 70982 121735 74114
rect 430 70866 121735 70982
rect 400 67734 121735 70866
rect 430 67618 121735 67734
rect 400 64486 121735 67618
rect 430 64370 121735 64486
rect 400 61238 121735 64370
rect 430 61122 121735 61238
rect 400 57990 121735 61122
rect 430 57874 121735 57990
rect 400 54742 121735 57874
rect 430 54626 121735 54742
rect 400 51494 121735 54626
rect 430 51378 121735 51494
rect 400 48246 121735 51378
rect 430 48130 121735 48246
rect 400 44998 121735 48130
rect 430 44882 121735 44998
rect 400 41750 121735 44882
rect 430 41634 121735 41750
rect 400 38502 121735 41634
rect 430 38386 121735 38502
rect 400 35254 121735 38386
rect 430 35138 121735 35254
rect 400 32006 121735 35138
rect 430 31890 121735 32006
rect 400 28758 121735 31890
rect 430 28642 121735 28758
rect 400 25510 121735 28642
rect 430 25394 121735 25510
rect 400 22262 121735 25394
rect 430 22146 121735 22262
rect 400 19014 121735 22146
rect 430 18898 121735 19014
rect 400 15766 121735 18898
rect 430 15650 121735 15766
rect 400 12518 121735 15650
rect 430 12402 121735 12518
rect 400 9270 121735 12402
rect 430 9154 121735 9270
rect 400 6022 121735 9154
rect 430 5906 121735 6022
rect 400 2774 121735 5906
rect 430 2658 121735 2774
rect 400 630 121735 2658
<< metal4 >>
rect 2224 1538 2384 120766
rect 9904 1538 10064 120766
rect 17584 1538 17744 120766
rect 25264 1538 25424 120766
rect 32944 1538 33104 120766
rect 40624 1538 40784 120766
rect 48304 1538 48464 120766
rect 55984 1538 56144 120766
rect 63664 1538 63824 120766
rect 71344 1538 71504 120766
rect 79024 1538 79184 120766
rect 86704 1538 86864 120766
rect 94384 1538 94544 120766
rect 102064 1538 102224 120766
rect 109744 1538 109904 120766
rect 117424 1538 117584 120766
<< obsm4 >>
rect 854 1508 2194 120447
rect 2414 1508 9874 120447
rect 10094 1508 17554 120447
rect 17774 1508 25234 120447
rect 25454 1508 32914 120447
rect 33134 1508 40594 120447
rect 40814 1508 48274 120447
rect 48494 1508 55954 120447
rect 56174 1508 63634 120447
rect 63854 1508 71314 120447
rect 71534 1508 78994 120447
rect 79214 1508 86674 120447
rect 86894 1508 94354 120447
rect 94574 1508 102034 120447
rect 102254 1508 109714 120447
rect 109934 1508 117394 120447
rect 117614 1508 120834 120447
rect 854 737 120834 1508
<< labels >>
rlabel metal3 s 0 9184 400 9240 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 15680 400 15736 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 0 48160 400 48216 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 0 51408 400 51464 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 0 54656 400 54712 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 0 57904 400 57960 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 0 61152 400 61208 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 0 64400 400 64456 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 0 67648 400 67704 6 io_in[16]
port 10 nsew signal input
rlabel metal3 s 0 70896 400 70952 6 io_in[17]
port 11 nsew signal input
rlabel metal3 s 0 74144 400 74200 6 io_in[18]
port 12 nsew signal input
rlabel metal3 s 0 77392 400 77448 6 io_in[19]
port 13 nsew signal input
rlabel metal3 s 0 18928 400 18984 6 io_in[1]
port 14 nsew signal input
rlabel metal3 s 0 80640 400 80696 6 io_in[20]
port 15 nsew signal input
rlabel metal3 s 0 83888 400 83944 6 io_in[21]
port 16 nsew signal input
rlabel metal3 s 0 87136 400 87192 6 io_in[22]
port 17 nsew signal input
rlabel metal3 s 0 90384 400 90440 6 io_in[23]
port 18 nsew signal input
rlabel metal3 s 0 93632 400 93688 6 io_in[24]
port 19 nsew signal input
rlabel metal3 s 0 96880 400 96936 6 io_in[25]
port 20 nsew signal input
rlabel metal3 s 0 100128 400 100184 6 io_in[26]
port 21 nsew signal input
rlabel metal3 s 0 103376 400 103432 6 io_in[27]
port 22 nsew signal input
rlabel metal3 s 0 106624 400 106680 6 io_in[28]
port 23 nsew signal input
rlabel metal3 s 0 109872 400 109928 6 io_in[29]
port 24 nsew signal input
rlabel metal3 s 0 22176 400 22232 6 io_in[2]
port 25 nsew signal input
rlabel metal3 s 0 113120 400 113176 6 io_in[30]
port 26 nsew signal input
rlabel metal3 s 0 116368 400 116424 6 io_in[31]
port 27 nsew signal input
rlabel metal3 s 0 119616 400 119672 6 io_in[32]
port 28 nsew signal input
rlabel metal3 s 0 25424 400 25480 6 io_in[3]
port 29 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 io_in[4]
port 30 nsew signal input
rlabel metal3 s 0 31920 400 31976 6 io_in[5]
port 31 nsew signal input
rlabel metal3 s 0 35168 400 35224 6 io_in[6]
port 32 nsew signal input
rlabel metal3 s 0 38416 400 38472 6 io_in[7]
port 33 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 io_in[8]
port 34 nsew signal input
rlabel metal3 s 0 44912 400 44968 6 io_in[9]
port 35 nsew signal input
rlabel metal2 s 2016 122100 2072 122500 6 io_oeb[0]
port 36 nsew signal output
rlabel metal2 s 38976 122100 39032 122500 6 io_oeb[10]
port 37 nsew signal output
rlabel metal2 s 42672 122100 42728 122500 6 io_oeb[11]
port 38 nsew signal output
rlabel metal2 s 46368 122100 46424 122500 6 io_oeb[12]
port 39 nsew signal output
rlabel metal2 s 50064 122100 50120 122500 6 io_oeb[13]
port 40 nsew signal output
rlabel metal2 s 53760 122100 53816 122500 6 io_oeb[14]
port 41 nsew signal output
rlabel metal2 s 57456 122100 57512 122500 6 io_oeb[15]
port 42 nsew signal output
rlabel metal2 s 61152 122100 61208 122500 6 io_oeb[16]
port 43 nsew signal output
rlabel metal2 s 64848 122100 64904 122500 6 io_oeb[17]
port 44 nsew signal output
rlabel metal2 s 68544 122100 68600 122500 6 io_oeb[18]
port 45 nsew signal output
rlabel metal2 s 72240 122100 72296 122500 6 io_oeb[19]
port 46 nsew signal output
rlabel metal2 s 5712 122100 5768 122500 6 io_oeb[1]
port 47 nsew signal output
rlabel metal2 s 75936 122100 75992 122500 6 io_oeb[20]
port 48 nsew signal output
rlabel metal2 s 79632 122100 79688 122500 6 io_oeb[21]
port 49 nsew signal output
rlabel metal2 s 83328 122100 83384 122500 6 io_oeb[22]
port 50 nsew signal output
rlabel metal2 s 87024 122100 87080 122500 6 io_oeb[23]
port 51 nsew signal output
rlabel metal2 s 90720 122100 90776 122500 6 io_oeb[24]
port 52 nsew signal output
rlabel metal2 s 94416 122100 94472 122500 6 io_oeb[25]
port 53 nsew signal output
rlabel metal2 s 98112 122100 98168 122500 6 io_oeb[26]
port 54 nsew signal output
rlabel metal2 s 101808 122100 101864 122500 6 io_oeb[27]
port 55 nsew signal output
rlabel metal2 s 105504 122100 105560 122500 6 io_oeb[28]
port 56 nsew signal output
rlabel metal2 s 109200 122100 109256 122500 6 io_oeb[29]
port 57 nsew signal output
rlabel metal2 s 9408 122100 9464 122500 6 io_oeb[2]
port 58 nsew signal output
rlabel metal2 s 112896 122100 112952 122500 6 io_oeb[30]
port 59 nsew signal output
rlabel metal2 s 116592 122100 116648 122500 6 io_oeb[31]
port 60 nsew signal output
rlabel metal2 s 120288 122100 120344 122500 6 io_oeb[32]
port 61 nsew signal output
rlabel metal2 s 13104 122100 13160 122500 6 io_oeb[3]
port 62 nsew signal output
rlabel metal2 s 16800 122100 16856 122500 6 io_oeb[4]
port 63 nsew signal output
rlabel metal2 s 20496 122100 20552 122500 6 io_oeb[5]
port 64 nsew signal output
rlabel metal2 s 24192 122100 24248 122500 6 io_oeb[6]
port 65 nsew signal output
rlabel metal2 s 27888 122100 27944 122500 6 io_oeb[7]
port 66 nsew signal output
rlabel metal2 s 31584 122100 31640 122500 6 io_oeb[8]
port 67 nsew signal output
rlabel metal2 s 35280 122100 35336 122500 6 io_oeb[9]
port 68 nsew signal output
rlabel metal2 s 2016 0 2072 400 6 io_out[0]
port 69 nsew signal output
rlabel metal2 s 38976 0 39032 400 6 io_out[10]
port 70 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 io_out[11]
port 71 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 io_out[12]
port 72 nsew signal output
rlabel metal2 s 50064 0 50120 400 6 io_out[13]
port 73 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 io_out[14]
port 74 nsew signal output
rlabel metal2 s 57456 0 57512 400 6 io_out[15]
port 75 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 io_out[16]
port 76 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 io_out[17]
port 77 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 io_out[18]
port 78 nsew signal output
rlabel metal2 s 72240 0 72296 400 6 io_out[19]
port 79 nsew signal output
rlabel metal2 s 5712 0 5768 400 6 io_out[1]
port 80 nsew signal output
rlabel metal2 s 75936 0 75992 400 6 io_out[20]
port 81 nsew signal output
rlabel metal2 s 79632 0 79688 400 6 io_out[21]
port 82 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 io_out[22]
port 83 nsew signal output
rlabel metal2 s 87024 0 87080 400 6 io_out[23]
port 84 nsew signal output
rlabel metal2 s 90720 0 90776 400 6 io_out[24]
port 85 nsew signal output
rlabel metal2 s 94416 0 94472 400 6 io_out[25]
port 86 nsew signal output
rlabel metal2 s 98112 0 98168 400 6 io_out[26]
port 87 nsew signal output
rlabel metal2 s 101808 0 101864 400 6 io_out[27]
port 88 nsew signal output
rlabel metal2 s 105504 0 105560 400 6 io_out[28]
port 89 nsew signal output
rlabel metal2 s 109200 0 109256 400 6 io_out[29]
port 90 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 io_out[2]
port 91 nsew signal output
rlabel metal2 s 112896 0 112952 400 6 io_out[30]
port 92 nsew signal output
rlabel metal2 s 116592 0 116648 400 6 io_out[31]
port 93 nsew signal output
rlabel metal2 s 120288 0 120344 400 6 io_out[32]
port 94 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 io_out[3]
port 95 nsew signal output
rlabel metal2 s 16800 0 16856 400 6 io_out[4]
port 96 nsew signal output
rlabel metal2 s 20496 0 20552 400 6 io_out[5]
port 97 nsew signal output
rlabel metal2 s 24192 0 24248 400 6 io_out[6]
port 98 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 io_out[7]
port 99 nsew signal output
rlabel metal2 s 31584 0 31640 400 6 io_out[8]
port 100 nsew signal output
rlabel metal2 s 35280 0 35336 400 6 io_out[9]
port 101 nsew signal output
rlabel metal3 s 0 5936 400 5992 6 rst_n
port 102 nsew signal input
rlabel metal4 s 2224 1538 2384 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 120766 6 vdd
port 103 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 120766 6 vss
port 104 nsew ground bidirectional
rlabel metal3 s 0 2688 400 2744 6 wb_clk_i
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 122500 122500
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 50409476
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_tholin_riscv/runs/25_08_01_12_59/results/signoff/wrapped_tholin_riscv.magic.gds
string GDS_START 307870
<< end >>

