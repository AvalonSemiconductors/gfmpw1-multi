magic
tech gf180mcuD
magscale 1 5
timestamp 1753967824
<< nwell >>
rect 629 20561 22331 20991
rect 629 19777 22331 20207
rect 629 18993 22331 19423
rect 629 18209 22331 18639
rect 629 17425 22331 17855
rect 629 16641 22331 17071
rect 629 15857 22331 16287
rect 629 15073 22331 15503
rect 629 14289 22331 14719
rect 629 13505 22331 13935
rect 629 12721 22331 13151
rect 629 11937 22331 12367
rect 629 11153 22331 11583
rect 629 10369 22331 10799
rect 629 9585 22331 10015
rect 629 8801 22331 9231
rect 629 8017 22331 8447
rect 629 7233 22331 7663
rect 629 6449 22331 6879
rect 629 5665 22331 6095
rect 629 4881 22331 5311
rect 629 4097 22331 4527
rect 629 3313 22331 3743
rect 629 2529 22331 2959
rect 629 1745 22331 2175
<< pwell >>
rect 629 20991 22331 21211
rect 629 20207 22331 20561
rect 629 19423 22331 19777
rect 629 18639 22331 18993
rect 629 17855 22331 18209
rect 629 17071 22331 17425
rect 629 16287 22331 16641
rect 629 15503 22331 15857
rect 629 14719 22331 15073
rect 629 13935 22331 14289
rect 629 13151 22331 13505
rect 629 12367 22331 12721
rect 629 11583 22331 11937
rect 629 10799 22331 11153
rect 629 10015 22331 10369
rect 629 9231 22331 9585
rect 629 8447 22331 8801
rect 629 7663 22331 8017
rect 629 6879 22331 7233
rect 629 6095 22331 6449
rect 629 5311 22331 5665
rect 629 4527 22331 4881
rect 629 3743 22331 4097
rect 629 2959 22331 3313
rect 629 2175 22331 2529
rect 629 1525 22331 1745
<< obsm1 >>
rect 672 1538 22288 21198
<< obsm2 >>
rect 2238 1353 22274 21551
<< metal3 >>
rect 22600 21504 23000 21560
rect 22600 19824 23000 19880
rect 22600 18144 23000 18200
rect 22600 16464 23000 16520
rect 22600 14784 23000 14840
rect 22600 13104 23000 13160
rect 22600 11424 23000 11480
rect 22600 9744 23000 9800
rect 22600 8064 23000 8120
rect 22600 6384 23000 6440
rect 22600 4704 23000 4760
rect 22600 3024 23000 3080
rect 22600 1344 23000 1400
<< obsm3 >>
rect 2233 21474 22570 21546
rect 2233 19910 22600 21474
rect 2233 19794 22570 19910
rect 2233 18230 22600 19794
rect 2233 18114 22570 18230
rect 2233 16550 22600 18114
rect 2233 16434 22570 16550
rect 2233 14870 22600 16434
rect 2233 14754 22570 14870
rect 2233 13190 22600 14754
rect 2233 13074 22570 13190
rect 2233 11510 22600 13074
rect 2233 11394 22570 11510
rect 2233 9830 22600 11394
rect 2233 9714 22570 9830
rect 2233 8150 22600 9714
rect 2233 8034 22570 8150
rect 2233 6470 22600 8034
rect 2233 6354 22570 6470
rect 2233 4790 22600 6354
rect 2233 4674 22570 4790
rect 2233 3110 22600 4674
rect 2233 2994 22570 3110
rect 2233 1430 22600 2994
rect 2233 1358 22570 1430
<< metal4 >>
rect 2224 1538 2384 21198
rect 9904 1538 10064 21198
rect 17584 1538 17744 21198
<< obsm4 >>
rect 8414 2137 9874 18807
rect 10094 2137 17554 18807
rect 17774 2137 21994 18807
<< labels >>
rlabel metal3 s 22600 1344 23000 1400 6 clk
port 1 nsew signal input
rlabel metal3 s 22600 4704 23000 4760 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 22600 6384 23000 6440 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 22600 8064 23000 8120 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 22600 9744 23000 9800 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 22600 11424 23000 11480 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 22600 13104 23000 13160 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 22600 14784 23000 14840 6 io_out[0]
port 8 nsew signal output
rlabel metal3 s 22600 16464 23000 16520 6 io_out[1]
port 9 nsew signal output
rlabel metal3 s 22600 18144 23000 18200 6 io_out[2]
port 10 nsew signal output
rlabel metal3 s 22600 19824 23000 19880 6 io_out[3]
port 11 nsew signal output
rlabel metal3 s 22600 21504 23000 21560 6 io_out[4]
port 12 nsew signal output
rlabel metal3 s 22600 3024 23000 3080 6 rst_n
port 13 nsew signal input
rlabel metal4 s 2224 1538 2384 21198 6 vdd
port 14 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 21198 6 vdd
port 14 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 21198 6 vss
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1291474
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/tbb1143/runs/25_07_31_15_15/results/signoff/tholin_avalonsemi_tbb1143.magic.gds
string GDS_START 193762
<< end >>

