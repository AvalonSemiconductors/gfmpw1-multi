magic
tech gf180mcuD
magscale 1 10
timestamp 1699956754
<< nwell >>
rect 1258 55257 58662 56096
rect 1258 55232 18333 55257
rect 1258 54503 18221 54528
rect 1258 53689 58662 54503
rect 1258 53664 33160 53689
rect 1258 52121 58662 52960
rect 1258 52096 15981 52121
rect 1258 51367 35021 51392
rect 1258 50553 58662 51367
rect 1258 50528 23485 50553
rect 1258 49799 13224 49824
rect 1258 48985 58662 49799
rect 1258 48960 16205 48985
rect 1258 48231 6909 48256
rect 1258 47417 58662 48231
rect 1258 47392 26539 47417
rect 1258 46663 6056 46688
rect 1258 45849 58662 46663
rect 1258 45824 48013 45849
rect 1258 45095 16101 45120
rect 1258 44281 58662 45095
rect 1258 44256 18221 44281
rect 1258 43527 6616 43552
rect 1258 42713 58662 43527
rect 1258 42688 25165 42713
rect 1258 41959 12733 41984
rect 1258 41145 58662 41959
rect 1258 41120 9261 41145
rect 1258 40391 12173 40416
rect 1258 39577 58662 40391
rect 1258 39552 2541 39577
rect 1258 38823 2541 38848
rect 1258 38009 58662 38823
rect 1258 37984 17101 38009
rect 1258 37255 13293 37280
rect 1258 36441 58662 37255
rect 1258 36416 2541 36441
rect 1258 35687 20685 35712
rect 1258 34873 58662 35687
rect 1258 34848 10312 34873
rect 1258 34119 12509 34144
rect 1258 33305 58662 34119
rect 1258 33280 2541 33305
rect 1258 32551 2541 32576
rect 1258 31737 58662 32551
rect 1258 31712 11880 31737
rect 1258 30983 13853 31008
rect 1258 30169 58662 30983
rect 1258 30144 2541 30169
rect 1258 29415 22141 29440
rect 1258 28601 58662 29415
rect 1258 28576 18445 28601
rect 1258 27847 2541 27872
rect 1258 27008 58662 27847
rect 1258 26279 12776 26304
rect 1258 25465 58662 26279
rect 1258 25440 8813 25465
rect 1258 24711 2541 24736
rect 1258 23897 58662 24711
rect 1258 23872 18669 23897
rect 1258 23143 2541 23168
rect 1258 22329 58662 23143
rect 1258 22304 7469 22329
rect 1258 21575 33901 21600
rect 1258 20761 58662 21575
rect 1258 20736 2541 20761
rect 1258 20007 10381 20032
rect 1258 19193 58662 20007
rect 1258 19168 16808 19193
rect 1258 18439 6392 18464
rect 1258 17625 58662 18439
rect 1258 17600 2541 17625
rect 1258 16871 21288 16896
rect 1258 16057 58662 16871
rect 1258 16032 10760 16057
rect 1258 15303 5565 15328
rect 1258 14489 58662 15303
rect 1258 14464 2541 14489
rect 1258 13735 11165 13760
rect 1258 12921 58662 13735
rect 1258 12896 7133 12921
rect 1258 12167 20013 12192
rect 1258 11353 58662 12167
rect 1258 11328 2541 11353
rect 1258 10599 19677 10624
rect 1258 9785 58662 10599
rect 1258 9760 2989 9785
rect 1258 9031 18221 9056
rect 1258 8217 58662 9031
rect 1258 8192 19160 8217
rect 1258 7463 12061 7488
rect 1258 6649 58662 7463
rect 1258 6624 7848 6649
rect 1258 5895 38269 5920
rect 1258 5081 58662 5895
rect 1258 5056 10717 5081
rect 1258 4327 10941 4352
rect 1258 3513 58662 4327
rect 1258 3488 44429 3513
<< pwell >>
rect 1258 56096 58662 56534
rect 1258 54528 58662 55232
rect 1258 52960 58662 53664
rect 1258 51392 58662 52096
rect 1258 49824 58662 50528
rect 1258 48256 58662 48960
rect 1258 46688 58662 47392
rect 1258 45120 58662 45824
rect 1258 43552 58662 44256
rect 1258 41984 58662 42688
rect 1258 40416 58662 41120
rect 1258 38848 58662 39552
rect 1258 37280 58662 37984
rect 1258 35712 58662 36416
rect 1258 34144 58662 34848
rect 1258 32576 58662 33280
rect 1258 31008 58662 31712
rect 1258 29440 58662 30144
rect 1258 27872 58662 28576
rect 1258 26304 58662 27008
rect 1258 24736 58662 25440
rect 1258 23168 58662 23872
rect 1258 21600 58662 22304
rect 1258 20032 58662 20736
rect 1258 18464 58662 19168
rect 1258 16896 58662 17600
rect 1258 15328 58662 16032
rect 1258 13760 58662 14464
rect 1258 12192 58662 12896
rect 1258 10624 58662 11328
rect 1258 9056 58662 9760
rect 1258 7488 58662 8192
rect 1258 5920 58662 6624
rect 1258 4352 58662 5056
rect 1258 3050 58662 3488
<< obsm1 >>
rect 1344 1710 58576 56508
<< metal2 >>
rect 7392 59200 7504 60000
rect 22400 59200 22512 60000
rect 37408 59200 37520 60000
rect 52416 59200 52528 60000
rect 2688 0 2800 800
rect 4704 0 4816 800
rect 6720 0 6832 800
rect 8736 0 8848 800
rect 10752 0 10864 800
rect 12768 0 12880 800
rect 14784 0 14896 800
rect 16800 0 16912 800
rect 18816 0 18928 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 24864 0 24976 800
rect 26880 0 26992 800
rect 28896 0 29008 800
rect 30912 0 31024 800
rect 32928 0 33040 800
rect 34944 0 35056 800
rect 36960 0 37072 800
rect 38976 0 39088 800
rect 40992 0 41104 800
rect 43008 0 43120 800
rect 45024 0 45136 800
rect 47040 0 47152 800
rect 49056 0 49168 800
rect 51072 0 51184 800
rect 53088 0 53200 800
rect 55104 0 55216 800
rect 57120 0 57232 800
<< obsm2 >>
rect 1820 59140 7332 59200
rect 7564 59140 22340 59200
rect 22572 59140 37348 59200
rect 37580 59140 52356 59200
rect 52588 59140 58324 59200
rect 1820 860 58324 59140
rect 1820 700 2628 860
rect 2860 700 4644 860
rect 4876 700 6660 860
rect 6892 700 8676 860
rect 8908 700 10692 860
rect 10924 700 12708 860
rect 12940 700 14724 860
rect 14956 700 16740 860
rect 16972 700 18756 860
rect 18988 700 20772 860
rect 21004 700 22788 860
rect 23020 700 24804 860
rect 25036 700 26820 860
rect 27052 700 28836 860
rect 29068 700 30852 860
rect 31084 700 32868 860
rect 33100 700 34884 860
rect 35116 700 36900 860
rect 37132 700 38916 860
rect 39148 700 40932 860
rect 41164 700 42948 860
rect 43180 700 44964 860
rect 45196 700 46980 860
rect 47212 700 48996 860
rect 49228 700 51012 860
rect 51244 700 53028 860
rect 53260 700 55044 860
rect 55276 700 57060 860
rect 57292 700 58324 860
<< metal3 >>
rect 59200 56000 60000 56112
rect 59200 50176 60000 50288
rect 59200 44352 60000 44464
rect 59200 38528 60000 38640
rect 59200 32704 60000 32816
rect 59200 26880 60000 26992
rect 59200 21056 60000 21168
rect 59200 15232 60000 15344
rect 59200 9408 60000 9520
rect 59200 3584 60000 3696
<< obsm3 >>
rect 1810 56172 59200 56476
rect 1810 55940 59140 56172
rect 1810 50348 59200 55940
rect 1810 50116 59140 50348
rect 1810 44524 59200 50116
rect 1810 44292 59140 44524
rect 1810 38700 59200 44292
rect 1810 38468 59140 38700
rect 1810 32876 59200 38468
rect 1810 32644 59140 32876
rect 1810 27052 59200 32644
rect 1810 26820 59140 27052
rect 1810 21228 59200 26820
rect 1810 20996 59140 21228
rect 1810 15404 59200 20996
rect 1810 15172 59140 15404
rect 1810 9580 59200 15172
rect 1810 9348 59140 9580
rect 1810 3756 59200 9348
rect 1810 3524 59140 3756
rect 1810 3108 59200 3524
<< metal4 >>
rect 4448 3076 4768 56508
rect 19808 3076 20128 56508
rect 35168 3076 35488 56508
rect 50528 3076 50848 56508
<< obsm4 >>
rect 8652 7186 19748 55982
rect 20188 7186 35108 55982
rect 35548 7186 50468 55982
rect 50908 7186 54516 55982
<< labels >>
rlabel metal3 s 59200 50176 60000 50288 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 59200 56000 60000 56112 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 59200 3584 60000 3696 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 59200 9408 60000 9520 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 59200 15232 60000 15344 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 59200 21056 60000 21168 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 59200 26880 60000 26992 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 59200 32704 60000 32816 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 59200 38528 60000 38640 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 59200 44352 60000 44464 6 io_in_1[7]
port 10 nsew signal input
rlabel metal2 s 37408 59200 37520 60000 6 io_in_2[0]
port 11 nsew signal input
rlabel metal2 s 52416 59200 52528 60000 6 io_in_2[1]
port 12 nsew signal input
rlabel metal2 s 2688 0 2800 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 22848 0 22960 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 24864 0 24976 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 26880 0 26992 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 28896 0 29008 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 30912 0 31024 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 32928 0 33040 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 34944 0 35056 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 36960 0 37072 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 38976 0 39088 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 40992 0 41104 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 4704 0 4816 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 43008 0 43120 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 45024 0 45136 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 47040 0 47152 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 49056 0 49168 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 51072 0 51184 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 53088 0 53200 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 55104 0 55216 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 57120 0 57232 800 6 io_out[27]
port 32 nsew signal output
rlabel metal2 s 6720 0 6832 800 6 io_out[2]
port 33 nsew signal output
rlabel metal2 s 8736 0 8848 800 6 io_out[3]
port 34 nsew signal output
rlabel metal2 s 10752 0 10864 800 6 io_out[4]
port 35 nsew signal output
rlabel metal2 s 12768 0 12880 800 6 io_out[5]
port 36 nsew signal output
rlabel metal2 s 14784 0 14896 800 6 io_out[6]
port 37 nsew signal output
rlabel metal2 s 16800 0 16912 800 6 io_out[7]
port 38 nsew signal output
rlabel metal2 s 18816 0 18928 800 6 io_out[8]
port 39 nsew signal output
rlabel metal2 s 20832 0 20944 800 6 io_out[9]
port 40 nsew signal output
rlabel metal2 s 22400 59200 22512 60000 6 rst_n
port 41 nsew signal input
rlabel metal4 s 4448 3076 4768 56508 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 56508 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 56508 6 vss
port 43 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 56508 6 vss
port 43 nsew ground bidirectional
rlabel metal2 s 7392 59200 7504 60000 6 wb_clk_i
port 44 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2340848
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_ay8913/runs/23_11_14_11_09/results/signoff/wrapped_ay8913.magic.gds
string GDS_START 289154
<< end >>

