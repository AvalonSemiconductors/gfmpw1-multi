magic
tech gf180mcuD
magscale 1 10
timestamp 1698916418
<< metal1 >>
rect 8754 66782 8766 66834
rect 8818 66831 8830 66834
rect 9314 66831 9326 66834
rect 8818 66785 9326 66831
rect 8818 66782 8830 66785
rect 9314 66782 9326 66785
rect 9378 66782 9390 66834
rect 1344 66666 58576 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 58576 66666
rect 1344 66580 58576 66614
rect 26126 66498 26178 66510
rect 26126 66434 26178 66446
rect 40798 66498 40850 66510
rect 40798 66434 40850 66446
rect 43822 66498 43874 66510
rect 43822 66434 43874 66446
rect 48414 66498 48466 66510
rect 48414 66434 48466 66446
rect 52222 66498 52274 66510
rect 52222 66434 52274 66446
rect 56030 66498 56082 66510
rect 56030 66434 56082 66446
rect 18834 66334 18846 66386
rect 18898 66334 18910 66386
rect 22866 66334 22878 66386
rect 22930 66334 22942 66386
rect 36978 66334 36990 66386
rect 37042 66334 37054 66386
rect 17602 66222 17614 66274
rect 17666 66222 17678 66274
rect 23538 66222 23550 66274
rect 23602 66222 23614 66274
rect 25106 66222 25118 66274
rect 25170 66222 25182 66274
rect 39218 66222 39230 66274
rect 39282 66222 39294 66274
rect 39778 66222 39790 66274
rect 39842 66222 39854 66274
rect 46162 66222 46174 66274
rect 46226 66222 46238 66274
rect 47394 66222 47406 66274
rect 47458 66222 47470 66274
rect 51202 66222 51214 66274
rect 51266 66222 51278 66274
rect 55010 66222 55022 66274
rect 55074 66222 55086 66274
rect 2942 66162 2994 66174
rect 2942 66098 2994 66110
rect 5518 66162 5570 66174
rect 5518 66098 5570 66110
rect 6974 66162 7026 66174
rect 6974 66098 7026 66110
rect 9326 66162 9378 66174
rect 9326 66098 9378 66110
rect 11006 66162 11058 66174
rect 11006 66098 11058 66110
rect 13134 66162 13186 66174
rect 13134 66098 13186 66110
rect 15038 66162 15090 66174
rect 15038 66098 15090 66110
rect 17054 66162 17106 66174
rect 17054 66098 17106 66110
rect 29150 66162 29202 66174
rect 29150 66098 29202 66110
rect 31166 66162 31218 66174
rect 31166 66098 31218 66110
rect 33182 66162 33234 66174
rect 33182 66098 33234 66110
rect 35198 66162 35250 66174
rect 35198 66098 35250 66110
rect 43038 66162 43090 66174
rect 43038 66098 43090 66110
rect 1344 65882 58576 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 58576 65882
rect 1344 65796 58576 65830
rect 34862 65602 34914 65614
rect 34862 65538 34914 65550
rect 57822 65602 57874 65614
rect 57822 65538 57874 65550
rect 35534 65490 35586 65502
rect 57598 65490 57650 65502
rect 20178 65438 20190 65490
rect 20242 65438 20254 65490
rect 21858 65438 21870 65490
rect 21922 65438 21934 65490
rect 29698 65438 29710 65490
rect 29762 65438 29774 65490
rect 36642 65438 36654 65490
rect 36706 65438 36718 65490
rect 44370 65438 44382 65490
rect 44434 65438 44446 65490
rect 44818 65438 44830 65490
rect 44882 65438 44894 65490
rect 48850 65438 48862 65490
rect 48914 65438 48926 65490
rect 54898 65438 54910 65490
rect 54962 65438 54974 65490
rect 35534 65426 35586 65438
rect 57598 65426 57650 65438
rect 58158 65490 58210 65502
rect 58158 65426 58210 65438
rect 12574 65378 12626 65390
rect 12574 65314 12626 65326
rect 13246 65378 13298 65390
rect 20862 65378 20914 65390
rect 25454 65378 25506 65390
rect 17378 65326 17390 65378
rect 17442 65326 17454 65378
rect 19506 65326 19518 65378
rect 19570 65326 19582 65378
rect 22530 65326 22542 65378
rect 22594 65326 22606 65378
rect 24658 65326 24670 65378
rect 24722 65326 24734 65378
rect 13246 65314 13298 65326
rect 20862 65314 20914 65326
rect 25454 65314 25506 65326
rect 27358 65378 27410 65390
rect 27358 65314 27410 65326
rect 30270 65378 30322 65390
rect 30270 65314 30322 65326
rect 34974 65378 35026 65390
rect 40126 65378 40178 65390
rect 37426 65326 37438 65378
rect 37490 65326 37502 65378
rect 39554 65326 39566 65378
rect 39618 65326 39630 65378
rect 34974 65314 35026 65326
rect 40126 65314 40178 65326
rect 41134 65378 41186 65390
rect 55470 65378 55522 65390
rect 41570 65326 41582 65378
rect 41634 65326 41646 65378
rect 43698 65326 43710 65378
rect 43762 65326 43774 65378
rect 45602 65326 45614 65378
rect 45666 65326 45678 65378
rect 47730 65326 47742 65378
rect 47794 65326 47806 65378
rect 49522 65326 49534 65378
rect 49586 65326 49598 65378
rect 51650 65326 51662 65378
rect 51714 65326 51726 65378
rect 51986 65326 51998 65378
rect 52050 65326 52062 65378
rect 54114 65326 54126 65378
rect 54178 65326 54190 65378
rect 41134 65314 41186 65326
rect 55470 65314 55522 65326
rect 35086 65266 35138 65278
rect 35086 65202 35138 65214
rect 1344 65098 58576 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 58576 65098
rect 1344 65012 58576 65046
rect 23550 64930 23602 64942
rect 23550 64866 23602 64878
rect 42702 64930 42754 64942
rect 42702 64866 42754 64878
rect 47518 64930 47570 64942
rect 47518 64866 47570 64878
rect 50206 64930 50258 64942
rect 50206 64866 50258 64878
rect 51774 64930 51826 64942
rect 51774 64866 51826 64878
rect 44942 64818 44994 64830
rect 8530 64766 8542 64818
rect 8594 64766 8606 64818
rect 10098 64766 10110 64818
rect 10162 64766 10174 64818
rect 12226 64766 12238 64818
rect 12290 64766 12302 64818
rect 12786 64766 12798 64818
rect 12850 64766 12862 64818
rect 16370 64766 16382 64818
rect 16434 64766 16446 64818
rect 20738 64766 20750 64818
rect 20802 64766 20814 64818
rect 26898 64766 26910 64818
rect 26962 64766 26974 64818
rect 33506 64766 33518 64818
rect 33570 64766 33582 64818
rect 35634 64766 35646 64818
rect 35698 64766 35710 64818
rect 41346 64766 41358 64818
rect 41410 64766 41422 64818
rect 44942 64754 44994 64766
rect 45390 64818 45442 64830
rect 45390 64754 45442 64766
rect 54910 64818 54962 64830
rect 55234 64766 55246 64818
rect 55298 64766 55310 64818
rect 54910 64754 54962 64766
rect 8878 64706 8930 64718
rect 16830 64706 16882 64718
rect 27918 64706 27970 64718
rect 5730 64654 5742 64706
rect 5794 64654 5806 64706
rect 9426 64654 9438 64706
rect 9490 64654 9502 64706
rect 13570 64654 13582 64706
rect 13634 64654 13646 64706
rect 17938 64654 17950 64706
rect 18002 64654 18014 64706
rect 23986 64654 23998 64706
rect 24050 64654 24062 64706
rect 8878 64642 8930 64654
rect 16830 64642 16882 64654
rect 27918 64642 27970 64654
rect 29038 64706 29090 64718
rect 29038 64642 29090 64654
rect 29486 64706 29538 64718
rect 29486 64642 29538 64654
rect 30382 64706 30434 64718
rect 37102 64706 37154 64718
rect 36418 64654 36430 64706
rect 36482 64654 36494 64706
rect 38546 64654 38558 64706
rect 38610 64654 38622 64706
rect 41682 64654 41694 64706
rect 41746 64654 41758 64706
rect 49410 64654 49422 64706
rect 49474 64654 49486 64706
rect 58146 64654 58158 64706
rect 58210 64654 58222 64706
rect 30382 64642 30434 64654
rect 37102 64642 37154 64654
rect 12574 64594 12626 64606
rect 23662 64594 23714 64606
rect 30942 64594 30994 64606
rect 6402 64542 6414 64594
rect 6466 64542 6478 64594
rect 14242 64542 14254 64594
rect 14306 64542 14318 64594
rect 18610 64542 18622 64594
rect 18674 64542 18686 64594
rect 24770 64542 24782 64594
rect 24834 64542 24846 64594
rect 12574 64530 12626 64542
rect 23662 64530 23714 64542
rect 30942 64530 30994 64542
rect 32510 64594 32562 64606
rect 32510 64530 32562 64542
rect 32622 64594 32674 64606
rect 32622 64530 32674 64542
rect 32958 64594 33010 64606
rect 50318 64594 50370 64606
rect 39218 64542 39230 64594
rect 39282 64542 39294 64594
rect 32958 64530 33010 64542
rect 50318 64530 50370 64542
rect 51662 64594 51714 64606
rect 57362 64542 57374 64594
rect 57426 64542 57438 64594
rect 51662 64530 51714 64542
rect 8990 64482 9042 64494
rect 8990 64418 9042 64430
rect 12798 64482 12850 64494
rect 12798 64418 12850 64430
rect 21422 64482 21474 64494
rect 21422 64418 21474 64430
rect 23214 64482 23266 64494
rect 23214 64418 23266 64430
rect 27246 64482 27298 64494
rect 27246 64418 27298 64430
rect 27358 64482 27410 64494
rect 27358 64418 27410 64430
rect 27470 64482 27522 64494
rect 27470 64418 27522 64430
rect 28702 64482 28754 64494
rect 28702 64418 28754 64430
rect 29598 64482 29650 64494
rect 29598 64418 29650 64430
rect 29710 64482 29762 64494
rect 29710 64418 29762 64430
rect 30830 64482 30882 64494
rect 30830 64418 30882 64430
rect 31054 64482 31106 64494
rect 31054 64418 31106 64430
rect 31502 64482 31554 64494
rect 31502 64418 31554 64430
rect 32286 64482 32338 64494
rect 32286 64418 32338 64430
rect 33070 64482 33122 64494
rect 33070 64418 33122 64430
rect 33294 64482 33346 64494
rect 33294 64418 33346 64430
rect 52782 64482 52834 64494
rect 52782 64418 52834 64430
rect 1344 64314 58576 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 58576 64314
rect 1344 64228 58576 64262
rect 8766 64146 8818 64158
rect 17614 64146 17666 64158
rect 11330 64094 11342 64146
rect 11394 64094 11406 64146
rect 8766 64082 8818 64094
rect 17614 64082 17666 64094
rect 27806 64146 27858 64158
rect 27806 64082 27858 64094
rect 32286 64146 32338 64158
rect 32286 64082 32338 64094
rect 41582 64146 41634 64158
rect 41582 64082 41634 64094
rect 42030 64146 42082 64158
rect 50430 64146 50482 64158
rect 46946 64094 46958 64146
rect 47010 64094 47022 64146
rect 42030 64082 42082 64094
rect 50430 64082 50482 64094
rect 52334 64146 52386 64158
rect 52334 64082 52386 64094
rect 54574 64146 54626 64158
rect 54574 64082 54626 64094
rect 13694 64034 13746 64046
rect 12898 63982 12910 64034
rect 12962 63982 12974 64034
rect 13694 63970 13746 63982
rect 13806 64034 13858 64046
rect 13806 63970 13858 63982
rect 14142 64034 14194 64046
rect 14142 63970 14194 63982
rect 27470 64034 27522 64046
rect 27470 63970 27522 63982
rect 27582 64034 27634 64046
rect 55246 64034 55298 64046
rect 31938 63982 31950 64034
rect 32002 63982 32014 64034
rect 35186 63982 35198 64034
rect 35250 63982 35262 64034
rect 46050 63982 46062 64034
rect 46114 63982 46126 64034
rect 50866 63982 50878 64034
rect 50930 64031 50942 64034
rect 51202 64031 51214 64034
rect 50930 63985 51214 64031
rect 50930 63982 50942 63985
rect 51202 63982 51214 63985
rect 51266 63982 51278 64034
rect 27582 63970 27634 63982
rect 55246 63970 55298 63982
rect 55806 64034 55858 64046
rect 55806 63970 55858 63982
rect 14254 63922 14306 63934
rect 11666 63870 11678 63922
rect 11730 63870 11742 63922
rect 12562 63870 12574 63922
rect 12626 63870 12638 63922
rect 14254 63858 14306 63870
rect 17278 63922 17330 63934
rect 17278 63858 17330 63870
rect 17614 63922 17666 63934
rect 17614 63858 17666 63870
rect 17838 63922 17890 63934
rect 23438 63922 23490 63934
rect 32510 63922 32562 63934
rect 39454 63922 39506 63934
rect 43822 63922 43874 63934
rect 49534 63922 49586 63934
rect 20178 63870 20190 63922
rect 20242 63870 20254 63922
rect 26674 63870 26686 63922
rect 26738 63870 26750 63922
rect 28018 63870 28030 63922
rect 28082 63870 28094 63922
rect 32050 63870 32062 63922
rect 32114 63870 32126 63922
rect 33506 63870 33518 63922
rect 33570 63870 33582 63922
rect 34626 63870 34638 63922
rect 34690 63870 34702 63922
rect 43362 63870 43374 63922
rect 43426 63870 43438 63922
rect 45938 63870 45950 63922
rect 46002 63870 46014 63922
rect 46946 63870 46958 63922
rect 47010 63870 47022 63922
rect 17838 63858 17890 63870
rect 23438 63858 23490 63870
rect 32510 63858 32562 63870
rect 39454 63858 39506 63870
rect 43822 63858 43874 63870
rect 49534 63858 49586 63870
rect 49646 63922 49698 63934
rect 49646 63858 49698 63870
rect 49982 63922 50034 63934
rect 49982 63858 50034 63870
rect 50094 63922 50146 63934
rect 54126 63922 54178 63934
rect 51314 63870 51326 63922
rect 51378 63870 51390 63922
rect 50094 63858 50146 63870
rect 54126 63858 54178 63870
rect 54798 63922 54850 63934
rect 54798 63858 54850 63870
rect 27134 63810 27186 63822
rect 32398 63810 32450 63822
rect 50430 63810 50482 63822
rect 20850 63758 20862 63810
rect 20914 63758 20926 63810
rect 22978 63758 22990 63810
rect 23042 63758 23054 63810
rect 26338 63758 26350 63810
rect 26402 63758 26414 63810
rect 28802 63758 28814 63810
rect 28866 63758 28878 63810
rect 30930 63758 30942 63810
rect 30994 63758 31006 63810
rect 33170 63758 33182 63810
rect 33234 63758 33246 63810
rect 27134 63746 27186 63758
rect 32398 63746 32450 63758
rect 50430 63746 50482 63758
rect 50766 63810 50818 63822
rect 50766 63746 50818 63758
rect 54686 63810 54738 63822
rect 54686 63746 54738 63758
rect 13694 63698 13746 63710
rect 13694 63634 13746 63646
rect 43038 63698 43090 63710
rect 43038 63634 43090 63646
rect 43374 63698 43426 63710
rect 43374 63634 43426 63646
rect 55582 63698 55634 63710
rect 55582 63634 55634 63646
rect 55918 63698 55970 63710
rect 55918 63634 55970 63646
rect 1344 63530 58576 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 58576 63530
rect 1344 63444 58576 63478
rect 19630 63362 19682 63374
rect 19630 63298 19682 63310
rect 22318 63362 22370 63374
rect 22318 63298 22370 63310
rect 53566 63362 53618 63374
rect 54450 63310 54462 63362
rect 54514 63310 54526 63362
rect 53566 63298 53618 63310
rect 6638 63250 6690 63262
rect 17502 63250 17554 63262
rect 12898 63198 12910 63250
rect 12962 63198 12974 63250
rect 6638 63186 6690 63198
rect 17502 63186 17554 63198
rect 26238 63250 26290 63262
rect 45166 63250 45218 63262
rect 32050 63198 32062 63250
rect 32114 63198 32126 63250
rect 26238 63186 26290 63198
rect 45166 63186 45218 63198
rect 47742 63250 47794 63262
rect 47742 63186 47794 63198
rect 51438 63250 51490 63262
rect 51438 63186 51490 63198
rect 51662 63250 51714 63262
rect 51662 63186 51714 63198
rect 53006 63250 53058 63262
rect 53006 63186 53058 63198
rect 53902 63250 53954 63262
rect 53902 63186 53954 63198
rect 54910 63250 54962 63262
rect 55234 63198 55246 63250
rect 55298 63198 55310 63250
rect 57362 63198 57374 63250
rect 57426 63198 57438 63250
rect 54910 63186 54962 63198
rect 6750 63138 6802 63150
rect 18062 63138 18114 63150
rect 26686 63138 26738 63150
rect 7858 63086 7870 63138
rect 7922 63086 7934 63138
rect 8082 63086 8094 63138
rect 8146 63086 8158 63138
rect 15474 63086 15486 63138
rect 15538 63086 15550 63138
rect 16258 63086 16270 63138
rect 16322 63086 16334 63138
rect 19618 63086 19630 63138
rect 19682 63086 19694 63138
rect 21298 63086 21310 63138
rect 21362 63086 21374 63138
rect 6750 63074 6802 63086
rect 18062 63074 18114 63086
rect 26686 63074 26738 63086
rect 27134 63138 27186 63150
rect 27806 63138 27858 63150
rect 27570 63086 27582 63138
rect 27634 63086 27646 63138
rect 27134 63074 27186 63086
rect 27806 63074 27858 63086
rect 28142 63138 28194 63150
rect 30382 63138 30434 63150
rect 32622 63138 32674 63150
rect 43486 63138 43538 63150
rect 30146 63086 30158 63138
rect 30210 63086 30222 63138
rect 32274 63086 32286 63138
rect 32338 63086 32350 63138
rect 41234 63086 41246 63138
rect 41298 63086 41310 63138
rect 28142 63074 28194 63086
rect 30382 63074 30434 63086
rect 32622 63074 32674 63086
rect 43486 63074 43538 63086
rect 44046 63138 44098 63150
rect 44046 63074 44098 63086
rect 44942 63138 44994 63150
rect 50654 63138 50706 63150
rect 46050 63086 46062 63138
rect 46114 63086 46126 63138
rect 46498 63086 46510 63138
rect 46562 63086 46574 63138
rect 44942 63074 44994 63086
rect 50654 63074 50706 63086
rect 50766 63138 50818 63150
rect 50766 63074 50818 63086
rect 51102 63138 51154 63150
rect 51102 63074 51154 63086
rect 51214 63138 51266 63150
rect 51214 63074 51266 63086
rect 51774 63138 51826 63150
rect 51774 63074 51826 63086
rect 53230 63138 53282 63150
rect 53230 63074 53282 63086
rect 54126 63138 54178 63150
rect 58146 63086 58158 63138
rect 58210 63086 58222 63138
rect 54126 63074 54178 63086
rect 6526 63026 6578 63038
rect 6526 62962 6578 62974
rect 7086 63026 7138 63038
rect 7086 62962 7138 62974
rect 7646 63026 7698 63038
rect 7646 62962 7698 62974
rect 12574 63026 12626 63038
rect 12574 62962 12626 62974
rect 12798 63026 12850 63038
rect 12798 62962 12850 62974
rect 14814 63026 14866 63038
rect 17614 63026 17666 63038
rect 16370 62974 16382 63026
rect 16434 62974 16446 63026
rect 14814 62962 14866 62974
rect 17614 62962 17666 62974
rect 19966 63026 20018 63038
rect 19966 62962 20018 62974
rect 26126 63026 26178 63038
rect 26126 62962 26178 62974
rect 26462 63026 26514 63038
rect 26462 62962 26514 62974
rect 28030 63026 28082 63038
rect 28030 62962 28082 62974
rect 29486 63026 29538 63038
rect 29486 62962 29538 62974
rect 31166 63026 31218 63038
rect 31166 62962 31218 62974
rect 31278 63026 31330 63038
rect 44158 63026 44210 63038
rect 41010 62974 41022 63026
rect 41074 62974 41086 63026
rect 42242 62974 42254 63026
rect 42306 62974 42318 63026
rect 31278 62962 31330 62974
rect 44158 62962 44210 62974
rect 45054 63026 45106 63038
rect 45054 62962 45106 62974
rect 45502 63026 45554 63038
rect 45502 62962 45554 62974
rect 45838 63026 45890 63038
rect 45838 62962 45890 62974
rect 17390 62914 17442 62926
rect 17390 62850 17442 62862
rect 18510 62914 18562 62926
rect 18510 62850 18562 62862
rect 27022 62914 27074 62926
rect 27022 62850 27074 62862
rect 27246 62914 27298 62926
rect 27246 62850 27298 62862
rect 28590 62914 28642 62926
rect 28590 62850 28642 62862
rect 31502 62914 31554 62926
rect 31502 62850 31554 62862
rect 32062 62914 32114 62926
rect 32062 62850 32114 62862
rect 32958 62914 33010 62926
rect 42926 62914 42978 62926
rect 42466 62862 42478 62914
rect 42530 62862 42542 62914
rect 32958 62850 33010 62862
rect 42926 62850 42978 62862
rect 44382 62914 44434 62926
rect 44382 62850 44434 62862
rect 45278 62914 45330 62926
rect 45278 62850 45330 62862
rect 47182 62914 47234 62926
rect 47182 62850 47234 62862
rect 1344 62746 58576 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 58576 62746
rect 1344 62660 58576 62694
rect 7198 62578 7250 62590
rect 7198 62514 7250 62526
rect 7310 62578 7362 62590
rect 7310 62514 7362 62526
rect 8542 62578 8594 62590
rect 14926 62578 14978 62590
rect 13122 62526 13134 62578
rect 13186 62526 13198 62578
rect 8542 62514 8594 62526
rect 14926 62514 14978 62526
rect 16494 62578 16546 62590
rect 16494 62514 16546 62526
rect 16718 62578 16770 62590
rect 16718 62514 16770 62526
rect 19406 62578 19458 62590
rect 19406 62514 19458 62526
rect 19966 62578 20018 62590
rect 19966 62514 20018 62526
rect 29038 62578 29090 62590
rect 29038 62514 29090 62526
rect 44046 62578 44098 62590
rect 44046 62514 44098 62526
rect 44718 62578 44770 62590
rect 44718 62514 44770 62526
rect 45502 62578 45554 62590
rect 45502 62514 45554 62526
rect 45614 62578 45666 62590
rect 45614 62514 45666 62526
rect 47182 62578 47234 62590
rect 47182 62514 47234 62526
rect 52110 62578 52162 62590
rect 52110 62514 52162 62526
rect 6862 62466 6914 62478
rect 6862 62402 6914 62414
rect 7870 62466 7922 62478
rect 7870 62402 7922 62414
rect 7982 62466 8034 62478
rect 14814 62466 14866 62478
rect 10882 62414 10894 62466
rect 10946 62414 10958 62466
rect 13570 62414 13582 62466
rect 13634 62414 13646 62466
rect 7982 62402 8034 62414
rect 14814 62402 14866 62414
rect 18958 62466 19010 62478
rect 18958 62402 19010 62414
rect 20862 62466 20914 62478
rect 20862 62402 20914 62414
rect 28926 62466 28978 62478
rect 28926 62402 28978 62414
rect 37886 62466 37938 62478
rect 37886 62402 37938 62414
rect 39454 62466 39506 62478
rect 39454 62402 39506 62414
rect 41918 62466 41970 62478
rect 41918 62402 41970 62414
rect 43262 62466 43314 62478
rect 43262 62402 43314 62414
rect 47294 62466 47346 62478
rect 47294 62402 47346 62414
rect 52446 62466 52498 62478
rect 52446 62402 52498 62414
rect 56590 62466 56642 62478
rect 56590 62402 56642 62414
rect 56702 62466 56754 62478
rect 56702 62402 56754 62414
rect 7086 62354 7138 62366
rect 7086 62290 7138 62302
rect 8206 62354 8258 62366
rect 8206 62290 8258 62302
rect 8430 62354 8482 62366
rect 8430 62290 8482 62302
rect 8766 62354 8818 62366
rect 16382 62354 16434 62366
rect 9426 62302 9438 62354
rect 9490 62302 9502 62354
rect 10210 62302 10222 62354
rect 10274 62302 10286 62354
rect 12898 62302 12910 62354
rect 12962 62302 12974 62354
rect 13682 62302 13694 62354
rect 13746 62302 13758 62354
rect 15138 62302 15150 62354
rect 15202 62302 15214 62354
rect 8766 62290 8818 62302
rect 16382 62290 16434 62302
rect 19182 62354 19234 62366
rect 19182 62290 19234 62302
rect 19518 62354 19570 62366
rect 19518 62290 19570 62302
rect 19854 62354 19906 62366
rect 19854 62290 19906 62302
rect 20078 62354 20130 62366
rect 29150 62354 29202 62366
rect 20402 62302 20414 62354
rect 20466 62302 20478 62354
rect 20078 62290 20130 62302
rect 29150 62290 29202 62302
rect 29374 62354 29426 62366
rect 43486 62354 43538 62366
rect 37202 62302 37214 62354
rect 37266 62302 37278 62354
rect 38770 62302 38782 62354
rect 38834 62302 38846 62354
rect 41234 62302 41246 62354
rect 41298 62302 41310 62354
rect 42802 62302 42814 62354
rect 42866 62302 42878 62354
rect 29374 62290 29426 62302
rect 43486 62290 43538 62302
rect 43934 62354 43986 62366
rect 43934 62290 43986 62302
rect 44158 62354 44210 62366
rect 44158 62290 44210 62302
rect 44606 62354 44658 62366
rect 44606 62290 44658 62302
rect 44942 62354 44994 62366
rect 44942 62290 44994 62302
rect 45054 62354 45106 62366
rect 45054 62290 45106 62302
rect 45726 62354 45778 62366
rect 45726 62290 45778 62302
rect 45950 62354 46002 62366
rect 45950 62290 46002 62302
rect 46286 62354 46338 62366
rect 46286 62290 46338 62302
rect 46510 62354 46562 62366
rect 56926 62354 56978 62366
rect 46946 62302 46958 62354
rect 47010 62302 47022 62354
rect 48850 62302 48862 62354
rect 48914 62302 48926 62354
rect 53442 62302 53454 62354
rect 53506 62302 53518 62354
rect 46510 62290 46562 62302
rect 56926 62290 56978 62302
rect 15598 62242 15650 62254
rect 10546 62190 10558 62242
rect 10610 62190 10622 62242
rect 15598 62178 15650 62190
rect 27694 62242 27746 62254
rect 27694 62178 27746 62190
rect 30830 62242 30882 62254
rect 30830 62178 30882 62190
rect 31278 62242 31330 62254
rect 46174 62242 46226 62254
rect 57262 62242 57314 62254
rect 37426 62190 37438 62242
rect 37490 62190 37502 62242
rect 38546 62190 38558 62242
rect 38610 62190 38622 62242
rect 41010 62190 41022 62242
rect 41074 62190 41086 62242
rect 42466 62190 42478 62242
rect 42530 62190 42542 62242
rect 49522 62190 49534 62242
rect 49586 62190 49598 62242
rect 51650 62190 51662 62242
rect 51714 62190 51726 62242
rect 52882 62190 52894 62242
rect 52946 62190 52958 62242
rect 55346 62190 55358 62242
rect 55410 62190 55422 62242
rect 31278 62178 31330 62190
rect 46174 62178 46226 62190
rect 57262 62178 57314 62190
rect 1344 61962 58576 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 58576 61962
rect 1344 61876 58576 61910
rect 20302 61794 20354 61806
rect 20302 61730 20354 61742
rect 43374 61794 43426 61806
rect 43374 61730 43426 61742
rect 49198 61794 49250 61806
rect 49198 61730 49250 61742
rect 56366 61794 56418 61806
rect 56366 61730 56418 61742
rect 12238 61682 12290 61694
rect 36318 61682 36370 61694
rect 24546 61630 24558 61682
rect 24610 61630 24622 61682
rect 35522 61630 35534 61682
rect 35586 61630 35598 61682
rect 12238 61618 12290 61630
rect 36318 61618 36370 61630
rect 37438 61682 37490 61694
rect 37438 61618 37490 61630
rect 38222 61682 38274 61694
rect 52770 61630 52782 61682
rect 52834 61630 52846 61682
rect 55010 61630 55022 61682
rect 55074 61630 55086 61682
rect 38222 61618 38274 61630
rect 21746 61518 21758 61570
rect 21810 61518 21822 61570
rect 38546 61518 38558 61570
rect 38610 61518 38622 61570
rect 43362 61518 43374 61570
rect 43426 61518 43438 61570
rect 53106 61518 53118 61570
rect 53170 61518 53182 61570
rect 54226 61518 54238 61570
rect 54290 61518 54302 61570
rect 55458 61518 55470 61570
rect 55522 61518 55534 61570
rect 6414 61458 6466 61470
rect 6414 61394 6466 61406
rect 6750 61458 6802 61470
rect 6750 61394 6802 61406
rect 19966 61458 20018 61470
rect 24894 61458 24946 61470
rect 20402 61406 20414 61458
rect 20466 61455 20478 61458
rect 20626 61455 20638 61458
rect 20466 61409 20638 61455
rect 20466 61406 20478 61409
rect 20626 61406 20638 61409
rect 20690 61406 20702 61458
rect 22418 61406 22430 61458
rect 22482 61406 22494 61458
rect 19966 61394 20018 61406
rect 24894 61394 24946 61406
rect 32734 61458 32786 61470
rect 32734 61394 32786 61406
rect 34638 61458 34690 61470
rect 34638 61394 34690 61406
rect 35198 61458 35250 61470
rect 35198 61394 35250 61406
rect 36430 61458 36482 61470
rect 36430 61394 36482 61406
rect 36990 61458 37042 61470
rect 36990 61394 37042 61406
rect 37214 61458 37266 61470
rect 37214 61394 37266 61406
rect 37550 61458 37602 61470
rect 37550 61394 37602 61406
rect 43710 61458 43762 61470
rect 43710 61394 43762 61406
rect 49086 61458 49138 61470
rect 49086 61394 49138 61406
rect 6190 61346 6242 61358
rect 6190 61282 6242 61294
rect 6302 61346 6354 61358
rect 6302 61282 6354 61294
rect 6862 61346 6914 61358
rect 6862 61282 6914 61294
rect 7086 61346 7138 61358
rect 7086 61282 7138 61294
rect 7534 61346 7586 61358
rect 7534 61282 7586 61294
rect 20190 61346 20242 61358
rect 20190 61282 20242 61294
rect 20750 61346 20802 61358
rect 20750 61282 20802 61294
rect 25006 61346 25058 61358
rect 25006 61282 25058 61294
rect 25566 61346 25618 61358
rect 25566 61282 25618 61294
rect 25902 61346 25954 61358
rect 25902 61282 25954 61294
rect 32398 61346 32450 61358
rect 32398 61282 32450 61294
rect 32622 61346 32674 61358
rect 32622 61282 32674 61294
rect 34750 61346 34802 61358
rect 34750 61282 34802 61294
rect 34974 61346 35026 61358
rect 34974 61282 35026 61294
rect 35422 61346 35474 61358
rect 35422 61282 35474 61294
rect 36206 61346 36258 61358
rect 36206 61282 36258 61294
rect 38334 61346 38386 61358
rect 38334 61282 38386 61294
rect 44942 61346 44994 61358
rect 44942 61282 44994 61294
rect 1344 61178 58576 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 58576 61178
rect 1344 61092 58576 61126
rect 25454 61010 25506 61022
rect 7858 60958 7870 61010
rect 7922 60958 7934 61010
rect 25454 60946 25506 60958
rect 26014 61010 26066 61022
rect 42702 61010 42754 61022
rect 32274 60958 32286 61010
rect 32338 60958 32350 61010
rect 40002 60958 40014 61010
rect 40066 60958 40078 61010
rect 26014 60946 26066 60958
rect 42702 60946 42754 60958
rect 49086 61010 49138 61022
rect 49086 60946 49138 60958
rect 49646 61010 49698 61022
rect 57934 61010 57986 61022
rect 50978 60958 50990 61010
rect 51042 60958 51054 61010
rect 57026 60958 57038 61010
rect 57090 60958 57102 61010
rect 49646 60946 49698 60958
rect 57934 60946 57986 60958
rect 11006 60898 11058 60910
rect 13246 60898 13298 60910
rect 6290 60846 6302 60898
rect 6354 60846 6366 60898
rect 11890 60846 11902 60898
rect 11954 60846 11966 60898
rect 11006 60834 11058 60846
rect 13246 60834 13298 60846
rect 17502 60898 17554 60910
rect 17502 60834 17554 60846
rect 17950 60898 18002 60910
rect 17950 60834 18002 60846
rect 18062 60898 18114 60910
rect 27246 60898 27298 60910
rect 20962 60846 20974 60898
rect 21026 60846 21038 60898
rect 18062 60834 18114 60846
rect 27246 60834 27298 60846
rect 27806 60898 27858 60910
rect 27806 60834 27858 60846
rect 29598 60898 29650 60910
rect 29598 60834 29650 60846
rect 35422 60898 35474 60910
rect 35422 60834 35474 60846
rect 36766 60898 36818 60910
rect 56590 60898 56642 60910
rect 39106 60846 39118 60898
rect 39170 60846 39182 60898
rect 54450 60846 54462 60898
rect 54514 60846 54526 60898
rect 55794 60846 55806 60898
rect 55858 60846 55870 60898
rect 36766 60834 36818 60846
rect 56590 60834 56642 60846
rect 10782 60786 10834 60798
rect 13022 60786 13074 60798
rect 2818 60734 2830 60786
rect 2882 60734 2894 60786
rect 6738 60734 6750 60786
rect 6802 60734 6814 60786
rect 7522 60734 7534 60786
rect 7586 60734 7598 60786
rect 11554 60734 11566 60786
rect 11618 60734 11630 60786
rect 11778 60734 11790 60786
rect 11842 60734 11854 60786
rect 12786 60734 12798 60786
rect 12850 60734 12862 60786
rect 10782 60722 10834 60734
rect 13022 60722 13074 60734
rect 13358 60786 13410 60798
rect 13358 60722 13410 60734
rect 17390 60786 17442 60798
rect 17390 60722 17442 60734
rect 17726 60786 17778 60798
rect 25902 60786 25954 60798
rect 21746 60734 21758 60786
rect 21810 60734 21822 60786
rect 22642 60734 22654 60786
rect 22706 60734 22718 60786
rect 17726 60722 17778 60734
rect 25902 60722 25954 60734
rect 26238 60786 26290 60798
rect 26238 60722 26290 60734
rect 27134 60786 27186 60798
rect 27134 60722 27186 60734
rect 27470 60786 27522 60798
rect 27470 60722 27522 60734
rect 27694 60786 27746 60798
rect 27694 60722 27746 60734
rect 27918 60786 27970 60798
rect 27918 60722 27970 60734
rect 28366 60786 28418 60798
rect 31950 60786 32002 60798
rect 35870 60786 35922 60798
rect 41358 60786 41410 60798
rect 50094 60786 50146 60798
rect 53006 60786 53058 60798
rect 56926 60786 56978 60798
rect 28914 60734 28926 60786
rect 28978 60734 28990 60786
rect 33394 60734 33406 60786
rect 33458 60734 33470 60786
rect 34738 60734 34750 60786
rect 34802 60734 34814 60786
rect 36082 60734 36094 60786
rect 36146 60734 36158 60786
rect 37762 60734 37774 60786
rect 37826 60734 37838 60786
rect 38994 60734 39006 60786
rect 39058 60734 39070 60786
rect 39890 60734 39902 60786
rect 39954 60734 39966 60786
rect 42466 60734 42478 60786
rect 42530 60734 42542 60786
rect 48850 60734 48862 60786
rect 48914 60734 48926 60786
rect 49298 60734 49310 60786
rect 49362 60734 49374 60786
rect 49634 60734 49646 60786
rect 49698 60734 49710 60786
rect 51202 60734 51214 60786
rect 51266 60734 51278 60786
rect 54674 60734 54686 60786
rect 54738 60734 54750 60786
rect 57250 60734 57262 60786
rect 57314 60734 57326 60786
rect 28366 60722 28418 60734
rect 31950 60722 32002 60734
rect 35870 60722 35922 60734
rect 41358 60722 41410 60734
rect 50094 60722 50146 60734
rect 53006 60722 53058 60734
rect 56926 60722 56978 60734
rect 13918 60674 13970 60686
rect 3490 60622 3502 60674
rect 3554 60622 3566 60674
rect 5618 60622 5630 60674
rect 5682 60622 5694 60674
rect 11106 60622 11118 60674
rect 11170 60622 11182 60674
rect 13918 60610 13970 60622
rect 14254 60674 14306 60686
rect 30046 60674 30098 60686
rect 18834 60622 18846 60674
rect 18898 60622 18910 60674
rect 23202 60622 23214 60674
rect 23266 60622 23278 60674
rect 28690 60622 28702 60674
rect 28754 60622 28766 60674
rect 14254 60610 14306 60622
rect 30046 60610 30098 60622
rect 30494 60674 30546 60686
rect 30494 60610 30546 60622
rect 31614 60674 31666 60686
rect 34078 60674 34130 60686
rect 37326 60674 37378 60686
rect 38558 60674 38610 60686
rect 33170 60622 33182 60674
rect 33234 60622 33246 60674
rect 34514 60622 34526 60674
rect 34578 60622 34590 60674
rect 37986 60622 37998 60674
rect 38050 60622 38062 60674
rect 31614 60610 31666 60622
rect 34078 60610 34130 60622
rect 37326 60610 37378 60622
rect 38558 60610 38610 60622
rect 41022 60674 41074 60686
rect 41022 60610 41074 60622
rect 49758 60674 49810 60686
rect 56030 60674 56082 60686
rect 53330 60622 53342 60674
rect 53394 60622 53406 60674
rect 49758 60610 49810 60622
rect 56030 60610 56082 60622
rect 57822 60674 57874 60686
rect 57822 60610 57874 60622
rect 18062 60562 18114 60574
rect 18062 60498 18114 60510
rect 25230 60562 25282 60574
rect 25230 60498 25282 60510
rect 25566 60562 25618 60574
rect 25566 60498 25618 60510
rect 29934 60562 29986 60574
rect 29934 60498 29986 60510
rect 41470 60562 41522 60574
rect 41470 60498 41522 60510
rect 42814 60562 42866 60574
rect 57710 60562 57762 60574
rect 57138 60510 57150 60562
rect 57202 60510 57214 60562
rect 42814 60498 42866 60510
rect 57710 60498 57762 60510
rect 1344 60394 58576 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 58576 60394
rect 1344 60308 58576 60342
rect 22654 60226 22706 60238
rect 6962 60174 6974 60226
rect 7026 60174 7038 60226
rect 17602 60174 17614 60226
rect 17666 60174 17678 60226
rect 18946 60174 18958 60226
rect 19010 60174 19022 60226
rect 22654 60162 22706 60174
rect 28366 60226 28418 60238
rect 28366 60162 28418 60174
rect 32510 60226 32562 60238
rect 32510 60162 32562 60174
rect 34414 60226 34466 60238
rect 44270 60226 44322 60238
rect 34738 60174 34750 60226
rect 34802 60174 34814 60226
rect 34414 60162 34466 60174
rect 44270 60162 44322 60174
rect 15710 60114 15762 60126
rect 27806 60114 27858 60126
rect 11218 60062 11230 60114
rect 11282 60062 11294 60114
rect 11778 60062 11790 60114
rect 11842 60062 11854 60114
rect 12786 60062 12798 60114
rect 12850 60062 12862 60114
rect 17042 60062 17054 60114
rect 17106 60062 17118 60114
rect 25442 60062 25454 60114
rect 25506 60062 25518 60114
rect 15710 60050 15762 60062
rect 27806 60050 27858 60062
rect 32062 60114 32114 60126
rect 32062 60050 32114 60062
rect 34190 60114 34242 60126
rect 34190 60050 34242 60062
rect 38670 60114 38722 60126
rect 54910 60114 54962 60126
rect 42466 60062 42478 60114
rect 42530 60062 42542 60114
rect 49858 60062 49870 60114
rect 49922 60062 49934 60114
rect 55234 60062 55246 60114
rect 55298 60062 55310 60114
rect 38670 60050 38722 60062
rect 54910 60050 54962 60062
rect 16494 60002 16546 60014
rect 19854 60002 19906 60014
rect 28030 60002 28082 60014
rect 6514 59950 6526 60002
rect 6578 59950 6590 60002
rect 7074 59950 7086 60002
rect 7138 59950 7150 60002
rect 7410 59950 7422 60002
rect 7474 59950 7486 60002
rect 8418 59950 8430 60002
rect 8482 59950 8494 60002
rect 9090 59950 9102 60002
rect 9154 59950 9166 60002
rect 11666 59950 11678 60002
rect 11730 59950 11742 60002
rect 12450 59950 12462 60002
rect 12514 59950 12526 60002
rect 14130 59950 14142 60002
rect 14194 59950 14206 60002
rect 15250 59950 15262 60002
rect 15314 59950 15326 60002
rect 16930 59950 16942 60002
rect 16994 59950 17006 60002
rect 18834 59950 18846 60002
rect 18898 59950 18910 60002
rect 20178 59950 20190 60002
rect 20242 59950 20254 60002
rect 23986 59950 23998 60002
rect 24050 59950 24062 60002
rect 25890 59950 25902 60002
rect 25954 59950 25966 60002
rect 26450 59950 26462 60002
rect 26514 59950 26526 60002
rect 16494 59938 16546 59950
rect 19854 59938 19906 59950
rect 28030 59938 28082 59950
rect 29038 60002 29090 60014
rect 29038 59938 29090 59950
rect 29374 60002 29426 60014
rect 29374 59938 29426 59950
rect 31166 60002 31218 60014
rect 32398 60002 32450 60014
rect 31602 59950 31614 60002
rect 31666 59950 31678 60002
rect 31166 59938 31218 59950
rect 32398 59938 32450 59950
rect 32846 60002 32898 60014
rect 32846 59938 32898 59950
rect 33182 60002 33234 60014
rect 33182 59938 33234 59950
rect 40238 60002 40290 60014
rect 50990 60002 51042 60014
rect 41234 59950 41246 60002
rect 41298 59950 41310 60002
rect 47058 59950 47070 60002
rect 47122 59950 47134 60002
rect 40238 59938 40290 59950
rect 50990 59938 51042 59950
rect 51214 60002 51266 60014
rect 51886 60002 51938 60014
rect 51650 59950 51662 60002
rect 51714 59950 51726 60002
rect 51214 59938 51266 59950
rect 51886 59938 51938 59950
rect 52110 60002 52162 60014
rect 58034 59950 58046 60002
rect 58098 59950 58110 60002
rect 52110 59938 52162 59950
rect 12014 59890 12066 59902
rect 16158 59890 16210 59902
rect 13794 59838 13806 59890
rect 13858 59838 13870 59890
rect 12014 59826 12066 59838
rect 16158 59826 16210 59838
rect 16270 59890 16322 59902
rect 16270 59826 16322 59838
rect 22990 59890 23042 59902
rect 22990 59826 23042 59838
rect 23326 59890 23378 59902
rect 29262 59890 29314 59902
rect 24882 59838 24894 59890
rect 24946 59838 24958 59890
rect 26562 59838 26574 59890
rect 26626 59838 26638 59890
rect 23326 59826 23378 59838
rect 29262 59826 29314 59838
rect 33070 59890 33122 59902
rect 33070 59826 33122 59838
rect 44158 59890 44210 59902
rect 47730 59838 47742 59890
rect 47794 59838 47806 59890
rect 50194 59838 50206 59890
rect 50258 59838 50270 59890
rect 57362 59838 57374 59890
rect 57426 59838 57438 59890
rect 44158 59826 44210 59838
rect 5854 59778 5906 59790
rect 5854 59714 5906 59726
rect 21982 59778 22034 59790
rect 21982 59714 22034 59726
rect 22766 59778 22818 59790
rect 27470 59778 27522 59790
rect 30718 59778 30770 59790
rect 26002 59726 26014 59778
rect 26066 59726 26078 59778
rect 30370 59726 30382 59778
rect 30434 59726 30446 59778
rect 22766 59714 22818 59726
rect 27470 59714 27522 59726
rect 30718 59714 30770 59726
rect 32510 59778 32562 59790
rect 32510 59714 32562 59726
rect 33630 59778 33682 59790
rect 33630 59714 33682 59726
rect 40014 59778 40066 59790
rect 40014 59714 40066 59726
rect 40686 59778 40738 59790
rect 40686 59714 40738 59726
rect 40798 59778 40850 59790
rect 40798 59714 40850 59726
rect 40910 59778 40962 59790
rect 40910 59714 40962 59726
rect 50542 59778 50594 59790
rect 50542 59714 50594 59726
rect 51102 59778 51154 59790
rect 51986 59726 51998 59778
rect 52050 59726 52062 59778
rect 51102 59714 51154 59726
rect 1344 59610 58576 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 58576 59610
rect 1344 59524 58576 59558
rect 7646 59442 7698 59454
rect 7646 59378 7698 59390
rect 11342 59442 11394 59454
rect 11342 59378 11394 59390
rect 15038 59442 15090 59454
rect 15038 59378 15090 59390
rect 15150 59442 15202 59454
rect 42254 59442 42306 59454
rect 15698 59390 15710 59442
rect 15762 59390 15774 59442
rect 16706 59390 16718 59442
rect 16770 59390 16782 59442
rect 27010 59390 27022 59442
rect 27074 59390 27086 59442
rect 15150 59378 15202 59390
rect 42254 59378 42306 59390
rect 48078 59442 48130 59454
rect 48078 59378 48130 59390
rect 48862 59442 48914 59454
rect 48862 59378 48914 59390
rect 48974 59442 49026 59454
rect 48974 59378 49026 59390
rect 49534 59442 49586 59454
rect 49534 59378 49586 59390
rect 50430 59442 50482 59454
rect 50430 59378 50482 59390
rect 54686 59442 54738 59454
rect 54686 59378 54738 59390
rect 56030 59442 56082 59454
rect 56030 59378 56082 59390
rect 56702 59442 56754 59454
rect 56702 59378 56754 59390
rect 7534 59330 7586 59342
rect 7534 59266 7586 59278
rect 7758 59330 7810 59342
rect 7758 59266 7810 59278
rect 8206 59330 8258 59342
rect 40350 59330 40402 59342
rect 17602 59278 17614 59330
rect 17666 59278 17678 59330
rect 37202 59278 37214 59330
rect 37266 59278 37278 59330
rect 8206 59266 8258 59278
rect 40350 59266 40402 59278
rect 40910 59330 40962 59342
rect 40910 59266 40962 59278
rect 41470 59330 41522 59342
rect 41470 59266 41522 59278
rect 42366 59330 42418 59342
rect 42366 59266 42418 59278
rect 43038 59330 43090 59342
rect 43038 59266 43090 59278
rect 48190 59330 48242 59342
rect 48190 59266 48242 59278
rect 56590 59330 56642 59342
rect 56590 59266 56642 59278
rect 56814 59330 56866 59342
rect 56814 59266 56866 59278
rect 14478 59218 14530 59230
rect 12226 59166 12238 59218
rect 12290 59166 12302 59218
rect 14478 59154 14530 59166
rect 14926 59218 14978 59230
rect 14926 59154 14978 59166
rect 16046 59218 16098 59230
rect 16046 59154 16098 59166
rect 16382 59218 16434 59230
rect 35422 59218 35474 59230
rect 17714 59166 17726 59218
rect 17778 59166 17790 59218
rect 27234 59166 27246 59218
rect 27298 59166 27310 59218
rect 16382 59154 16434 59166
rect 35422 59154 35474 59166
rect 35982 59218 36034 59230
rect 41246 59218 41298 59230
rect 42142 59218 42194 59230
rect 42926 59218 42978 59230
rect 39890 59166 39902 59218
rect 39954 59166 39966 59218
rect 41906 59166 41918 59218
rect 41970 59166 41982 59218
rect 42578 59166 42590 59218
rect 42642 59166 42654 59218
rect 35982 59154 36034 59166
rect 41246 59154 41298 59166
rect 42142 59154 42194 59166
rect 42926 59154 42978 59166
rect 43262 59218 43314 59230
rect 45726 59218 45778 59230
rect 45266 59166 45278 59218
rect 45330 59166 45342 59218
rect 43262 59154 43314 59166
rect 45726 59154 45778 59166
rect 49310 59218 49362 59230
rect 49310 59154 49362 59166
rect 49422 59218 49474 59230
rect 49422 59154 49474 59166
rect 49982 59218 50034 59230
rect 58158 59218 58210 59230
rect 51426 59166 51438 59218
rect 51490 59166 51502 59218
rect 49982 59154 50034 59166
rect 58158 59154 58210 59166
rect 1822 59106 1874 59118
rect 27806 59106 27858 59118
rect 12786 59054 12798 59106
rect 12850 59054 12862 59106
rect 18050 59054 18062 59106
rect 18114 59054 18126 59106
rect 1822 59042 1874 59054
rect 27806 59042 27858 59054
rect 30942 59106 30994 59118
rect 30942 59042 30994 59054
rect 32286 59106 32338 59118
rect 41022 59106 41074 59118
rect 36866 59054 36878 59106
rect 36930 59054 36942 59106
rect 39442 59054 39454 59106
rect 39506 59054 39518 59106
rect 32286 59042 32338 59054
rect 41022 59042 41074 59054
rect 49646 59106 49698 59118
rect 52098 59054 52110 59106
rect 52162 59054 52174 59106
rect 54226 59054 54238 59106
rect 54290 59054 54302 59106
rect 57698 59054 57710 59106
rect 57762 59054 57774 59106
rect 49646 59042 49698 59054
rect 35646 58994 35698 59006
rect 35646 58930 35698 58942
rect 44942 58994 44994 59006
rect 44942 58930 44994 58942
rect 45278 58994 45330 59006
rect 45278 58930 45330 58942
rect 1344 58826 58576 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 58576 58826
rect 1344 58740 58576 58774
rect 16718 58658 16770 58670
rect 16718 58594 16770 58606
rect 43150 58658 43202 58670
rect 43150 58594 43202 58606
rect 52110 58658 52162 58670
rect 52110 58594 52162 58606
rect 41806 58546 41858 58558
rect 48190 58546 48242 58558
rect 10210 58494 10222 58546
rect 10274 58494 10286 58546
rect 27570 58494 27582 58546
rect 27634 58494 27646 58546
rect 36194 58494 36206 58546
rect 36258 58494 36270 58546
rect 39218 58494 39230 58546
rect 39282 58494 39294 58546
rect 41346 58494 41358 58546
rect 41410 58494 41422 58546
rect 44818 58494 44830 58546
rect 44882 58494 44894 58546
rect 46946 58494 46958 58546
rect 47010 58494 47022 58546
rect 41806 58482 41858 58494
rect 48190 58482 48242 58494
rect 51998 58546 52050 58558
rect 58270 58546 58322 58558
rect 54674 58494 54686 58546
rect 54738 58494 54750 58546
rect 51998 58482 52050 58494
rect 58270 58482 58322 58494
rect 2270 58434 2322 58446
rect 2270 58370 2322 58382
rect 4062 58434 4114 58446
rect 4062 58370 4114 58382
rect 4286 58434 4338 58446
rect 13806 58434 13858 58446
rect 11778 58382 11790 58434
rect 11842 58382 11854 58434
rect 4286 58370 4338 58382
rect 13806 58370 13858 58382
rect 16382 58434 16434 58446
rect 43262 58434 43314 58446
rect 26674 58382 26686 58434
rect 26738 58382 26750 58434
rect 27458 58382 27470 58434
rect 27522 58382 27534 58434
rect 38546 58382 38558 58434
rect 38610 58382 38622 58434
rect 47730 58382 47742 58434
rect 47794 58382 47806 58434
rect 52994 58382 53006 58434
rect 53058 58382 53070 58434
rect 16382 58370 16434 58382
rect 43262 58370 43314 58382
rect 1710 58322 1762 58334
rect 1710 58258 1762 58270
rect 3838 58322 3890 58334
rect 3838 58258 3890 58270
rect 5630 58322 5682 58334
rect 16158 58322 16210 58334
rect 29822 58322 29874 58334
rect 10658 58270 10670 58322
rect 10722 58270 10734 58322
rect 13458 58270 13470 58322
rect 13522 58270 13534 58322
rect 28130 58270 28142 58322
rect 28194 58270 28206 58322
rect 5630 58258 5682 58270
rect 16158 58258 16210 58270
rect 29822 58258 29874 58270
rect 30494 58322 30546 58334
rect 30494 58258 30546 58270
rect 35982 58322 36034 58334
rect 35982 58258 36034 58270
rect 43150 58322 43202 58334
rect 43150 58258 43202 58270
rect 3950 58210 4002 58222
rect 3950 58146 4002 58158
rect 4846 58210 4898 58222
rect 4846 58146 4898 58158
rect 5742 58210 5794 58222
rect 5742 58146 5794 58158
rect 5966 58210 6018 58222
rect 14478 58210 14530 58222
rect 12002 58158 12014 58210
rect 12066 58158 12078 58210
rect 5966 58146 6018 58158
rect 14478 58146 14530 58158
rect 15374 58210 15426 58222
rect 15374 58146 15426 58158
rect 15822 58210 15874 58222
rect 15822 58146 15874 58158
rect 26574 58210 26626 58222
rect 26574 58146 26626 58158
rect 29934 58210 29986 58222
rect 29934 58146 29986 58158
rect 30046 58210 30098 58222
rect 30046 58146 30098 58158
rect 30606 58210 30658 58222
rect 30606 58146 30658 58158
rect 30830 58210 30882 58222
rect 30830 58146 30882 58158
rect 36206 58210 36258 58222
rect 36206 58146 36258 58158
rect 1344 58042 58576 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 58576 58042
rect 1344 57956 58576 57990
rect 9886 57874 9938 57886
rect 6850 57822 6862 57874
rect 6914 57822 6926 57874
rect 9886 57810 9938 57822
rect 10558 57874 10610 57886
rect 10558 57810 10610 57822
rect 13806 57874 13858 57886
rect 13806 57810 13858 57822
rect 20526 57874 20578 57886
rect 20526 57810 20578 57822
rect 25230 57874 25282 57886
rect 51662 57874 51714 57886
rect 44930 57822 44942 57874
rect 44994 57822 45006 57874
rect 25230 57810 25282 57822
rect 51662 57810 51714 57822
rect 52558 57874 52610 57886
rect 52558 57810 52610 57822
rect 4958 57762 5010 57774
rect 2482 57710 2494 57762
rect 2546 57710 2558 57762
rect 4958 57698 5010 57710
rect 7982 57762 8034 57774
rect 7982 57698 8034 57710
rect 19630 57762 19682 57774
rect 19630 57698 19682 57710
rect 19742 57762 19794 57774
rect 19742 57698 19794 57710
rect 22878 57762 22930 57774
rect 25454 57762 25506 57774
rect 23986 57710 23998 57762
rect 24050 57710 24062 57762
rect 22878 57698 22930 57710
rect 25454 57698 25506 57710
rect 25566 57762 25618 57774
rect 32286 57762 32338 57774
rect 25890 57710 25902 57762
rect 25954 57710 25966 57762
rect 28242 57710 28254 57762
rect 28306 57710 28318 57762
rect 30034 57710 30046 57762
rect 30098 57710 30110 57762
rect 36418 57710 36430 57762
rect 36482 57710 36494 57762
rect 38994 57710 39006 57762
rect 39058 57710 39070 57762
rect 43250 57710 43262 57762
rect 43314 57710 43326 57762
rect 25566 57698 25618 57710
rect 32286 57698 32338 57710
rect 6302 57650 6354 57662
rect 1810 57598 1822 57650
rect 1874 57598 1886 57650
rect 5618 57598 5630 57650
rect 5682 57598 5694 57650
rect 6302 57586 6354 57598
rect 8318 57650 8370 57662
rect 8318 57586 8370 57598
rect 8542 57650 8594 57662
rect 8542 57586 8594 57598
rect 9438 57650 9490 57662
rect 9438 57586 9490 57598
rect 10110 57650 10162 57662
rect 10110 57586 10162 57598
rect 10334 57650 10386 57662
rect 10334 57586 10386 57598
rect 10670 57650 10722 57662
rect 10670 57586 10722 57598
rect 13918 57650 13970 57662
rect 13918 57586 13970 57598
rect 19406 57650 19458 57662
rect 19406 57586 19458 57598
rect 20078 57650 20130 57662
rect 20078 57586 20130 57598
rect 20302 57650 20354 57662
rect 20302 57586 20354 57598
rect 20750 57650 20802 57662
rect 20750 57586 20802 57598
rect 22766 57650 22818 57662
rect 26238 57650 26290 57662
rect 51438 57650 51490 57662
rect 23650 57598 23662 57650
rect 23714 57598 23726 57650
rect 24658 57598 24670 57650
rect 24722 57598 24734 57650
rect 27010 57598 27022 57650
rect 27074 57598 27086 57650
rect 27570 57598 27582 57650
rect 27634 57598 27646 57650
rect 30258 57598 30270 57650
rect 30322 57598 30334 57650
rect 30930 57598 30942 57650
rect 30994 57598 31006 57650
rect 37650 57598 37662 57650
rect 37714 57598 37726 57650
rect 42130 57598 42142 57650
rect 42194 57598 42206 57650
rect 44482 57598 44494 57650
rect 44546 57598 44558 57650
rect 51986 57598 51998 57650
rect 52050 57598 52062 57650
rect 22766 57586 22818 57598
rect 26238 57586 26290 57598
rect 51438 57586 51490 57598
rect 8094 57538 8146 57550
rect 4610 57486 4622 57538
rect 4674 57486 4686 57538
rect 5842 57486 5854 57538
rect 5906 57486 5918 57538
rect 8094 57474 8146 57486
rect 9998 57538 10050 57550
rect 9998 57474 10050 57486
rect 13358 57538 13410 57550
rect 31614 57538 31666 57550
rect 23762 57486 23774 57538
rect 23826 57486 23838 57538
rect 13358 57474 13410 57486
rect 31614 57474 31666 57486
rect 32062 57538 32114 57550
rect 32062 57474 32114 57486
rect 33182 57538 33234 57550
rect 42590 57538 42642 57550
rect 36194 57486 36206 57538
rect 36258 57486 36270 57538
rect 33182 57474 33234 57486
rect 42590 57474 42642 57486
rect 43150 57538 43202 57550
rect 43150 57474 43202 57486
rect 51102 57538 51154 57550
rect 51102 57474 51154 57486
rect 51550 57538 51602 57550
rect 51550 57474 51602 57486
rect 6526 57426 6578 57438
rect 6526 57362 6578 57374
rect 13806 57426 13858 57438
rect 13806 57362 13858 57374
rect 22654 57426 22706 57438
rect 22654 57362 22706 57374
rect 32398 57426 32450 57438
rect 32398 57362 32450 57374
rect 1344 57258 58576 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 58576 57258
rect 1344 57172 58576 57206
rect 12238 57090 12290 57102
rect 12238 57026 12290 57038
rect 24670 57090 24722 57102
rect 24670 57026 24722 57038
rect 27246 57090 27298 57102
rect 43598 57090 43650 57102
rect 29810 57038 29822 57090
rect 29874 57038 29886 57090
rect 27246 57026 27298 57038
rect 43598 57026 43650 57038
rect 4398 56978 4450 56990
rect 4398 56914 4450 56926
rect 6078 56978 6130 56990
rect 14142 56978 14194 56990
rect 7410 56926 7422 56978
rect 7474 56926 7486 56978
rect 9538 56926 9550 56978
rect 9602 56926 9614 56978
rect 10658 56926 10670 56978
rect 10722 56926 10734 56978
rect 6078 56914 6130 56926
rect 14142 56914 14194 56926
rect 15038 56978 15090 56990
rect 15038 56914 15090 56926
rect 16158 56978 16210 56990
rect 20190 56978 20242 56990
rect 34974 56978 35026 56990
rect 19394 56926 19406 56978
rect 19458 56926 19470 56978
rect 22082 56926 22094 56978
rect 22146 56926 22158 56978
rect 24210 56926 24222 56978
rect 24274 56926 24286 56978
rect 29922 56926 29934 56978
rect 29986 56926 29998 56978
rect 31602 56926 31614 56978
rect 31666 56926 31678 56978
rect 33730 56926 33742 56978
rect 33794 56926 33806 56978
rect 16158 56914 16210 56926
rect 20190 56914 20242 56926
rect 34974 56914 35026 56926
rect 36318 56978 36370 56990
rect 36318 56914 36370 56926
rect 42366 56978 42418 56990
rect 42366 56914 42418 56926
rect 42702 56978 42754 56990
rect 50430 56978 50482 56990
rect 47058 56926 47070 56978
rect 47122 56926 47134 56978
rect 55346 56926 55358 56978
rect 55410 56926 55422 56978
rect 42702 56914 42754 56926
rect 50430 56914 50482 56926
rect 4510 56866 4562 56878
rect 4510 56802 4562 56814
rect 4958 56866 5010 56878
rect 4958 56802 5010 56814
rect 5518 56866 5570 56878
rect 5518 56802 5570 56814
rect 5966 56866 6018 56878
rect 20302 56866 20354 56878
rect 6738 56814 6750 56866
rect 6802 56814 6814 56866
rect 10546 56814 10558 56866
rect 10610 56814 10622 56866
rect 14578 56814 14590 56866
rect 14642 56814 14654 56866
rect 16482 56814 16494 56866
rect 16546 56814 16558 56866
rect 5966 56802 6018 56814
rect 20302 56802 20354 56814
rect 20750 56866 20802 56878
rect 25454 56866 25506 56878
rect 26686 56866 26738 56878
rect 35982 56866 36034 56878
rect 21298 56814 21310 56866
rect 21362 56814 21374 56866
rect 26114 56814 26126 56866
rect 26178 56814 26190 56866
rect 30146 56814 30158 56866
rect 30210 56814 30222 56866
rect 30818 56814 30830 56866
rect 30882 56814 30894 56866
rect 34514 56814 34526 56866
rect 34578 56814 34590 56866
rect 20750 56802 20802 56814
rect 25454 56802 25506 56814
rect 26686 56802 26738 56814
rect 35982 56802 36034 56814
rect 37102 56866 37154 56878
rect 37998 56866 38050 56878
rect 37314 56814 37326 56866
rect 37378 56814 37390 56866
rect 37102 56802 37154 56814
rect 37998 56802 38050 56814
rect 42254 56866 42306 56878
rect 42254 56802 42306 56814
rect 42926 56866 42978 56878
rect 49970 56814 49982 56866
rect 50034 56814 50046 56866
rect 42926 56802 42978 56814
rect 4286 56754 4338 56766
rect 4286 56690 4338 56702
rect 9886 56754 9938 56766
rect 9886 56690 9938 56702
rect 12014 56754 12066 56766
rect 13918 56754 13970 56766
rect 13794 56702 13806 56754
rect 13858 56702 13870 56754
rect 12014 56690 12066 56702
rect 13918 56690 13970 56702
rect 14254 56754 14306 56766
rect 14254 56690 14306 56702
rect 15150 56754 15202 56766
rect 19854 56754 19906 56766
rect 17266 56702 17278 56754
rect 17330 56702 17342 56754
rect 15150 56690 15202 56702
rect 19854 56690 19906 56702
rect 24782 56754 24834 56766
rect 26798 56754 26850 56766
rect 25106 56702 25118 56754
rect 25170 56702 25182 56754
rect 24782 56690 24834 56702
rect 26798 56690 26850 56702
rect 27134 56754 27186 56766
rect 27134 56690 27186 56702
rect 36094 56754 36146 56766
rect 36094 56690 36146 56702
rect 36430 56754 36482 56766
rect 36430 56690 36482 56702
rect 42478 56754 42530 56766
rect 42478 56690 42530 56702
rect 43262 56754 43314 56766
rect 43262 56690 43314 56702
rect 43486 56754 43538 56766
rect 55582 56754 55634 56766
rect 49186 56702 49198 56754
rect 49250 56702 49262 56754
rect 43486 56690 43538 56702
rect 55582 56690 55634 56702
rect 6190 56642 6242 56654
rect 14030 56642 14082 56654
rect 12562 56590 12574 56642
rect 12626 56590 12638 56642
rect 6190 56578 6242 56590
rect 14030 56578 14082 56590
rect 14926 56642 14978 56654
rect 14926 56578 14978 56590
rect 20078 56642 20130 56654
rect 20078 56578 20130 56590
rect 24670 56642 24722 56654
rect 24670 56578 24722 56590
rect 27694 56642 27746 56654
rect 27694 56578 27746 56590
rect 55358 56642 55410 56654
rect 55358 56578 55410 56590
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 8654 56306 8706 56318
rect 8654 56242 8706 56254
rect 8766 56306 8818 56318
rect 8766 56242 8818 56254
rect 9774 56306 9826 56318
rect 13694 56306 13746 56318
rect 10770 56254 10782 56306
rect 10834 56254 10846 56306
rect 11218 56254 11230 56306
rect 11282 56254 11294 56306
rect 12114 56254 12126 56306
rect 12178 56254 12190 56306
rect 9774 56242 9826 56254
rect 13694 56242 13746 56254
rect 14590 56306 14642 56318
rect 28478 56306 28530 56318
rect 22642 56254 22654 56306
rect 22706 56254 22718 56306
rect 14590 56242 14642 56254
rect 28478 56242 28530 56254
rect 46958 56306 47010 56318
rect 46958 56242 47010 56254
rect 48190 56306 48242 56318
rect 48190 56242 48242 56254
rect 48862 56306 48914 56318
rect 54238 56306 54290 56318
rect 49970 56254 49982 56306
rect 50034 56254 50046 56306
rect 48862 56242 48914 56254
rect 54238 56242 54290 56254
rect 8318 56194 8370 56206
rect 8318 56130 8370 56142
rect 12910 56194 12962 56206
rect 12910 56130 12962 56142
rect 13134 56194 13186 56206
rect 13134 56130 13186 56142
rect 13358 56194 13410 56206
rect 13358 56130 13410 56142
rect 13470 56194 13522 56206
rect 13470 56130 13522 56142
rect 13918 56194 13970 56206
rect 13918 56130 13970 56142
rect 14030 56194 14082 56206
rect 14030 56130 14082 56142
rect 17950 56194 18002 56206
rect 48750 56194 48802 56206
rect 19058 56142 19070 56194
rect 19122 56142 19134 56194
rect 20290 56142 20302 56194
rect 20354 56142 20366 56194
rect 23874 56142 23886 56194
rect 23938 56142 23950 56194
rect 31826 56142 31838 56194
rect 31890 56142 31902 56194
rect 32498 56142 32510 56194
rect 32562 56142 32574 56194
rect 35186 56142 35198 56194
rect 35250 56142 35262 56194
rect 35634 56142 35646 56194
rect 35698 56142 35710 56194
rect 37314 56142 37326 56194
rect 37378 56142 37390 56194
rect 51650 56142 51662 56194
rect 51714 56142 51726 56194
rect 17950 56130 18002 56142
rect 48750 56130 48802 56142
rect 8542 56082 8594 56094
rect 8542 56018 8594 56030
rect 10222 56082 10274 56094
rect 10222 56018 10274 56030
rect 10446 56082 10498 56094
rect 10446 56018 10498 56030
rect 11566 56082 11618 56094
rect 11566 56018 11618 56030
rect 12462 56082 12514 56094
rect 12462 56018 12514 56030
rect 12798 56082 12850 56094
rect 12798 56018 12850 56030
rect 14254 56082 14306 56094
rect 38222 56082 38274 56094
rect 47070 56082 47122 56094
rect 15138 56030 15150 56082
rect 15202 56030 15214 56082
rect 22978 56030 22990 56082
rect 23042 56030 23054 56082
rect 32274 56030 32286 56082
rect 32338 56030 32350 56082
rect 33618 56030 33630 56082
rect 33682 56030 33694 56082
rect 34178 56030 34190 56082
rect 34242 56030 34254 56082
rect 35858 56030 35870 56082
rect 35922 56030 35934 56082
rect 37202 56030 37214 56082
rect 37266 56030 37278 56082
rect 38994 56030 39006 56082
rect 39058 56030 39070 56082
rect 14254 56018 14306 56030
rect 38222 56018 38274 56030
rect 47070 56018 47122 56030
rect 47182 56082 47234 56094
rect 48078 56082 48130 56094
rect 47618 56030 47630 56082
rect 47682 56030 47694 56082
rect 47182 56018 47234 56030
rect 48078 56018 48130 56030
rect 50318 56082 50370 56094
rect 50866 56030 50878 56082
rect 50930 56030 50942 56082
rect 54898 56030 54910 56082
rect 54962 56030 54974 56082
rect 50318 56018 50370 56030
rect 4510 55970 4562 55982
rect 4510 55906 4562 55918
rect 5070 55970 5122 55982
rect 18174 55970 18226 55982
rect 15250 55918 15262 55970
rect 15314 55918 15326 55970
rect 17826 55918 17838 55970
rect 17890 55918 17902 55970
rect 5070 55906 5122 55918
rect 18174 55906 18226 55918
rect 18734 55970 18786 55982
rect 18734 55906 18786 55918
rect 20750 55970 20802 55982
rect 25342 55970 25394 55982
rect 24434 55918 24446 55970
rect 24498 55918 24510 55970
rect 20750 55906 20802 55918
rect 25342 55906 25394 55918
rect 31390 55970 31442 55982
rect 31390 55906 31442 55918
rect 45502 55970 45554 55982
rect 45502 55906 45554 55918
rect 47854 55970 47906 55982
rect 53778 55918 53790 55970
rect 53842 55918 53854 55970
rect 55122 55918 55134 55970
rect 55186 55918 55198 55970
rect 47854 55906 47906 55918
rect 45614 55858 45666 55870
rect 15922 55806 15934 55858
rect 15986 55806 15998 55858
rect 55570 55806 55582 55858
rect 55634 55806 55646 55858
rect 45614 55794 45666 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 4734 55522 4786 55534
rect 4734 55458 4786 55470
rect 23550 55522 23602 55534
rect 23550 55458 23602 55470
rect 32286 55522 32338 55534
rect 43150 55522 43202 55534
rect 35186 55470 35198 55522
rect 35250 55470 35262 55522
rect 32286 55458 32338 55470
rect 43150 55458 43202 55470
rect 11790 55410 11842 55422
rect 23762 55358 23774 55410
rect 23826 55358 23838 55410
rect 33170 55358 33182 55410
rect 33234 55358 33246 55410
rect 34850 55358 34862 55410
rect 34914 55358 34926 55410
rect 40450 55358 40462 55410
rect 40514 55358 40526 55410
rect 41570 55358 41582 55410
rect 41634 55358 41646 55410
rect 42130 55358 42142 55410
rect 42194 55358 42206 55410
rect 45602 55358 45614 55410
rect 45666 55358 45678 55410
rect 47730 55358 47742 55410
rect 47794 55358 47806 55410
rect 52770 55358 52782 55410
rect 52834 55358 52846 55410
rect 55570 55358 55582 55410
rect 55634 55358 55646 55410
rect 57698 55358 57710 55410
rect 57762 55358 57774 55410
rect 11790 55346 11842 55358
rect 3390 55298 3442 55310
rect 3390 55234 3442 55246
rect 3838 55298 3890 55310
rect 3838 55234 3890 55246
rect 4398 55298 4450 55310
rect 4398 55234 4450 55246
rect 11006 55298 11058 55310
rect 11006 55234 11058 55246
rect 11342 55298 11394 55310
rect 11342 55234 11394 55246
rect 14478 55298 14530 55310
rect 28366 55298 28418 55310
rect 31726 55298 31778 55310
rect 33854 55298 33906 55310
rect 42814 55298 42866 55310
rect 58158 55298 58210 55310
rect 23874 55246 23886 55298
rect 23938 55246 23950 55298
rect 29250 55246 29262 55298
rect 29314 55246 29326 55298
rect 30146 55246 30158 55298
rect 30210 55246 30222 55298
rect 32946 55246 32958 55298
rect 33010 55246 33022 55298
rect 34738 55246 34750 55298
rect 34802 55246 34814 55298
rect 37650 55246 37662 55298
rect 37714 55246 37726 55298
rect 41458 55246 41470 55298
rect 41522 55246 41534 55298
rect 42354 55246 42366 55298
rect 42418 55246 42430 55298
rect 44930 55246 44942 55298
rect 44994 55246 45006 55298
rect 53330 55246 53342 55298
rect 53394 55246 53406 55298
rect 54898 55246 54910 55298
rect 54962 55246 54974 55298
rect 14478 55234 14530 55246
rect 28366 55234 28418 55246
rect 31726 55234 31778 55246
rect 33854 55234 33906 55246
rect 42814 55234 42866 55246
rect 58158 55234 58210 55246
rect 2830 55186 2882 55198
rect 2830 55122 2882 55134
rect 3166 55186 3218 55198
rect 3166 55122 3218 55134
rect 4846 55186 4898 55198
rect 31390 55186 31442 55198
rect 29362 55134 29374 55186
rect 29426 55134 29438 55186
rect 30706 55134 30718 55186
rect 30770 55134 30782 55186
rect 4846 55122 4898 55134
rect 31390 55122 31442 55134
rect 31502 55186 31554 55198
rect 31502 55122 31554 55134
rect 32286 55186 32338 55198
rect 32286 55122 32338 55134
rect 32398 55186 32450 55198
rect 40798 55186 40850 55198
rect 38322 55134 38334 55186
rect 38386 55134 38398 55186
rect 49970 55134 49982 55186
rect 50034 55134 50046 55186
rect 32398 55122 32450 55134
rect 40798 55122 40850 55134
rect 2942 55074 2994 55086
rect 2942 55010 2994 55022
rect 3726 55074 3778 55086
rect 3726 55010 3778 55022
rect 3950 55074 4002 55086
rect 3950 55010 4002 55022
rect 4734 55074 4786 55086
rect 4734 55010 4786 55022
rect 11118 55074 11170 55086
rect 11118 55010 11170 55022
rect 12686 55074 12738 55086
rect 12686 55010 12738 55022
rect 13582 55074 13634 55086
rect 13582 55010 13634 55022
rect 14590 55074 14642 55086
rect 14590 55010 14642 55022
rect 18398 55074 18450 55086
rect 18398 55010 18450 55022
rect 27694 55074 27746 55086
rect 27694 55010 27746 55022
rect 27806 55074 27858 55086
rect 27806 55010 27858 55022
rect 27918 55074 27970 55086
rect 31054 55074 31106 55086
rect 30146 55022 30158 55074
rect 30210 55022 30222 55074
rect 27918 55010 27970 55022
rect 31054 55010 31106 55022
rect 43038 55074 43090 55086
rect 43038 55010 43090 55022
rect 44270 55074 44322 55086
rect 49534 55074 49586 55086
rect 49186 55022 49198 55074
rect 49250 55022 49262 55074
rect 44270 55010 44322 55022
rect 49534 55010 49586 55022
rect 50318 55074 50370 55086
rect 50318 55010 50370 55022
rect 52782 55074 52834 55086
rect 52782 55010 52834 55022
rect 52894 55074 52946 55086
rect 52894 55010 52946 55022
rect 53118 55074 53170 55086
rect 53118 55010 53170 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 5070 54738 5122 54750
rect 14590 54738 14642 54750
rect 39566 54738 39618 54750
rect 10994 54686 11006 54738
rect 11058 54686 11070 54738
rect 29474 54686 29486 54738
rect 29538 54686 29550 54738
rect 5070 54674 5122 54686
rect 14590 54674 14642 54686
rect 39566 54674 39618 54686
rect 41022 54738 41074 54750
rect 41022 54674 41074 54686
rect 41582 54738 41634 54750
rect 41582 54674 41634 54686
rect 41694 54738 41746 54750
rect 41694 54674 41746 54686
rect 41806 54738 41858 54750
rect 41806 54674 41858 54686
rect 42478 54738 42530 54750
rect 42478 54674 42530 54686
rect 45502 54738 45554 54750
rect 45502 54674 45554 54686
rect 45950 54738 46002 54750
rect 45950 54674 46002 54686
rect 46622 54738 46674 54750
rect 51874 54686 51886 54738
rect 51938 54686 51950 54738
rect 46622 54674 46674 54686
rect 5406 54626 5458 54638
rect 2482 54574 2494 54626
rect 2546 54574 2558 54626
rect 5406 54562 5458 54574
rect 26686 54626 26738 54638
rect 26686 54562 26738 54574
rect 27022 54626 27074 54638
rect 27022 54562 27074 54574
rect 31502 54626 31554 54638
rect 31502 54562 31554 54574
rect 39454 54626 39506 54638
rect 39454 54562 39506 54574
rect 39790 54626 39842 54638
rect 39790 54562 39842 54574
rect 42366 54626 42418 54638
rect 55806 54626 55858 54638
rect 51202 54574 51214 54626
rect 51266 54574 51278 54626
rect 42366 54562 42418 54574
rect 55806 54562 55858 54574
rect 4958 54514 5010 54526
rect 1810 54462 1822 54514
rect 1874 54462 1886 54514
rect 4958 54450 5010 54462
rect 5182 54514 5234 54526
rect 5182 54450 5234 54462
rect 11342 54514 11394 54526
rect 11342 54450 11394 54462
rect 14254 54514 14306 54526
rect 14254 54450 14306 54462
rect 14478 54514 14530 54526
rect 14478 54450 14530 54462
rect 14814 54514 14866 54526
rect 14814 54450 14866 54462
rect 15150 54514 15202 54526
rect 18286 54514 18338 54526
rect 15362 54462 15374 54514
rect 15426 54462 15438 54514
rect 15150 54450 15202 54462
rect 18286 54450 18338 54462
rect 27246 54514 27298 54526
rect 27246 54450 27298 54462
rect 27582 54514 27634 54526
rect 39902 54514 39954 54526
rect 28130 54462 28142 54514
rect 28194 54462 28206 54514
rect 31042 54462 31054 54514
rect 31106 54462 31118 54514
rect 27582 54450 27634 54462
rect 39902 54450 39954 54462
rect 41470 54514 41522 54526
rect 46062 54514 46114 54526
rect 42018 54462 42030 54514
rect 42082 54462 42094 54514
rect 41470 54450 41522 54462
rect 46062 54450 46114 54462
rect 46398 54514 46450 54526
rect 50878 54514 50930 54526
rect 56478 54514 56530 54526
rect 46610 54462 46622 54514
rect 46674 54462 46686 54514
rect 51650 54462 51662 54514
rect 51714 54462 51726 54514
rect 46398 54450 46450 54462
rect 50878 54450 50930 54462
rect 56478 54450 56530 54462
rect 56814 54514 56866 54526
rect 56814 54450 56866 54462
rect 57150 54514 57202 54526
rect 57150 54450 57202 54462
rect 16046 54402 16098 54414
rect 4610 54350 4622 54402
rect 4674 54350 4686 54402
rect 16046 54338 16098 54350
rect 26798 54402 26850 54414
rect 28926 54402 28978 54414
rect 28466 54350 28478 54402
rect 28530 54350 28542 54402
rect 26798 54338 26850 54350
rect 28926 54338 28978 54350
rect 29150 54402 29202 54414
rect 31950 54402 32002 54414
rect 30594 54350 30606 54402
rect 30658 54350 30670 54402
rect 29150 54338 29202 54350
rect 31950 54338 32002 54350
rect 32510 54402 32562 54414
rect 32510 54338 32562 54350
rect 33182 54402 33234 54414
rect 33182 54338 33234 54350
rect 46846 54402 46898 54414
rect 46846 54338 46898 54350
rect 47182 54402 47234 54414
rect 47182 54338 47234 54350
rect 55134 54402 55186 54414
rect 55134 54338 55186 54350
rect 55918 54402 55970 54414
rect 55918 54338 55970 54350
rect 56702 54402 56754 54414
rect 56702 54338 56754 54350
rect 54910 54290 54962 54302
rect 54562 54238 54574 54290
rect 54626 54238 54638 54290
rect 54910 54226 54962 54238
rect 56030 54290 56082 54302
rect 56030 54226 56082 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 8990 53954 9042 53966
rect 8990 53890 9042 53902
rect 23326 53954 23378 53966
rect 23326 53890 23378 53902
rect 29374 53954 29426 53966
rect 29374 53890 29426 53902
rect 29710 53954 29762 53966
rect 52670 53954 52722 53966
rect 36306 53902 36318 53954
rect 36370 53902 36382 53954
rect 29710 53890 29762 53902
rect 52670 53890 52722 53902
rect 2942 53842 2994 53854
rect 2942 53778 2994 53790
rect 5070 53842 5122 53854
rect 5070 53778 5122 53790
rect 18734 53842 18786 53854
rect 29150 53842 29202 53854
rect 39902 53842 39954 53854
rect 22306 53790 22318 53842
rect 22370 53790 22382 53842
rect 24098 53790 24110 53842
rect 24162 53790 24174 53842
rect 26002 53790 26014 53842
rect 26066 53790 26078 53842
rect 28130 53790 28142 53842
rect 28194 53790 28206 53842
rect 36082 53790 36094 53842
rect 36146 53790 36158 53842
rect 37090 53790 37102 53842
rect 37154 53790 37166 53842
rect 18734 53778 18786 53790
rect 29150 53778 29202 53790
rect 39902 53778 39954 53790
rect 53006 53842 53058 53854
rect 53006 53778 53058 53790
rect 53902 53842 53954 53854
rect 56018 53790 56030 53842
rect 56082 53790 56094 53842
rect 58146 53790 58158 53842
rect 58210 53790 58222 53842
rect 53902 53778 53954 53790
rect 3838 53730 3890 53742
rect 3378 53678 3390 53730
rect 3442 53678 3454 53730
rect 3838 53666 3890 53678
rect 4622 53730 4674 53742
rect 4622 53666 4674 53678
rect 8430 53730 8482 53742
rect 8430 53666 8482 53678
rect 8878 53730 8930 53742
rect 8878 53666 8930 53678
rect 17838 53730 17890 53742
rect 17838 53666 17890 53678
rect 18398 53730 18450 53742
rect 18398 53666 18450 53678
rect 19854 53730 19906 53742
rect 19854 53666 19906 53678
rect 19966 53730 20018 53742
rect 37998 53730 38050 53742
rect 23874 53678 23886 53730
rect 23938 53678 23950 53730
rect 24770 53678 24782 53730
rect 24834 53678 24846 53730
rect 25330 53678 25342 53730
rect 25394 53678 25406 53730
rect 34514 53678 34526 53730
rect 34578 53678 34590 53730
rect 35970 53678 35982 53730
rect 36034 53678 36046 53730
rect 37314 53678 37326 53730
rect 37378 53678 37390 53730
rect 19966 53666 20018 53678
rect 37998 53666 38050 53678
rect 39790 53730 39842 53742
rect 39790 53666 39842 53678
rect 40014 53730 40066 53742
rect 51426 53678 51438 53730
rect 51490 53678 51502 53730
rect 54898 53678 54910 53730
rect 54962 53678 54974 53730
rect 55234 53678 55246 53730
rect 55298 53678 55310 53730
rect 40014 53666 40066 53678
rect 4286 53618 4338 53630
rect 4286 53554 4338 53566
rect 4398 53618 4450 53630
rect 4398 53554 4450 53566
rect 7086 53618 7138 53630
rect 7086 53554 7138 53566
rect 7422 53618 7474 53630
rect 7422 53554 7474 53566
rect 7646 53618 7698 53630
rect 17950 53618 18002 53630
rect 10322 53566 10334 53618
rect 10386 53566 10398 53618
rect 7646 53554 7698 53566
rect 17950 53554 18002 53566
rect 19070 53618 19122 53630
rect 19070 53554 19122 53566
rect 20638 53618 20690 53630
rect 20638 53554 20690 53566
rect 22654 53618 22706 53630
rect 22654 53554 22706 53566
rect 23102 53618 23154 53630
rect 40238 53618 40290 53630
rect 24322 53566 24334 53618
rect 24386 53566 24398 53618
rect 30370 53566 30382 53618
rect 30434 53566 30446 53618
rect 23102 53554 23154 53566
rect 40238 53554 40290 53566
rect 40910 53618 40962 53630
rect 40910 53554 40962 53566
rect 41246 53618 41298 53630
rect 41246 53554 41298 53566
rect 41582 53618 41634 53630
rect 41582 53554 41634 53566
rect 41694 53618 41746 53630
rect 54226 53566 54238 53618
rect 54290 53566 54302 53618
rect 54786 53566 54798 53618
rect 54850 53566 54862 53618
rect 41694 53554 41746 53566
rect 7198 53506 7250 53518
rect 7198 53442 7250 53454
rect 8094 53506 8146 53518
rect 8094 53442 8146 53454
rect 8318 53506 8370 53518
rect 8318 53442 8370 53454
rect 8542 53506 8594 53518
rect 8542 53442 8594 53454
rect 8990 53506 9042 53518
rect 8990 53442 9042 53454
rect 10670 53506 10722 53518
rect 10670 53442 10722 53454
rect 18174 53506 18226 53518
rect 18174 53442 18226 53454
rect 18622 53506 18674 53518
rect 18622 53442 18674 53454
rect 18846 53506 18898 53518
rect 18846 53442 18898 53454
rect 19630 53506 19682 53518
rect 19630 53442 19682 53454
rect 20078 53506 20130 53518
rect 20078 53442 20130 53454
rect 20302 53506 20354 53518
rect 20302 53442 20354 53454
rect 20526 53506 20578 53518
rect 20526 53442 20578 53454
rect 22430 53506 22482 53518
rect 22430 53442 22482 53454
rect 23214 53506 23266 53518
rect 23214 53442 23266 53454
rect 30046 53506 30098 53518
rect 30046 53442 30098 53454
rect 33182 53506 33234 53518
rect 33182 53442 33234 53454
rect 39566 53506 39618 53518
rect 39566 53442 39618 53454
rect 41022 53506 41074 53518
rect 41022 53442 41074 53454
rect 41358 53506 41410 53518
rect 52782 53506 52834 53518
rect 51650 53454 51662 53506
rect 51714 53454 51726 53506
rect 41358 53442 41410 53454
rect 52782 53442 52834 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 8542 53170 8594 53182
rect 14590 53170 14642 53182
rect 13122 53118 13134 53170
rect 13186 53118 13198 53170
rect 8542 53106 8594 53118
rect 14590 53106 14642 53118
rect 23998 53170 24050 53182
rect 23998 53106 24050 53118
rect 24670 53170 24722 53182
rect 24670 53106 24722 53118
rect 25342 53170 25394 53182
rect 25342 53106 25394 53118
rect 31278 53170 31330 53182
rect 31278 53106 31330 53118
rect 36430 53170 36482 53182
rect 36430 53106 36482 53118
rect 41022 53170 41074 53182
rect 41022 53106 41074 53118
rect 45838 53170 45890 53182
rect 45838 53106 45890 53118
rect 46622 53170 46674 53182
rect 46622 53106 46674 53118
rect 46846 53170 46898 53182
rect 46846 53106 46898 53118
rect 47518 53170 47570 53182
rect 47518 53106 47570 53118
rect 47966 53170 48018 53182
rect 47966 53106 48018 53118
rect 55022 53170 55074 53182
rect 55022 53106 55074 53118
rect 12014 53058 12066 53070
rect 5954 53006 5966 53058
rect 6018 53006 6030 53058
rect 12014 52994 12066 53006
rect 12574 53058 12626 53070
rect 12574 52994 12626 53006
rect 14814 53058 14866 53070
rect 23886 53058 23938 53070
rect 18162 53006 18174 53058
rect 18226 53006 18238 53058
rect 21410 53006 21422 53058
rect 21474 53006 21486 53058
rect 14814 52994 14866 53006
rect 23886 52994 23938 53006
rect 36206 53058 36258 53070
rect 36206 52994 36258 53006
rect 36654 53058 36706 53070
rect 51538 53006 51550 53058
rect 51602 53006 51614 53058
rect 36654 52994 36706 53006
rect 8430 52946 8482 52958
rect 5282 52894 5294 52946
rect 5346 52894 5358 52946
rect 8430 52882 8482 52894
rect 8654 52946 8706 52958
rect 8654 52882 8706 52894
rect 9102 52946 9154 52958
rect 12686 52946 12738 52958
rect 11554 52894 11566 52946
rect 11618 52894 11630 52946
rect 12338 52894 12350 52946
rect 12402 52894 12414 52946
rect 9102 52882 9154 52894
rect 12686 52882 12738 52894
rect 14926 52946 14978 52958
rect 32174 52946 32226 52958
rect 34414 52946 34466 52958
rect 36766 52946 36818 52958
rect 54126 52946 54178 52958
rect 17490 52894 17502 52946
rect 17554 52894 17566 52946
rect 20626 52894 20638 52946
rect 20690 52894 20702 52946
rect 24210 52894 24222 52946
rect 24274 52894 24286 52946
rect 31490 52894 31502 52946
rect 31554 52894 31566 52946
rect 33730 52894 33742 52946
rect 33794 52894 33806 52946
rect 35634 52894 35646 52946
rect 35698 52894 35710 52946
rect 35970 52894 35982 52946
rect 36034 52894 36046 52946
rect 42466 52894 42478 52946
rect 42530 52894 42542 52946
rect 46386 52894 46398 52946
rect 46450 52894 46462 52946
rect 47058 52894 47070 52946
rect 47122 52894 47134 52946
rect 50754 52894 50766 52946
rect 50818 52894 50830 52946
rect 14926 52882 14978 52894
rect 32174 52882 32226 52894
rect 34414 52882 34466 52894
rect 36766 52882 36818 52894
rect 54126 52882 54178 52894
rect 54462 52946 54514 52958
rect 54462 52882 54514 52894
rect 58158 52946 58210 52958
rect 58158 52882 58210 52894
rect 9774 52834 9826 52846
rect 8082 52782 8094 52834
rect 8146 52782 8158 52834
rect 9774 52770 9826 52782
rect 10110 52834 10162 52846
rect 10110 52770 10162 52782
rect 10670 52834 10722 52846
rect 13694 52834 13746 52846
rect 31950 52834 32002 52846
rect 57374 52834 57426 52846
rect 11106 52782 11118 52834
rect 11170 52782 11182 52834
rect 20290 52782 20302 52834
rect 20354 52782 20366 52834
rect 23538 52782 23550 52834
rect 23602 52782 23614 52834
rect 33506 52782 33518 52834
rect 33570 52782 33582 52834
rect 43250 52782 43262 52834
rect 43314 52782 43326 52834
rect 45378 52782 45390 52834
rect 45442 52782 45454 52834
rect 46498 52782 46510 52834
rect 46562 52782 46574 52834
rect 53666 52782 53678 52834
rect 53730 52782 53742 52834
rect 10670 52770 10722 52782
rect 13694 52770 13746 52782
rect 31950 52770 32002 52782
rect 57374 52770 57426 52782
rect 57598 52834 57650 52846
rect 57598 52770 57650 52782
rect 10334 52722 10386 52734
rect 54014 52722 54066 52734
rect 32498 52670 32510 52722
rect 32562 52670 32574 52722
rect 45602 52670 45614 52722
rect 45666 52719 45678 52722
rect 46162 52719 46174 52722
rect 45666 52673 46174 52719
rect 45666 52670 45678 52673
rect 46162 52670 46174 52673
rect 46226 52670 46238 52722
rect 47282 52670 47294 52722
rect 47346 52719 47358 52722
rect 47618 52719 47630 52722
rect 47346 52673 47630 52719
rect 47346 52670 47358 52673
rect 47618 52670 47630 52673
rect 47682 52670 47694 52722
rect 10334 52658 10386 52670
rect 54014 52658 54066 52670
rect 54350 52722 54402 52734
rect 54350 52658 54402 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 8766 52386 8818 52398
rect 8766 52322 8818 52334
rect 15710 52386 15762 52398
rect 15710 52322 15762 52334
rect 16158 52386 16210 52398
rect 20414 52386 20466 52398
rect 55918 52386 55970 52398
rect 16482 52334 16494 52386
rect 16546 52334 16558 52386
rect 36082 52334 36094 52386
rect 36146 52334 36158 52386
rect 16158 52322 16210 52334
rect 20414 52322 20466 52334
rect 55918 52322 55970 52334
rect 56142 52386 56194 52398
rect 56142 52322 56194 52334
rect 56254 52386 56306 52398
rect 56254 52322 56306 52334
rect 4622 52274 4674 52286
rect 4622 52210 4674 52222
rect 7310 52274 7362 52286
rect 12350 52274 12402 52286
rect 18510 52274 18562 52286
rect 20190 52274 20242 52286
rect 21534 52274 21586 52286
rect 32398 52274 32450 52286
rect 35982 52274 36034 52286
rect 8194 52222 8206 52274
rect 8258 52222 8270 52274
rect 13682 52222 13694 52274
rect 13746 52222 13758 52274
rect 19394 52222 19406 52274
rect 19458 52222 19470 52274
rect 20738 52222 20750 52274
rect 20802 52222 20814 52274
rect 24546 52222 24558 52274
rect 24610 52222 24622 52274
rect 33618 52222 33630 52274
rect 33682 52222 33694 52274
rect 7310 52210 7362 52222
rect 12350 52210 12402 52222
rect 18510 52210 18562 52222
rect 20190 52210 20242 52222
rect 21534 52210 21586 52222
rect 32398 52210 32450 52222
rect 35982 52210 36034 52222
rect 39454 52274 39506 52286
rect 39454 52210 39506 52222
rect 43262 52274 43314 52286
rect 51774 52274 51826 52286
rect 46722 52222 46734 52274
rect 46786 52222 46798 52274
rect 47618 52222 47630 52274
rect 47682 52222 47694 52274
rect 51202 52222 51214 52274
rect 51266 52222 51278 52274
rect 43262 52210 43314 52222
rect 51774 52210 51826 52222
rect 8654 52162 8706 52174
rect 7970 52110 7982 52162
rect 8034 52110 8046 52162
rect 8654 52098 8706 52110
rect 10334 52162 10386 52174
rect 10334 52098 10386 52110
rect 10782 52162 10834 52174
rect 10782 52098 10834 52110
rect 12910 52162 12962 52174
rect 14478 52162 14530 52174
rect 13794 52110 13806 52162
rect 13858 52110 13870 52162
rect 12910 52098 12962 52110
rect 14478 52098 14530 52110
rect 14814 52162 14866 52174
rect 14814 52098 14866 52110
rect 15038 52162 15090 52174
rect 15038 52098 15090 52110
rect 15262 52162 15314 52174
rect 15262 52098 15314 52110
rect 15934 52162 15986 52174
rect 31502 52162 31554 52174
rect 38894 52162 38946 52174
rect 19170 52110 19182 52162
rect 19234 52110 19246 52162
rect 23090 52110 23102 52162
rect 23154 52110 23166 52162
rect 30930 52110 30942 52162
rect 30994 52110 31006 52162
rect 31826 52110 31838 52162
rect 31890 52110 31902 52162
rect 32722 52110 32734 52162
rect 32786 52110 32798 52162
rect 33282 52110 33294 52162
rect 33346 52110 33358 52162
rect 35634 52110 35646 52162
rect 35698 52110 35710 52162
rect 15934 52098 15986 52110
rect 31502 52098 31554 52110
rect 38894 52098 38946 52110
rect 43822 52162 43874 52174
rect 54126 52162 54178 52174
rect 46610 52110 46622 52162
rect 46674 52110 46686 52162
rect 50530 52110 50542 52162
rect 50594 52110 50606 52162
rect 50978 52110 50990 52162
rect 51042 52110 51054 52162
rect 43822 52098 43874 52110
rect 54126 52098 54178 52110
rect 8766 52050 8818 52062
rect 43150 52050 43202 52062
rect 9986 51998 9998 52050
rect 10050 51998 10062 52050
rect 11442 51998 11454 52050
rect 11506 51998 11518 52050
rect 24322 51998 24334 52050
rect 24386 51998 24398 52050
rect 30706 51998 30718 52050
rect 30770 51998 30782 52050
rect 33730 51998 33742 52050
rect 33794 51998 33806 52050
rect 8766 51986 8818 51998
rect 43150 51986 43202 51998
rect 44158 52050 44210 52062
rect 44158 51986 44210 51998
rect 47070 52050 47122 52062
rect 47070 51986 47122 51998
rect 47294 52050 47346 52062
rect 49746 51998 49758 52050
rect 49810 51998 49822 52050
rect 47294 51986 47346 51998
rect 11790 51938 11842 51950
rect 11790 51874 11842 51886
rect 12238 51938 12290 51950
rect 12238 51874 12290 51886
rect 12462 51938 12514 51950
rect 43374 51938 43426 51950
rect 22530 51886 22542 51938
rect 22594 51886 22606 51938
rect 12462 51874 12514 51886
rect 43374 51874 43426 51886
rect 46846 51938 46898 51950
rect 56254 51938 56306 51950
rect 54450 51886 54462 51938
rect 54514 51886 54526 51938
rect 46846 51874 46898 51886
rect 56254 51874 56306 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 3950 51602 4002 51614
rect 3950 51538 4002 51550
rect 12798 51602 12850 51614
rect 12798 51538 12850 51550
rect 13022 51602 13074 51614
rect 13022 51538 13074 51550
rect 13246 51602 13298 51614
rect 13246 51538 13298 51550
rect 15150 51602 15202 51614
rect 15150 51538 15202 51550
rect 32510 51602 32562 51614
rect 43262 51602 43314 51614
rect 36306 51550 36318 51602
rect 36370 51550 36382 51602
rect 32510 51538 32562 51550
rect 43262 51538 43314 51550
rect 47182 51602 47234 51614
rect 47182 51538 47234 51550
rect 48302 51602 48354 51614
rect 48302 51538 48354 51550
rect 48862 51602 48914 51614
rect 48862 51538 48914 51550
rect 51886 51602 51938 51614
rect 56702 51602 56754 51614
rect 52770 51550 52782 51602
rect 52834 51550 52846 51602
rect 55906 51550 55918 51602
rect 55970 51550 55982 51602
rect 51886 51538 51938 51550
rect 56702 51538 56754 51550
rect 3390 51490 3442 51502
rect 38670 51490 38722 51502
rect 5394 51438 5406 51490
rect 5458 51438 5470 51490
rect 37314 51438 37326 51490
rect 37378 51438 37390 51490
rect 3390 51426 3442 51438
rect 38670 51426 38722 51438
rect 41022 51490 41074 51502
rect 41022 51426 41074 51438
rect 41694 51490 41746 51502
rect 41694 51426 41746 51438
rect 48750 51490 48802 51502
rect 48750 51426 48802 51438
rect 53230 51490 53282 51502
rect 53230 51426 53282 51438
rect 55470 51490 55522 51502
rect 55470 51426 55522 51438
rect 3278 51378 3330 51390
rect 3278 51314 3330 51326
rect 3614 51378 3666 51390
rect 3614 51314 3666 51326
rect 4174 51378 4226 51390
rect 4174 51314 4226 51326
rect 4398 51378 4450 51390
rect 13358 51378 13410 51390
rect 5058 51326 5070 51378
rect 5122 51326 5134 51378
rect 5730 51326 5742 51378
rect 5794 51326 5806 51378
rect 4398 51314 4450 51326
rect 13358 51314 13410 51326
rect 14590 51378 14642 51390
rect 14590 51314 14642 51326
rect 15038 51378 15090 51390
rect 15038 51314 15090 51326
rect 15262 51378 15314 51390
rect 15262 51314 15314 51326
rect 28366 51378 28418 51390
rect 28366 51314 28418 51326
rect 28478 51378 28530 51390
rect 41582 51378 41634 51390
rect 47294 51378 47346 51390
rect 29138 51326 29150 51378
rect 29202 51326 29214 51378
rect 30146 51326 30158 51378
rect 30210 51326 30222 51378
rect 36194 51326 36206 51378
rect 36258 51326 36270 51378
rect 36754 51326 36766 51378
rect 36818 51326 36830 51378
rect 37986 51326 37998 51378
rect 38050 51326 38062 51378
rect 43698 51326 43710 51378
rect 43762 51326 43774 51378
rect 46946 51326 46958 51378
rect 47010 51326 47022 51378
rect 28478 51314 28530 51326
rect 41582 51314 41634 51326
rect 47294 51314 47346 51326
rect 47630 51378 47682 51390
rect 52446 51378 52498 51390
rect 55358 51378 55410 51390
rect 52098 51326 52110 51378
rect 52162 51326 52174 51378
rect 55122 51326 55134 51378
rect 55186 51326 55198 51378
rect 47630 51314 47682 51326
rect 52446 51314 52498 51326
rect 55358 51314 55410 51326
rect 56478 51378 56530 51390
rect 56478 51314 56530 51326
rect 56814 51378 56866 51390
rect 56814 51314 56866 51326
rect 57038 51378 57090 51390
rect 57038 51314 57090 51326
rect 4286 51266 4338 51278
rect 29038 51266 29090 51278
rect 42254 51266 42306 51278
rect 47854 51266 47906 51278
rect 5506 51214 5518 51266
rect 5570 51214 5582 51266
rect 29810 51214 29822 51266
rect 29874 51214 29886 51266
rect 37762 51214 37774 51266
rect 37826 51214 37838 51266
rect 44370 51214 44382 51266
rect 44434 51214 44446 51266
rect 46498 51214 46510 51266
rect 46562 51214 46574 51266
rect 4286 51202 4338 51214
rect 29038 51202 29090 51214
rect 42254 51202 42306 51214
rect 47854 51202 47906 51214
rect 48190 51266 48242 51278
rect 48190 51202 48242 51214
rect 40910 51154 40962 51166
rect 40910 51090 40962 51102
rect 41246 51154 41298 51166
rect 41246 51090 41298 51102
rect 41694 51154 41746 51166
rect 41694 51090 41746 51102
rect 51774 51154 51826 51166
rect 51774 51090 51826 51102
rect 53118 51154 53170 51166
rect 53118 51090 53170 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 5070 50818 5122 50830
rect 5070 50754 5122 50766
rect 5742 50818 5794 50830
rect 5742 50754 5794 50766
rect 14366 50818 14418 50830
rect 14366 50754 14418 50766
rect 33406 50818 33458 50830
rect 11678 50706 11730 50718
rect 28354 50710 28366 50762
rect 28418 50710 28430 50762
rect 33406 50754 33458 50766
rect 41806 50818 41858 50830
rect 41806 50754 41858 50766
rect 44942 50706 44994 50718
rect 4610 50654 4622 50706
rect 4674 50654 4686 50706
rect 9314 50654 9326 50706
rect 9378 50654 9390 50706
rect 35186 50654 35198 50706
rect 35250 50654 35262 50706
rect 36306 50654 36318 50706
rect 36370 50654 36382 50706
rect 38546 50654 38558 50706
rect 38610 50654 38622 50706
rect 40674 50654 40686 50706
rect 40738 50654 40750 50706
rect 56018 50654 56030 50706
rect 56082 50654 56094 50706
rect 58146 50654 58158 50706
rect 58210 50654 58222 50706
rect 11678 50642 11730 50654
rect 44942 50642 44994 50654
rect 4958 50594 5010 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 4958 50530 5010 50542
rect 5630 50594 5682 50606
rect 14030 50594 14082 50606
rect 29262 50594 29314 50606
rect 30158 50594 30210 50606
rect 9090 50542 9102 50594
rect 9154 50542 9166 50594
rect 9762 50542 9774 50594
rect 9826 50542 9838 50594
rect 25442 50542 25454 50594
rect 25506 50542 25518 50594
rect 29474 50542 29486 50594
rect 29538 50542 29550 50594
rect 5630 50530 5682 50542
rect 14030 50530 14082 50542
rect 29262 50530 29314 50542
rect 30158 50530 30210 50542
rect 30382 50594 30434 50606
rect 30382 50530 30434 50542
rect 30942 50594 30994 50606
rect 41918 50594 41970 50606
rect 32274 50542 32286 50594
rect 32338 50542 32350 50594
rect 32498 50542 32510 50594
rect 32562 50542 32574 50594
rect 33282 50542 33294 50594
rect 33346 50542 33358 50594
rect 35074 50542 35086 50594
rect 35138 50542 35150 50594
rect 41458 50542 41470 50594
rect 41522 50542 41534 50594
rect 30942 50530 30994 50542
rect 41918 50530 41970 50542
rect 42142 50594 42194 50606
rect 42142 50530 42194 50542
rect 42254 50594 42306 50606
rect 42254 50530 42306 50542
rect 42814 50594 42866 50606
rect 42814 50530 42866 50542
rect 44830 50594 44882 50606
rect 44830 50530 44882 50542
rect 45502 50594 45554 50606
rect 45502 50530 45554 50542
rect 45838 50594 45890 50606
rect 47182 50594 47234 50606
rect 46722 50542 46734 50594
rect 46786 50542 46798 50594
rect 47394 50542 47406 50594
rect 47458 50542 47470 50594
rect 55234 50542 55246 50594
rect 55298 50542 55310 50594
rect 45838 50530 45890 50542
rect 47182 50530 47234 50542
rect 5742 50482 5794 50494
rect 10782 50482 10834 50494
rect 2482 50430 2494 50482
rect 2546 50430 2558 50482
rect 8754 50430 8766 50482
rect 8818 50430 8830 50482
rect 5742 50418 5794 50430
rect 10782 50418 10834 50430
rect 11118 50482 11170 50494
rect 11118 50418 11170 50430
rect 19630 50482 19682 50494
rect 19630 50418 19682 50430
rect 25118 50482 25170 50494
rect 30606 50482 30658 50494
rect 26226 50430 26238 50482
rect 26290 50430 26302 50482
rect 25118 50418 25170 50430
rect 30606 50418 30658 50430
rect 30830 50482 30882 50494
rect 30830 50418 30882 50430
rect 47854 50482 47906 50494
rect 47854 50418 47906 50430
rect 13694 50370 13746 50382
rect 13694 50306 13746 50318
rect 14254 50370 14306 50382
rect 14254 50306 14306 50318
rect 19742 50370 19794 50382
rect 19742 50306 19794 50318
rect 45054 50370 45106 50382
rect 45054 50306 45106 50318
rect 46958 50370 47010 50382
rect 46958 50306 47010 50318
rect 47070 50370 47122 50382
rect 47070 50306 47122 50318
rect 54910 50370 54962 50382
rect 54910 50306 54962 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 4510 50034 4562 50046
rect 4510 49970 4562 49982
rect 9438 50034 9490 50046
rect 9438 49970 9490 49982
rect 12350 50034 12402 50046
rect 12350 49970 12402 49982
rect 28478 50034 28530 50046
rect 28478 49970 28530 49982
rect 28702 50034 28754 50046
rect 28702 49970 28754 49982
rect 29374 50034 29426 50046
rect 29374 49970 29426 49982
rect 29486 50034 29538 50046
rect 29486 49970 29538 49982
rect 30158 50034 30210 50046
rect 41022 50034 41074 50046
rect 35410 49982 35422 50034
rect 35474 49982 35486 50034
rect 30158 49970 30210 49982
rect 41022 49970 41074 49982
rect 41358 50034 41410 50046
rect 41358 49970 41410 49982
rect 51102 50034 51154 50046
rect 51102 49970 51154 49982
rect 4062 49922 4114 49934
rect 4062 49858 4114 49870
rect 9662 49922 9714 49934
rect 9662 49858 9714 49870
rect 10222 49922 10274 49934
rect 10222 49858 10274 49870
rect 19294 49922 19346 49934
rect 21534 49922 21586 49934
rect 20290 49870 20302 49922
rect 20354 49870 20366 49922
rect 19294 49858 19346 49870
rect 21534 49858 21586 49870
rect 28366 49922 28418 49934
rect 28366 49858 28418 49870
rect 29038 49922 29090 49934
rect 29038 49858 29090 49870
rect 29822 49922 29874 49934
rect 29822 49858 29874 49870
rect 29934 49922 29986 49934
rect 29934 49858 29986 49870
rect 34078 49922 34130 49934
rect 39342 49922 39394 49934
rect 37650 49870 37662 49922
rect 37714 49870 37726 49922
rect 34078 49858 34130 49870
rect 39342 49858 39394 49870
rect 41918 49922 41970 49934
rect 41918 49858 41970 49870
rect 47294 49922 47346 49934
rect 47294 49858 47346 49870
rect 50878 49922 50930 49934
rect 50878 49858 50930 49870
rect 51662 49922 51714 49934
rect 51662 49858 51714 49870
rect 51998 49922 52050 49934
rect 51998 49858 52050 49870
rect 52222 49922 52274 49934
rect 52222 49858 52274 49870
rect 3950 49810 4002 49822
rect 3378 49758 3390 49810
rect 3442 49758 3454 49810
rect 3950 49746 4002 49758
rect 4286 49810 4338 49822
rect 4286 49746 4338 49758
rect 4734 49810 4786 49822
rect 4734 49746 4786 49758
rect 4846 49810 4898 49822
rect 8878 49810 8930 49822
rect 8642 49758 8654 49810
rect 8706 49758 8718 49810
rect 4846 49746 4898 49758
rect 8878 49746 8930 49758
rect 9774 49810 9826 49822
rect 9774 49746 9826 49758
rect 9998 49810 10050 49822
rect 9998 49746 10050 49758
rect 10334 49810 10386 49822
rect 10334 49746 10386 49758
rect 12686 49810 12738 49822
rect 12686 49746 12738 49758
rect 13246 49810 13298 49822
rect 19182 49810 19234 49822
rect 14242 49758 14254 49810
rect 14306 49758 14318 49810
rect 13246 49746 13298 49758
rect 19182 49746 19234 49758
rect 19518 49810 19570 49822
rect 21422 49810 21474 49822
rect 29262 49810 29314 49822
rect 20178 49758 20190 49810
rect 20242 49758 20254 49810
rect 21186 49758 21198 49810
rect 21250 49758 21262 49810
rect 23762 49758 23774 49810
rect 23826 49758 23838 49810
rect 19518 49746 19570 49758
rect 21422 49746 21474 49758
rect 29262 49746 29314 49758
rect 31614 49810 31666 49822
rect 35086 49810 35138 49822
rect 41246 49810 41298 49822
rect 32050 49758 32062 49810
rect 32114 49758 32126 49810
rect 33394 49758 33406 49810
rect 33458 49758 33470 49810
rect 38658 49758 38670 49810
rect 38722 49758 38734 49810
rect 31614 49746 31666 49758
rect 35086 49746 35138 49758
rect 41246 49746 41298 49758
rect 41470 49810 41522 49822
rect 41470 49746 41522 49758
rect 50766 49810 50818 49822
rect 50766 49746 50818 49758
rect 52670 49810 52722 49822
rect 52670 49746 52722 49758
rect 5406 49698 5458 49710
rect 5406 49634 5458 49646
rect 7982 49698 8034 49710
rect 30494 49698 30546 49710
rect 14018 49646 14030 49698
rect 14082 49646 14094 49698
rect 20514 49646 20526 49698
rect 20578 49646 20590 49698
rect 23650 49646 23662 49698
rect 23714 49646 23726 49698
rect 7982 49634 8034 49646
rect 30494 49634 30546 49646
rect 31054 49698 31106 49710
rect 34862 49698 34914 49710
rect 42142 49698 42194 49710
rect 32386 49646 32398 49698
rect 32450 49646 32462 49698
rect 33170 49646 33182 49698
rect 33234 49646 33246 49698
rect 37202 49646 37214 49698
rect 37266 49646 37278 49698
rect 41794 49646 41806 49698
rect 41858 49646 41870 49698
rect 31054 49634 31106 49646
rect 34862 49634 34914 49646
rect 42142 49634 42194 49646
rect 49870 49698 49922 49710
rect 49870 49634 49922 49646
rect 50430 49698 50482 49710
rect 50430 49634 50482 49646
rect 52446 49698 52498 49710
rect 52446 49634 52498 49646
rect 21534 49586 21586 49598
rect 14690 49534 14702 49586
rect 14754 49534 14766 49586
rect 21534 49522 21586 49534
rect 23438 49586 23490 49598
rect 23438 49522 23490 49534
rect 47406 49586 47458 49598
rect 47406 49522 47458 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 32958 49250 33010 49262
rect 32958 49186 33010 49198
rect 33294 49250 33346 49262
rect 33294 49186 33346 49198
rect 53006 49250 53058 49262
rect 53006 49186 53058 49198
rect 10222 49138 10274 49150
rect 16270 49138 16322 49150
rect 20078 49138 20130 49150
rect 32734 49138 32786 49150
rect 8866 49086 8878 49138
rect 8930 49086 8942 49138
rect 15810 49086 15822 49138
rect 15874 49086 15886 49138
rect 17378 49086 17390 49138
rect 17442 49086 17454 49138
rect 19506 49086 19518 49138
rect 19570 49086 19582 49138
rect 23650 49086 23662 49138
rect 23714 49086 23726 49138
rect 25778 49086 25790 49138
rect 25842 49086 25854 49138
rect 10222 49074 10274 49086
rect 16270 49074 16322 49086
rect 20078 49074 20130 49086
rect 32734 49074 32786 49086
rect 33742 49138 33794 49150
rect 33742 49074 33794 49086
rect 42142 49138 42194 49150
rect 46722 49086 46734 49138
rect 46786 49086 46798 49138
rect 48850 49086 48862 49138
rect 48914 49086 48926 49138
rect 58146 49086 58158 49138
rect 58210 49086 58222 49138
rect 42142 49074 42194 49086
rect 9102 49026 9154 49038
rect 6066 48974 6078 49026
rect 6130 48974 6142 49026
rect 9102 48962 9154 48974
rect 9662 49026 9714 49038
rect 21982 49026 22034 49038
rect 15586 48974 15598 49026
rect 15650 48974 15662 49026
rect 16706 48974 16718 49026
rect 16770 48974 16782 49026
rect 9662 48962 9714 48974
rect 21982 48962 22034 48974
rect 22542 49026 22594 49038
rect 32174 49026 32226 49038
rect 22978 48974 22990 49026
rect 23042 48974 23054 49026
rect 31714 48974 31726 49026
rect 31778 48974 31790 49026
rect 22542 48962 22594 48974
rect 32174 48962 32226 48974
rect 32398 49026 32450 49038
rect 32398 48962 32450 48974
rect 41918 49026 41970 49038
rect 41918 48962 41970 48974
rect 42030 49026 42082 49038
rect 42030 48962 42082 48974
rect 42254 49026 42306 49038
rect 42254 48962 42306 48974
rect 42814 49026 42866 49038
rect 51102 49026 51154 49038
rect 49634 48974 49646 49026
rect 49698 48974 49710 49026
rect 50866 48974 50878 49026
rect 50930 48974 50942 49026
rect 42814 48962 42866 48974
rect 51102 48962 51154 48974
rect 51550 49026 51602 49038
rect 51550 48962 51602 48974
rect 52782 49026 52834 49038
rect 54910 49026 54962 49038
rect 53218 48974 53230 49026
rect 53282 48974 53294 49026
rect 54114 48974 54126 49026
rect 54178 48974 54190 49026
rect 54450 48974 54462 49026
rect 54514 48974 54526 49026
rect 55234 48974 55246 49026
rect 55298 48974 55310 49026
rect 52782 48962 52834 48974
rect 54910 48962 54962 48974
rect 9326 48914 9378 48926
rect 6738 48862 6750 48914
rect 6802 48862 6814 48914
rect 9326 48850 9378 48862
rect 9550 48914 9602 48926
rect 9550 48850 9602 48862
rect 11118 48914 11170 48926
rect 11118 48850 11170 48862
rect 19966 48914 20018 48926
rect 19966 48850 20018 48862
rect 20302 48914 20354 48926
rect 20302 48850 20354 48862
rect 20526 48914 20578 48926
rect 20526 48850 20578 48862
rect 21422 48914 21474 48926
rect 21422 48850 21474 48862
rect 43150 48914 43202 48926
rect 43150 48850 43202 48862
rect 54686 48914 54738 48926
rect 56018 48862 56030 48914
rect 56082 48862 56094 48914
rect 54686 48850 54738 48862
rect 11230 48802 11282 48814
rect 11230 48738 11282 48750
rect 11342 48802 11394 48814
rect 11342 48738 11394 48750
rect 21310 48802 21362 48814
rect 21310 48738 21362 48750
rect 21534 48802 21586 48814
rect 21534 48738 21586 48750
rect 42366 48802 42418 48814
rect 42366 48738 42418 48750
rect 43038 48802 43090 48814
rect 43038 48738 43090 48750
rect 50990 48802 51042 48814
rect 50990 48738 51042 48750
rect 52110 48802 52162 48814
rect 52110 48738 52162 48750
rect 53118 48802 53170 48814
rect 53118 48738 53170 48750
rect 53902 48802 53954 48814
rect 53902 48738 53954 48750
rect 54798 48802 54850 48814
rect 54798 48738 54850 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 8318 48466 8370 48478
rect 8318 48402 8370 48414
rect 8430 48466 8482 48478
rect 8430 48402 8482 48414
rect 8542 48466 8594 48478
rect 8542 48402 8594 48414
rect 8990 48466 9042 48478
rect 8990 48402 9042 48414
rect 19070 48466 19122 48478
rect 19070 48402 19122 48414
rect 20974 48466 21026 48478
rect 24446 48466 24498 48478
rect 22082 48414 22094 48466
rect 22146 48414 22158 48466
rect 20974 48402 21026 48414
rect 24446 48402 24498 48414
rect 27358 48466 27410 48478
rect 27358 48402 27410 48414
rect 32510 48466 32562 48478
rect 32510 48402 32562 48414
rect 41694 48466 41746 48478
rect 41694 48402 41746 48414
rect 42478 48466 42530 48478
rect 42478 48402 42530 48414
rect 55918 48466 55970 48478
rect 55918 48402 55970 48414
rect 5854 48354 5906 48366
rect 4834 48302 4846 48354
rect 4898 48302 4910 48354
rect 5854 48290 5906 48302
rect 6078 48354 6130 48366
rect 6078 48290 6130 48302
rect 8094 48354 8146 48366
rect 8094 48290 8146 48302
rect 8878 48354 8930 48366
rect 13918 48354 13970 48366
rect 20414 48354 20466 48366
rect 42366 48354 42418 48366
rect 10546 48302 10558 48354
rect 10610 48302 10622 48354
rect 14578 48302 14590 48354
rect 14642 48302 14654 48354
rect 15250 48302 15262 48354
rect 15314 48302 15326 48354
rect 23538 48302 23550 48354
rect 23602 48302 23614 48354
rect 37202 48302 37214 48354
rect 37266 48302 37278 48354
rect 8878 48290 8930 48302
rect 13918 48290 13970 48302
rect 20414 48290 20466 48302
rect 42366 48290 42418 48302
rect 43374 48354 43426 48366
rect 55470 48354 55522 48366
rect 52994 48302 53006 48354
rect 53058 48302 53070 48354
rect 43374 48290 43426 48302
rect 55470 48290 55522 48302
rect 55694 48354 55746 48366
rect 55694 48290 55746 48302
rect 6190 48242 6242 48254
rect 14030 48242 14082 48254
rect 19518 48242 19570 48254
rect 27246 48242 27298 48254
rect 4610 48190 4622 48242
rect 4674 48190 4686 48242
rect 5506 48190 5518 48242
rect 5570 48190 5582 48242
rect 11106 48190 11118 48242
rect 11170 48190 11182 48242
rect 11778 48190 11790 48242
rect 11842 48190 11854 48242
rect 14914 48190 14926 48242
rect 14978 48190 14990 48242
rect 15474 48190 15486 48242
rect 15538 48190 15550 48242
rect 19954 48190 19966 48242
rect 20018 48190 20030 48242
rect 22418 48190 22430 48242
rect 22482 48190 22494 48242
rect 6190 48178 6242 48190
rect 14030 48178 14082 48190
rect 19518 48178 19570 48190
rect 27246 48178 27298 48190
rect 27470 48242 27522 48254
rect 27470 48178 27522 48190
rect 27918 48242 27970 48254
rect 43262 48242 43314 48254
rect 35970 48190 35982 48242
rect 36034 48190 36046 48242
rect 37090 48190 37102 48242
rect 37154 48190 37166 48242
rect 27918 48178 27970 48190
rect 43262 48178 43314 48190
rect 43486 48242 43538 48254
rect 43486 48178 43538 48190
rect 43934 48242 43986 48254
rect 43934 48178 43986 48190
rect 49198 48242 49250 48254
rect 49198 48178 49250 48190
rect 50094 48242 50146 48254
rect 54238 48242 54290 48254
rect 53666 48190 53678 48242
rect 53730 48190 53742 48242
rect 50094 48178 50146 48190
rect 54238 48178 54290 48190
rect 54910 48242 54962 48254
rect 54910 48178 54962 48190
rect 56142 48242 56194 48254
rect 56142 48178 56194 48190
rect 12462 48130 12514 48142
rect 4946 48078 4958 48130
rect 5010 48078 5022 48130
rect 12462 48066 12514 48078
rect 13022 48130 13074 48142
rect 13022 48066 13074 48078
rect 14142 48130 14194 48142
rect 24670 48130 24722 48142
rect 41582 48130 41634 48142
rect 15362 48078 15374 48130
rect 15426 48078 15438 48130
rect 23874 48078 23886 48130
rect 23938 48078 23950 48130
rect 36642 48078 36654 48130
rect 36706 48078 36718 48130
rect 14142 48066 14194 48078
rect 24670 48066 24722 48078
rect 41582 48066 41634 48078
rect 48862 48130 48914 48142
rect 49634 48078 49646 48130
rect 49698 48078 49710 48130
rect 50866 48078 50878 48130
rect 50930 48078 50942 48130
rect 48862 48066 48914 48078
rect 24334 48018 24386 48030
rect 24334 47954 24386 47966
rect 42478 48018 42530 48030
rect 42478 47954 42530 47966
rect 50206 48018 50258 48030
rect 50206 47954 50258 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 5630 47682 5682 47694
rect 12462 47682 12514 47694
rect 28366 47682 28418 47694
rect 11106 47630 11118 47682
rect 11170 47630 11182 47682
rect 22642 47630 22654 47682
rect 22706 47630 22718 47682
rect 35410 47630 35422 47682
rect 35474 47630 35486 47682
rect 5630 47618 5682 47630
rect 12462 47618 12514 47630
rect 28366 47618 28418 47630
rect 5070 47570 5122 47582
rect 15486 47570 15538 47582
rect 25902 47570 25954 47582
rect 37998 47570 38050 47582
rect 4610 47518 4622 47570
rect 4674 47518 4686 47570
rect 11218 47518 11230 47570
rect 11282 47518 11294 47570
rect 17490 47518 17502 47570
rect 17554 47518 17566 47570
rect 23090 47518 23102 47570
rect 23154 47518 23166 47570
rect 29698 47518 29710 47570
rect 29762 47518 29774 47570
rect 34626 47518 34638 47570
rect 34690 47518 34702 47570
rect 37426 47518 37438 47570
rect 37490 47518 37502 47570
rect 5070 47506 5122 47518
rect 15486 47506 15538 47518
rect 25902 47506 25954 47518
rect 37998 47506 38050 47518
rect 44270 47570 44322 47582
rect 56254 47570 56306 47582
rect 47730 47518 47742 47570
rect 47794 47518 47806 47570
rect 44270 47506 44322 47518
rect 56254 47506 56306 47518
rect 12574 47458 12626 47470
rect 1810 47406 1822 47458
rect 1874 47406 1886 47458
rect 11106 47406 11118 47458
rect 11170 47406 11182 47458
rect 12226 47406 12238 47458
rect 12290 47406 12302 47458
rect 12574 47394 12626 47406
rect 15934 47458 15986 47470
rect 24558 47458 24610 47470
rect 17826 47406 17838 47458
rect 17890 47406 17902 47458
rect 22866 47406 22878 47458
rect 22930 47406 22942 47458
rect 23650 47406 23662 47458
rect 23714 47406 23726 47458
rect 15934 47394 15986 47406
rect 24558 47394 24610 47406
rect 24894 47458 24946 47470
rect 27918 47458 27970 47470
rect 27346 47406 27358 47458
rect 27410 47406 27422 47458
rect 34738 47406 34750 47458
rect 34802 47406 34814 47458
rect 37650 47406 37662 47458
rect 37714 47406 37726 47458
rect 38434 47406 38446 47458
rect 38498 47406 38510 47458
rect 38994 47406 39006 47458
rect 39058 47406 39070 47458
rect 41682 47406 41694 47458
rect 41746 47406 41758 47458
rect 42466 47406 42478 47458
rect 42530 47406 42542 47458
rect 44818 47406 44830 47458
rect 44882 47406 44894 47458
rect 52658 47406 52670 47458
rect 52722 47406 52734 47458
rect 24894 47394 24946 47406
rect 27918 47394 27970 47406
rect 5742 47346 5794 47358
rect 2482 47294 2494 47346
rect 2546 47294 2558 47346
rect 5742 47282 5794 47294
rect 5966 47346 6018 47358
rect 15374 47346 15426 47358
rect 13794 47294 13806 47346
rect 13858 47294 13870 47346
rect 15026 47294 15038 47346
rect 15090 47294 15102 47346
rect 5966 47282 6018 47294
rect 15374 47282 15426 47294
rect 15710 47346 15762 47358
rect 15710 47282 15762 47294
rect 18286 47346 18338 47358
rect 24782 47346 24834 47358
rect 28254 47346 28306 47358
rect 23986 47294 23998 47346
rect 24050 47294 24062 47346
rect 26114 47294 26126 47346
rect 26178 47294 26190 47346
rect 18286 47282 18338 47294
rect 24782 47282 24834 47294
rect 28254 47282 28306 47294
rect 29374 47346 29426 47358
rect 39106 47294 39118 47346
rect 39170 47294 39182 47346
rect 42578 47294 42590 47346
rect 42642 47294 42654 47346
rect 45602 47294 45614 47346
rect 45666 47294 45678 47346
rect 53442 47294 53454 47346
rect 53506 47294 53518 47346
rect 29374 47282 29426 47294
rect 12686 47234 12738 47246
rect 12686 47170 12738 47182
rect 14142 47234 14194 47246
rect 14142 47170 14194 47182
rect 14702 47234 14754 47246
rect 14702 47170 14754 47182
rect 24334 47234 24386 47246
rect 24334 47170 24386 47182
rect 25454 47234 25506 47246
rect 25454 47170 25506 47182
rect 28366 47234 28418 47246
rect 28366 47170 28418 47182
rect 29598 47234 29650 47246
rect 48526 47234 48578 47246
rect 38546 47182 38558 47234
rect 38610 47182 38622 47234
rect 41122 47182 41134 47234
rect 41186 47182 41198 47234
rect 29598 47170 29650 47182
rect 48526 47170 48578 47182
rect 49758 47234 49810 47246
rect 55682 47182 55694 47234
rect 55746 47182 55758 47234
rect 49758 47170 49810 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 2606 46898 2658 46910
rect 2606 46834 2658 46846
rect 12574 46898 12626 46910
rect 12574 46834 12626 46846
rect 13358 46898 13410 46910
rect 36094 46898 36146 46910
rect 13682 46846 13694 46898
rect 13746 46846 13758 46898
rect 24546 46846 24558 46898
rect 24610 46846 24622 46898
rect 27234 46846 27246 46898
rect 27298 46846 27310 46898
rect 35298 46846 35310 46898
rect 35362 46846 35374 46898
rect 13358 46834 13410 46846
rect 36094 46834 36146 46846
rect 36430 46898 36482 46910
rect 36430 46834 36482 46846
rect 45950 46898 46002 46910
rect 45950 46834 46002 46846
rect 53566 46898 53618 46910
rect 53566 46834 53618 46846
rect 2494 46786 2546 46798
rect 8878 46786 8930 46798
rect 5282 46734 5294 46786
rect 5346 46734 5358 46786
rect 2494 46722 2546 46734
rect 8878 46722 8930 46734
rect 12798 46786 12850 46798
rect 12798 46722 12850 46734
rect 12910 46786 12962 46798
rect 28590 46786 28642 46798
rect 23650 46734 23662 46786
rect 23714 46734 23726 46786
rect 12910 46722 12962 46734
rect 28590 46722 28642 46734
rect 28702 46786 28754 46798
rect 31950 46786 32002 46798
rect 29810 46734 29822 46786
rect 29874 46734 29886 46786
rect 31042 46734 31054 46786
rect 31106 46734 31118 46786
rect 28702 46722 28754 46734
rect 31950 46722 32002 46734
rect 34750 46786 34802 46798
rect 34750 46722 34802 46734
rect 35870 46786 35922 46798
rect 41022 46786 41074 46798
rect 37426 46734 37438 46786
rect 37490 46734 37502 46786
rect 39890 46734 39902 46786
rect 39954 46734 39966 46786
rect 35870 46722 35922 46734
rect 41022 46722 41074 46734
rect 41246 46786 41298 46798
rect 41246 46722 41298 46734
rect 46174 46786 46226 46798
rect 46174 46722 46226 46734
rect 48750 46786 48802 46798
rect 48750 46722 48802 46734
rect 8766 46674 8818 46686
rect 4050 46622 4062 46674
rect 4114 46622 4126 46674
rect 8766 46610 8818 46622
rect 9102 46674 9154 46686
rect 14030 46674 14082 46686
rect 28926 46674 28978 46686
rect 12338 46622 12350 46674
rect 12402 46622 12414 46674
rect 14690 46622 14702 46674
rect 14754 46622 14766 46674
rect 17826 46622 17838 46674
rect 17890 46622 17902 46674
rect 19394 46622 19406 46674
rect 19458 46622 19470 46674
rect 23538 46622 23550 46674
rect 23602 46622 23614 46674
rect 24434 46622 24446 46674
rect 24498 46622 24510 46674
rect 26002 46622 26014 46674
rect 26066 46622 26078 46674
rect 27458 46622 27470 46674
rect 27522 46622 27534 46674
rect 9102 46610 9154 46622
rect 14030 46610 14082 46622
rect 28926 46610 28978 46622
rect 34974 46674 35026 46686
rect 34974 46610 35026 46622
rect 35758 46674 35810 46686
rect 44494 46674 44546 46686
rect 45390 46674 45442 46686
rect 36642 46622 36654 46674
rect 36706 46622 36718 46674
rect 38882 46622 38894 46674
rect 38946 46622 38958 46674
rect 44818 46622 44830 46674
rect 44882 46622 44894 46674
rect 35758 46610 35810 46622
rect 44494 46610 44546 46622
rect 45390 46610 45442 46622
rect 45726 46674 45778 46686
rect 49310 46674 49362 46686
rect 50542 46674 50594 46686
rect 53678 46674 53730 46686
rect 48066 46622 48078 46674
rect 48130 46622 48142 46674
rect 49746 46622 49758 46674
rect 49810 46622 49822 46674
rect 53330 46622 53342 46674
rect 53394 46622 53406 46674
rect 45726 46610 45778 46622
rect 49310 46610 49362 46622
rect 50542 46610 50594 46622
rect 53678 46610 53730 46622
rect 54126 46674 54178 46686
rect 55010 46622 55022 46674
rect 55074 46622 55086 46674
rect 54126 46610 54178 46622
rect 2718 46562 2770 46574
rect 2718 46498 2770 46510
rect 3390 46562 3442 46574
rect 3390 46498 3442 46510
rect 5406 46562 5458 46574
rect 15374 46562 15426 46574
rect 26798 46562 26850 46574
rect 10098 46510 10110 46562
rect 10162 46510 10174 46562
rect 14914 46510 14926 46562
rect 14978 46510 14990 46562
rect 17714 46510 17726 46562
rect 17778 46510 17790 46562
rect 26226 46510 26238 46562
rect 26290 46510 26302 46562
rect 5406 46498 5458 46510
rect 15374 46498 15426 46510
rect 26798 46498 26850 46510
rect 29374 46562 29426 46574
rect 29374 46498 29426 46510
rect 31390 46562 31442 46574
rect 31390 46498 31442 46510
rect 31726 46562 31778 46574
rect 31726 46498 31778 46510
rect 32510 46562 32562 46574
rect 41694 46562 41746 46574
rect 37090 46510 37102 46562
rect 37154 46510 37166 46562
rect 32510 46498 32562 46510
rect 41694 46498 41746 46510
rect 45838 46562 45890 46574
rect 45838 46498 45890 46510
rect 47630 46562 47682 46574
rect 47630 46498 47682 46510
rect 50206 46562 50258 46574
rect 50206 46498 50258 46510
rect 51102 46562 51154 46574
rect 51102 46498 51154 46510
rect 53006 46562 53058 46574
rect 54786 46510 54798 46562
rect 54850 46510 54862 46562
rect 53006 46498 53058 46510
rect 32062 46450 32114 46462
rect 19730 46398 19742 46450
rect 19794 46398 19806 46450
rect 32062 46386 32114 46398
rect 36318 46450 36370 46462
rect 36318 46386 36370 46398
rect 40910 46450 40962 46462
rect 40910 46386 40962 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 29262 46114 29314 46126
rect 9650 46062 9662 46114
rect 9714 46062 9726 46114
rect 27570 46062 27582 46114
rect 27634 46062 27646 46114
rect 29262 46050 29314 46062
rect 2942 46002 2994 46014
rect 2942 45938 2994 45950
rect 9102 46002 9154 46014
rect 20190 46002 20242 46014
rect 42142 46002 42194 46014
rect 9986 45950 9998 46002
rect 10050 45950 10062 46002
rect 12114 45950 12126 46002
rect 12178 45950 12190 46002
rect 17714 45950 17726 46002
rect 17778 45950 17790 46002
rect 30034 45950 30046 46002
rect 30098 45950 30110 46002
rect 31042 45950 31054 46002
rect 31106 45950 31118 46002
rect 39554 45950 39566 46002
rect 39618 45950 39630 46002
rect 41682 45950 41694 46002
rect 41746 45950 41758 46002
rect 50866 45950 50878 46002
rect 50930 45950 50942 46002
rect 55234 45950 55246 46002
rect 55298 45950 55310 46002
rect 9102 45938 9154 45950
rect 20190 45938 20242 45950
rect 42142 45938 42194 45950
rect 8094 45890 8146 45902
rect 8094 45826 8146 45838
rect 9326 45890 9378 45902
rect 15822 45890 15874 45902
rect 27246 45890 27298 45902
rect 37550 45890 37602 45902
rect 45054 45890 45106 45902
rect 12786 45838 12798 45890
rect 12850 45838 12862 45890
rect 15026 45838 15038 45890
rect 15090 45838 15102 45890
rect 17042 45838 17054 45890
rect 17106 45838 17118 45890
rect 17826 45838 17838 45890
rect 17890 45838 17902 45890
rect 27906 45838 27918 45890
rect 27970 45838 27982 45890
rect 29026 45838 29038 45890
rect 29090 45838 29102 45890
rect 30146 45838 30158 45890
rect 30210 45838 30222 45890
rect 33954 45838 33966 45890
rect 34018 45838 34030 45890
rect 37986 45838 37998 45890
rect 38050 45838 38062 45890
rect 38882 45838 38894 45890
rect 38946 45838 38958 45890
rect 9326 45826 9378 45838
rect 15822 45826 15874 45838
rect 27246 45826 27298 45838
rect 37550 45826 37602 45838
rect 45054 45826 45106 45838
rect 45278 45890 45330 45902
rect 45278 45826 45330 45838
rect 45502 45890 45554 45902
rect 45502 45826 45554 45838
rect 48414 45890 48466 45902
rect 54910 45890 54962 45902
rect 49298 45838 49310 45890
rect 49362 45838 49374 45890
rect 58034 45838 58046 45890
rect 58098 45838 58110 45890
rect 48414 45826 48466 45838
rect 54910 45826 54962 45838
rect 15486 45778 15538 45790
rect 49534 45778 49586 45790
rect 14802 45726 14814 45778
rect 14866 45726 14878 45778
rect 18386 45726 18398 45778
rect 18450 45726 18462 45778
rect 33170 45726 33182 45778
rect 33234 45726 33246 45778
rect 15486 45714 15538 45726
rect 49534 45714 49586 45726
rect 49982 45778 50034 45790
rect 49982 45714 50034 45726
rect 51214 45778 51266 45790
rect 57362 45726 57374 45778
rect 57426 45726 57438 45778
rect 51214 45714 51266 45726
rect 7982 45666 8034 45678
rect 7982 45602 8034 45614
rect 8206 45666 8258 45678
rect 8206 45602 8258 45614
rect 8430 45666 8482 45678
rect 8430 45602 8482 45614
rect 13582 45666 13634 45678
rect 13582 45602 13634 45614
rect 15598 45666 15650 45678
rect 15598 45602 15650 45614
rect 20750 45666 20802 45678
rect 20750 45602 20802 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 23102 45666 23154 45678
rect 23102 45602 23154 45614
rect 28590 45666 28642 45678
rect 28590 45602 28642 45614
rect 34414 45666 34466 45678
rect 34414 45602 34466 45614
rect 45390 45666 45442 45678
rect 45390 45602 45442 45614
rect 45950 45666 46002 45678
rect 50654 45666 50706 45678
rect 48066 45614 48078 45666
rect 48130 45614 48142 45666
rect 45950 45602 46002 45614
rect 50654 45602 50706 45614
rect 50990 45666 51042 45678
rect 50990 45602 51042 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 3054 45330 3106 45342
rect 3054 45266 3106 45278
rect 9662 45330 9714 45342
rect 9662 45266 9714 45278
rect 9774 45330 9826 45342
rect 9774 45266 9826 45278
rect 22318 45330 22370 45342
rect 36654 45330 36706 45342
rect 23650 45278 23662 45330
rect 23714 45278 23726 45330
rect 24098 45278 24110 45330
rect 24162 45278 24174 45330
rect 28690 45278 28702 45330
rect 28754 45278 28766 45330
rect 22318 45266 22370 45278
rect 36654 45266 36706 45278
rect 38446 45330 38498 45342
rect 38446 45266 38498 45278
rect 48302 45330 48354 45342
rect 48302 45266 48354 45278
rect 48750 45330 48802 45342
rect 48750 45266 48802 45278
rect 53342 45330 53394 45342
rect 53342 45266 53394 45278
rect 55918 45330 55970 45342
rect 55918 45266 55970 45278
rect 58158 45330 58210 45342
rect 58158 45266 58210 45278
rect 4958 45218 5010 45230
rect 4958 45154 5010 45166
rect 14590 45218 14642 45230
rect 21758 45218 21810 45230
rect 15586 45166 15598 45218
rect 15650 45166 15662 45218
rect 14590 45154 14642 45166
rect 21758 45154 21810 45166
rect 22206 45218 22258 45230
rect 22206 45154 22258 45166
rect 25230 45218 25282 45230
rect 55134 45218 55186 45230
rect 31490 45166 31502 45218
rect 31554 45166 31566 45218
rect 49074 45166 49086 45218
rect 49138 45166 49150 45218
rect 50754 45166 50766 45218
rect 50818 45166 50830 45218
rect 25230 45154 25282 45166
rect 55134 45154 55186 45166
rect 57150 45218 57202 45230
rect 57150 45154 57202 45166
rect 5070 45106 5122 45118
rect 9550 45106 9602 45118
rect 21646 45106 21698 45118
rect 6066 45054 6078 45106
rect 6130 45054 6142 45106
rect 10098 45054 10110 45106
rect 10162 45054 10174 45106
rect 14914 45054 14926 45106
rect 14978 45054 14990 45106
rect 15810 45054 15822 45106
rect 15874 45054 15886 45106
rect 5070 45042 5122 45054
rect 9550 45042 9602 45054
rect 21646 45042 21698 45054
rect 21982 45106 22034 45118
rect 21982 45042 22034 45054
rect 22430 45106 22482 45118
rect 22430 45042 22482 45054
rect 22878 45106 22930 45118
rect 22878 45042 22930 45054
rect 23326 45106 23378 45118
rect 23326 45042 23378 45054
rect 25342 45106 25394 45118
rect 43822 45106 43874 45118
rect 55470 45106 55522 45118
rect 25778 45054 25790 45106
rect 25842 45054 25854 45106
rect 28466 45054 28478 45106
rect 28530 45054 28542 45106
rect 31714 45054 31726 45106
rect 31778 45054 31790 45106
rect 32498 45054 32510 45106
rect 32562 45054 32574 45106
rect 36194 45054 36206 45106
rect 36258 45054 36270 45106
rect 49970 45054 49982 45106
rect 50034 45054 50046 45106
rect 25342 45042 25394 45054
rect 43822 45042 43874 45054
rect 55470 45042 55522 45054
rect 55694 45106 55746 45118
rect 55694 45042 55746 45054
rect 56030 45106 56082 45118
rect 56814 45106 56866 45118
rect 56578 45054 56590 45106
rect 56642 45054 56654 45106
rect 56030 45042 56082 45054
rect 56814 45042 56866 45054
rect 57038 45106 57090 45118
rect 57038 45042 57090 45054
rect 20974 44994 21026 45006
rect 6738 44942 6750 44994
rect 6802 44942 6814 44994
rect 8866 44942 8878 44994
rect 8930 44942 8942 44994
rect 15698 44942 15710 44994
rect 15762 44942 15774 44994
rect 20974 44930 21026 44942
rect 23102 44994 23154 45006
rect 23102 44930 23154 44942
rect 24670 44994 24722 45006
rect 24670 44930 24722 44942
rect 29150 44994 29202 45006
rect 31938 44942 31950 44994
rect 32002 44942 32014 44994
rect 33282 44942 33294 44994
rect 33346 44942 33358 44994
rect 35410 44942 35422 44994
rect 35474 44942 35486 44994
rect 52882 44942 52894 44994
rect 52946 44942 52958 44994
rect 57698 44942 57710 44994
rect 57762 44942 57774 44994
rect 29150 44930 29202 44942
rect 4958 44882 5010 44894
rect 4958 44818 5010 44830
rect 24446 44882 24498 44894
rect 24446 44818 24498 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 3502 44546 3554 44558
rect 31726 44546 31778 44558
rect 54574 44546 54626 44558
rect 9314 44494 9326 44546
rect 9378 44543 9390 44546
rect 9650 44543 9662 44546
rect 9378 44497 9662 44543
rect 9378 44494 9390 44497
rect 9650 44494 9662 44497
rect 9714 44494 9726 44546
rect 16258 44494 16270 44546
rect 16322 44494 16334 44546
rect 45378 44494 45390 44546
rect 45442 44494 45454 44546
rect 51202 44494 51214 44546
rect 51266 44494 51278 44546
rect 3502 44482 3554 44494
rect 31726 44482 31778 44494
rect 54574 44482 54626 44494
rect 55246 44546 55298 44558
rect 56130 44494 56142 44546
rect 56194 44494 56206 44546
rect 55246 44482 55298 44494
rect 5630 44434 5682 44446
rect 4050 44382 4062 44434
rect 4114 44382 4126 44434
rect 5630 44370 5682 44382
rect 5966 44434 6018 44446
rect 5966 44370 6018 44382
rect 7310 44434 7362 44446
rect 7310 44370 7362 44382
rect 8094 44434 8146 44446
rect 9550 44434 9602 44446
rect 24110 44434 24162 44446
rect 8978 44382 8990 44434
rect 9042 44382 9054 44434
rect 16818 44382 16830 44434
rect 16882 44382 16894 44434
rect 19618 44382 19630 44434
rect 19682 44382 19694 44434
rect 8094 44370 8146 44382
rect 9550 44370 9602 44382
rect 24110 44370 24162 44382
rect 31390 44434 31442 44446
rect 57598 44434 57650 44446
rect 32274 44382 32286 44434
rect 32338 44382 32350 44434
rect 43586 44382 43598 44434
rect 43650 44382 43662 44434
rect 45490 44382 45502 44434
rect 45554 44382 45566 44434
rect 51762 44382 51774 44434
rect 51826 44382 51838 44434
rect 54226 44382 54238 44434
rect 54290 44382 54302 44434
rect 31390 44370 31442 44382
rect 57598 44370 57650 44382
rect 58270 44434 58322 44446
rect 58270 44370 58322 44382
rect 6190 44322 6242 44334
rect 2482 44270 2494 44322
rect 2546 44270 2558 44322
rect 4498 44270 4510 44322
rect 4562 44270 4574 44322
rect 4946 44270 4958 44322
rect 5010 44270 5022 44322
rect 6190 44258 6242 44270
rect 7534 44322 7586 44334
rect 7534 44258 7586 44270
rect 7758 44322 7810 44334
rect 16158 44322 16210 44334
rect 23326 44322 23378 44334
rect 8754 44270 8766 44322
rect 8818 44270 8830 44322
rect 15474 44270 15486 44322
rect 15538 44270 15550 44322
rect 17266 44270 17278 44322
rect 17330 44270 17342 44322
rect 17826 44270 17838 44322
rect 17890 44270 17902 44322
rect 18498 44270 18510 44322
rect 18562 44270 18574 44322
rect 21746 44270 21758 44322
rect 21810 44270 21822 44322
rect 22082 44270 22094 44322
rect 22146 44270 22158 44322
rect 7758 44258 7810 44270
rect 16158 44258 16210 44270
rect 23326 44258 23378 44270
rect 24782 44322 24834 44334
rect 31166 44322 31218 44334
rect 33070 44322 33122 44334
rect 25778 44270 25790 44322
rect 25842 44270 25854 44322
rect 32386 44270 32398 44322
rect 32450 44270 32462 44322
rect 24782 44258 24834 44270
rect 31166 44258 31218 44270
rect 33070 44258 33122 44270
rect 33742 44322 33794 44334
rect 33742 44258 33794 44270
rect 34302 44322 34354 44334
rect 34302 44258 34354 44270
rect 34750 44322 34802 44334
rect 34750 44258 34802 44270
rect 35310 44322 35362 44334
rect 44270 44322 44322 44334
rect 46510 44322 46562 44334
rect 40786 44270 40798 44322
rect 40850 44270 40862 44322
rect 44706 44270 44718 44322
rect 44770 44270 44782 44322
rect 45602 44270 45614 44322
rect 45666 44270 45678 44322
rect 35310 44258 35362 44270
rect 44270 44258 44322 44270
rect 46510 44258 46562 44270
rect 46958 44322 47010 44334
rect 55470 44322 55522 44334
rect 51874 44270 51886 44322
rect 51938 44270 51950 44322
rect 46958 44258 47010 44270
rect 55470 44258 55522 44270
rect 56590 44322 56642 44334
rect 56590 44258 56642 44270
rect 2830 44210 2882 44222
rect 2830 44146 2882 44158
rect 3502 44210 3554 44222
rect 3502 44146 3554 44158
rect 3614 44210 3666 44222
rect 7198 44210 7250 44222
rect 22318 44210 22370 44222
rect 3938 44158 3950 44210
rect 4002 44158 4014 44210
rect 13458 44158 13470 44210
rect 13522 44158 13534 44210
rect 16930 44158 16942 44210
rect 16994 44158 17006 44210
rect 3614 44146 3666 44158
rect 7198 44146 7250 44158
rect 22318 44146 22370 44158
rect 22654 44210 22706 44222
rect 25566 44210 25618 44222
rect 24434 44158 24446 44210
rect 24498 44158 24510 44210
rect 22654 44146 22706 44158
rect 25566 44146 25618 44158
rect 34078 44210 34130 44222
rect 43934 44210 43986 44222
rect 41458 44158 41470 44210
rect 41522 44158 41534 44210
rect 34078 44146 34130 44158
rect 43934 44146 43986 44158
rect 44046 44210 44098 44222
rect 44046 44146 44098 44158
rect 46846 44210 46898 44222
rect 46846 44146 46898 44158
rect 56702 44210 56754 44222
rect 56702 44146 56754 44158
rect 56814 44210 56866 44222
rect 56814 44146 56866 44158
rect 2718 44098 2770 44110
rect 2718 44034 2770 44046
rect 13806 44098 13858 44110
rect 13806 44034 13858 44046
rect 22766 44098 22818 44110
rect 22766 44034 22818 44046
rect 22878 44098 22930 44110
rect 22878 44034 22930 44046
rect 23662 44098 23714 44110
rect 23662 44034 23714 44046
rect 33966 44098 34018 44110
rect 33966 44034 34018 44046
rect 34638 44098 34690 44110
rect 34638 44034 34690 44046
rect 34862 44098 34914 44110
rect 34862 44034 34914 44046
rect 35646 44098 35698 44110
rect 35646 44034 35698 44046
rect 37886 44098 37938 44110
rect 37886 44034 37938 44046
rect 46622 44098 46674 44110
rect 46622 44034 46674 44046
rect 54350 44098 54402 44110
rect 54898 44046 54910 44098
rect 54962 44046 54974 44098
rect 54350 44034 54402 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 4958 43762 5010 43774
rect 4958 43698 5010 43710
rect 23214 43762 23266 43774
rect 32386 43710 32398 43762
rect 32450 43710 32462 43762
rect 37650 43710 37662 43762
rect 37714 43710 37726 43762
rect 23214 43698 23266 43710
rect 5070 43650 5122 43662
rect 2482 43598 2494 43650
rect 2546 43598 2558 43650
rect 5070 43586 5122 43598
rect 5518 43650 5570 43662
rect 5518 43586 5570 43598
rect 15374 43650 15426 43662
rect 15374 43586 15426 43598
rect 15598 43650 15650 43662
rect 15598 43586 15650 43598
rect 16382 43650 16434 43662
rect 22206 43650 22258 43662
rect 17714 43598 17726 43650
rect 17778 43598 17790 43650
rect 18274 43598 18286 43650
rect 18338 43598 18350 43650
rect 16382 43586 16434 43598
rect 22206 43586 22258 43598
rect 22542 43650 22594 43662
rect 22542 43586 22594 43598
rect 22766 43650 22818 43662
rect 22766 43586 22818 43598
rect 29822 43650 29874 43662
rect 57374 43650 57426 43662
rect 36642 43598 36654 43650
rect 36706 43598 36718 43650
rect 38546 43598 38558 43650
rect 38610 43598 38622 43650
rect 46050 43598 46062 43650
rect 46114 43598 46126 43650
rect 29822 43586 29874 43598
rect 57374 43586 57426 43598
rect 57822 43650 57874 43662
rect 57822 43586 57874 43598
rect 15710 43538 15762 43550
rect 1810 43486 1822 43538
rect 1874 43486 1886 43538
rect 15710 43474 15762 43486
rect 17614 43538 17666 43550
rect 29710 43538 29762 43550
rect 19058 43486 19070 43538
rect 19122 43486 19134 43538
rect 17614 43474 17666 43486
rect 29710 43474 29762 43486
rect 29934 43538 29986 43550
rect 31838 43538 31890 43550
rect 30258 43486 30270 43538
rect 30322 43486 30334 43538
rect 29934 43474 29986 43486
rect 31838 43474 31890 43486
rect 32062 43538 32114 43550
rect 41022 43538 41074 43550
rect 52782 43538 52834 43550
rect 37090 43486 37102 43538
rect 37154 43486 37166 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 39666 43486 39678 43538
rect 39730 43486 39742 43538
rect 41458 43486 41470 43538
rect 41522 43486 41534 43538
rect 45378 43486 45390 43538
rect 45442 43486 45454 43538
rect 53218 43486 53230 43538
rect 53282 43486 53294 43538
rect 32062 43474 32114 43486
rect 41022 43474 41074 43486
rect 52782 43474 52834 43486
rect 17390 43426 17442 43438
rect 22318 43426 22370 43438
rect 40350 43426 40402 43438
rect 44942 43426 44994 43438
rect 4610 43374 4622 43426
rect 4674 43374 4686 43426
rect 16482 43374 16494 43426
rect 16546 43374 16558 43426
rect 19730 43374 19742 43426
rect 19794 43374 19806 43426
rect 21858 43374 21870 43426
rect 21922 43374 21934 43426
rect 38210 43374 38222 43426
rect 38274 43374 38286 43426
rect 42466 43374 42478 43426
rect 42530 43374 42542 43426
rect 48178 43374 48190 43426
rect 48242 43374 48254 43426
rect 54786 43374 54798 43426
rect 54850 43374 54862 43426
rect 57138 43374 57150 43426
rect 57202 43374 57214 43426
rect 17390 43362 17442 43374
rect 22318 43362 22370 43374
rect 40350 43362 40402 43374
rect 44942 43362 44994 43374
rect 16158 43314 16210 43326
rect 57586 43262 57598 43314
rect 57650 43311 57662 43314
rect 57810 43311 57822 43314
rect 57650 43265 57822 43311
rect 57650 43262 57662 43265
rect 57810 43262 57822 43265
rect 57874 43311 57886 43314
rect 58146 43311 58158 43314
rect 57874 43265 58158 43311
rect 57874 43262 57886 43265
rect 58146 43262 58158 43265
rect 58210 43262 58222 43314
rect 16158 43250 16210 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 20190 42978 20242 42990
rect 37102 42978 37154 42990
rect 10098 42926 10110 42978
rect 10162 42926 10174 42978
rect 33170 42926 33182 42978
rect 33234 42975 33246 42978
rect 34066 42975 34078 42978
rect 33234 42929 34078 42975
rect 33234 42926 33246 42929
rect 34066 42926 34078 42929
rect 34130 42926 34142 42978
rect 20190 42914 20242 42926
rect 37102 42914 37154 42926
rect 45614 42978 45666 42990
rect 45614 42914 45666 42926
rect 50094 42978 50146 42990
rect 50094 42914 50146 42926
rect 53566 42978 53618 42990
rect 53566 42914 53618 42926
rect 53678 42978 53730 42990
rect 53678 42914 53730 42926
rect 53902 42978 53954 42990
rect 53902 42914 53954 42926
rect 2942 42866 2994 42878
rect 13022 42866 13074 42878
rect 22094 42866 22146 42878
rect 33182 42866 33234 42878
rect 3714 42814 3726 42866
rect 3778 42814 3790 42866
rect 16818 42814 16830 42866
rect 16882 42814 16894 42866
rect 25330 42814 25342 42866
rect 25394 42814 25406 42866
rect 31042 42814 31054 42866
rect 31106 42814 31118 42866
rect 2942 42802 2994 42814
rect 13022 42802 13074 42814
rect 22094 42802 22146 42814
rect 33182 42802 33234 42814
rect 34078 42866 34130 42878
rect 34078 42802 34130 42814
rect 40126 42866 40178 42878
rect 40126 42802 40178 42814
rect 41582 42866 41634 42878
rect 46734 42866 46786 42878
rect 44146 42814 44158 42866
rect 44210 42814 44222 42866
rect 41582 42802 41634 42814
rect 46734 42802 46786 42814
rect 51662 42866 51714 42878
rect 51662 42802 51714 42814
rect 53118 42866 53170 42878
rect 57026 42814 57038 42866
rect 57090 42814 57102 42866
rect 53118 42802 53170 42814
rect 8430 42754 8482 42766
rect 15710 42754 15762 42766
rect 3602 42702 3614 42754
rect 3666 42702 3678 42754
rect 8754 42702 8766 42754
rect 8818 42702 8830 42754
rect 9650 42702 9662 42754
rect 9714 42702 9726 42754
rect 10098 42702 10110 42754
rect 10162 42702 10174 42754
rect 10546 42702 10558 42754
rect 10610 42702 10622 42754
rect 14018 42702 14030 42754
rect 14082 42702 14094 42754
rect 14466 42702 14478 42754
rect 14530 42702 14542 42754
rect 15362 42702 15374 42754
rect 15426 42702 15438 42754
rect 8430 42690 8482 42702
rect 15710 42690 15762 42702
rect 15934 42754 15986 42766
rect 27470 42754 27522 42766
rect 16482 42702 16494 42754
rect 16546 42702 16558 42754
rect 18162 42702 18174 42754
rect 18226 42702 18238 42754
rect 19394 42702 19406 42754
rect 19458 42702 19470 42754
rect 25218 42702 25230 42754
rect 25282 42702 25294 42754
rect 26002 42702 26014 42754
rect 26066 42702 26078 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 27122 42702 27134 42754
rect 27186 42702 27198 42754
rect 15934 42690 15986 42702
rect 27470 42690 27522 42702
rect 27694 42754 27746 42766
rect 27694 42690 27746 42702
rect 28366 42754 28418 42766
rect 39230 42754 39282 42766
rect 46622 42754 46674 42766
rect 56478 42754 56530 42766
rect 29138 42702 29150 42754
rect 29202 42702 29214 42754
rect 30034 42702 30046 42754
rect 30098 42702 30110 42754
rect 30930 42702 30942 42754
rect 30994 42702 31006 42754
rect 37538 42702 37550 42754
rect 37602 42702 37614 42754
rect 38098 42702 38110 42754
rect 38162 42702 38174 42754
rect 39442 42702 39454 42754
rect 39506 42702 39518 42754
rect 51538 42702 51550 42754
rect 51602 42702 51614 42754
rect 51762 42702 51774 42754
rect 51826 42702 51838 42754
rect 55906 42702 55918 42754
rect 55970 42702 55982 42754
rect 28366 42690 28418 42702
rect 39230 42690 39282 42702
rect 46622 42690 46674 42702
rect 56478 42690 56530 42702
rect 9102 42642 9154 42654
rect 20302 42642 20354 42654
rect 13906 42590 13918 42642
rect 13970 42590 13982 42642
rect 16818 42590 16830 42642
rect 16882 42590 16894 42642
rect 9102 42578 9154 42590
rect 20302 42578 20354 42590
rect 20750 42642 20802 42654
rect 31278 42642 31330 42654
rect 25106 42590 25118 42642
rect 25170 42590 25182 42642
rect 30482 42590 30494 42642
rect 30546 42590 30558 42642
rect 20750 42578 20802 42590
rect 31278 42578 31330 42590
rect 37214 42642 37266 42654
rect 41694 42642 41746 42654
rect 38546 42590 38558 42642
rect 38610 42590 38622 42642
rect 37214 42578 37266 42590
rect 41694 42578 41746 42590
rect 42030 42642 42082 42654
rect 45614 42642 45666 42654
rect 42242 42590 42254 42642
rect 42306 42590 42318 42642
rect 43922 42590 43934 42642
rect 43986 42590 43998 42642
rect 42030 42578 42082 42590
rect 45614 42578 45666 42590
rect 45726 42642 45778 42654
rect 45726 42578 45778 42590
rect 50206 42642 50258 42654
rect 50206 42578 50258 42590
rect 54014 42642 54066 42654
rect 54014 42578 54066 42590
rect 55470 42642 55522 42654
rect 55470 42578 55522 42590
rect 56926 42642 56978 42654
rect 56926 42578 56978 42590
rect 8990 42530 9042 42542
rect 20526 42530 20578 42542
rect 14354 42478 14366 42530
rect 14418 42478 14430 42530
rect 8990 42466 9042 42478
rect 20526 42466 20578 42478
rect 21422 42530 21474 42542
rect 21422 42466 21474 42478
rect 28478 42530 28530 42542
rect 28478 42466 28530 42478
rect 28702 42530 28754 42542
rect 33630 42530 33682 42542
rect 29250 42478 29262 42530
rect 29314 42478 29326 42530
rect 29474 42478 29486 42530
rect 29538 42478 29550 42530
rect 28702 42466 28754 42478
rect 33630 42466 33682 42478
rect 36430 42530 36482 42542
rect 36430 42466 36482 42478
rect 37102 42530 37154 42542
rect 41022 42530 41074 42542
rect 37650 42478 37662 42530
rect 37714 42478 37726 42530
rect 37102 42466 37154 42478
rect 41022 42466 41074 42478
rect 41470 42530 41522 42542
rect 41470 42466 41522 42478
rect 45166 42530 45218 42542
rect 45166 42466 45218 42478
rect 46398 42530 46450 42542
rect 46398 42466 46450 42478
rect 46846 42530 46898 42542
rect 46846 42466 46898 42478
rect 49646 42530 49698 42542
rect 49646 42466 49698 42478
rect 50094 42530 50146 42542
rect 50094 42466 50146 42478
rect 51998 42530 52050 42542
rect 51998 42466 52050 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 14478 42194 14530 42206
rect 28030 42194 28082 42206
rect 20962 42142 20974 42194
rect 21026 42142 21038 42194
rect 14478 42130 14530 42142
rect 28030 42130 28082 42142
rect 28478 42194 28530 42206
rect 28478 42130 28530 42142
rect 58158 42194 58210 42206
rect 58158 42130 58210 42142
rect 8766 42082 8818 42094
rect 8766 42018 8818 42030
rect 9662 42082 9714 42094
rect 23886 42082 23938 42094
rect 11554 42030 11566 42082
rect 11618 42030 11630 42082
rect 15586 42030 15598 42082
rect 15650 42030 15662 42082
rect 18386 42030 18398 42082
rect 18450 42030 18462 42082
rect 20514 42030 20526 42082
rect 20578 42030 20590 42082
rect 9662 42018 9714 42030
rect 23886 42018 23938 42030
rect 24110 42082 24162 42094
rect 24110 42018 24162 42030
rect 24446 42082 24498 42094
rect 24446 42018 24498 42030
rect 24558 42082 24610 42094
rect 34078 42082 34130 42094
rect 27234 42030 27246 42082
rect 27298 42030 27310 42082
rect 24558 42018 24610 42030
rect 34078 42018 34130 42030
rect 35534 42082 35586 42094
rect 35534 42018 35586 42030
rect 43486 42082 43538 42094
rect 57038 42082 57090 42094
rect 53778 42030 53790 42082
rect 53842 42030 53854 42082
rect 43486 42018 43538 42030
rect 57038 42018 57090 42030
rect 57598 42082 57650 42094
rect 57598 42018 57650 42030
rect 8878 41970 8930 41982
rect 5394 41918 5406 41970
rect 5458 41918 5470 41970
rect 6066 41918 6078 41970
rect 6130 41918 6142 41970
rect 8878 41906 8930 41918
rect 9550 41970 9602 41982
rect 9550 41906 9602 41918
rect 9886 41970 9938 41982
rect 9886 41906 9938 41918
rect 10222 41970 10274 41982
rect 14142 41970 14194 41982
rect 12786 41918 12798 41970
rect 12850 41918 12862 41970
rect 10222 41906 10274 41918
rect 14142 41906 14194 41918
rect 14478 41970 14530 41982
rect 14478 41906 14530 41918
rect 14814 41970 14866 41982
rect 14814 41906 14866 41918
rect 15262 41970 15314 41982
rect 19854 41970 19906 41982
rect 23550 41970 23602 41982
rect 15474 41918 15486 41970
rect 15538 41918 15550 41970
rect 15922 41918 15934 41970
rect 15986 41918 15998 41970
rect 16706 41918 16718 41970
rect 16770 41918 16782 41970
rect 18274 41918 18286 41970
rect 18338 41918 18350 41970
rect 20626 41918 20638 41970
rect 20690 41918 20702 41970
rect 21410 41918 21422 41970
rect 21474 41918 21486 41970
rect 15262 41906 15314 41918
rect 19854 41906 19906 41918
rect 23550 41906 23602 41918
rect 24782 41970 24834 41982
rect 26910 41970 26962 41982
rect 25106 41918 25118 41970
rect 25170 41918 25182 41970
rect 25890 41918 25902 41970
rect 25954 41918 25966 41970
rect 24782 41906 24834 41918
rect 26910 41906 26962 41918
rect 27918 41970 27970 41982
rect 28590 41970 28642 41982
rect 28130 41918 28142 41970
rect 28194 41918 28206 41970
rect 27918 41906 27970 41918
rect 28590 41906 28642 41918
rect 28702 41970 28754 41982
rect 29486 41970 29538 41982
rect 30382 41970 30434 41982
rect 40350 41970 40402 41982
rect 29026 41918 29038 41970
rect 29090 41918 29102 41970
rect 29698 41918 29710 41970
rect 29762 41918 29774 41970
rect 33730 41918 33742 41970
rect 33794 41918 33806 41970
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 36866 41918 36878 41970
rect 36930 41918 36942 41970
rect 38770 41918 38782 41970
rect 38834 41918 38846 41970
rect 28702 41906 28754 41918
rect 29486 41906 29538 41918
rect 30382 41906 30434 41918
rect 40350 41906 40402 41918
rect 41134 41970 41186 41982
rect 41134 41906 41186 41918
rect 41358 41970 41410 41982
rect 41358 41906 41410 41918
rect 41806 41970 41858 41982
rect 52446 41970 52498 41982
rect 56702 41970 56754 41982
rect 43810 41918 43822 41970
rect 43874 41918 43886 41970
rect 49186 41918 49198 41970
rect 49250 41918 49262 41970
rect 53106 41918 53118 41970
rect 53170 41918 53182 41970
rect 41806 41906 41858 41918
rect 52446 41906 52498 41918
rect 56702 41906 56754 41918
rect 57374 41970 57426 41982
rect 57374 41906 57426 41918
rect 3278 41858 3330 41870
rect 21198 41858 21250 41870
rect 32510 41858 32562 41870
rect 39454 41858 39506 41870
rect 8194 41806 8206 41858
rect 8258 41806 8270 41858
rect 10994 41806 11006 41858
rect 11058 41806 11070 41858
rect 25778 41806 25790 41858
rect 25842 41806 25854 41858
rect 34402 41806 34414 41858
rect 34466 41806 34478 41858
rect 37202 41806 37214 41858
rect 37266 41806 37278 41858
rect 38098 41806 38110 41858
rect 38162 41806 38174 41858
rect 38882 41806 38894 41858
rect 38946 41806 38958 41858
rect 3278 41794 3330 41806
rect 21198 41794 21250 41806
rect 32510 41794 32562 41806
rect 39454 41794 39506 41806
rect 41246 41858 41298 41870
rect 41246 41794 41298 41806
rect 44494 41858 44546 41870
rect 57486 41858 57538 41870
rect 49858 41806 49870 41858
rect 49922 41806 49934 41858
rect 51986 41806 51998 41858
rect 52050 41806 52062 41858
rect 55906 41806 55918 41858
rect 55970 41806 55982 41858
rect 44494 41794 44546 41806
rect 57486 41794 57538 41806
rect 8990 41746 9042 41758
rect 8990 41682 9042 41694
rect 13806 41746 13858 41758
rect 24222 41746 24274 41758
rect 19954 41694 19966 41746
rect 20018 41694 20030 41746
rect 13806 41682 13858 41694
rect 24222 41682 24274 41694
rect 25678 41746 25730 41758
rect 25678 41682 25730 41694
rect 27694 41746 27746 41758
rect 27694 41682 27746 41694
rect 33406 41746 33458 41758
rect 33406 41682 33458 41694
rect 33742 41746 33794 41758
rect 43822 41746 43874 41758
rect 34626 41694 34638 41746
rect 34690 41694 34702 41746
rect 33742 41682 33794 41694
rect 43822 41682 43874 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 14030 41410 14082 41422
rect 27358 41410 27410 41422
rect 44158 41410 44210 41422
rect 27122 41358 27134 41410
rect 27186 41358 27198 41410
rect 32162 41358 32174 41410
rect 32226 41358 32238 41410
rect 33506 41358 33518 41410
rect 33570 41358 33582 41410
rect 14030 41346 14082 41358
rect 27358 41346 27410 41358
rect 44158 41346 44210 41358
rect 50318 41410 50370 41422
rect 50318 41346 50370 41358
rect 52894 41410 52946 41422
rect 52894 41346 52946 41358
rect 9998 41298 10050 41310
rect 20078 41298 20130 41310
rect 2706 41246 2718 41298
rect 2770 41246 2782 41298
rect 4498 41246 4510 41298
rect 4562 41246 4574 41298
rect 14690 41246 14702 41298
rect 14754 41246 14766 41298
rect 9998 41234 10050 41246
rect 20078 41234 20130 41246
rect 21310 41298 21362 41310
rect 23774 41298 23826 41310
rect 34862 41298 34914 41310
rect 23202 41246 23214 41298
rect 23266 41246 23278 41298
rect 25554 41246 25566 41298
rect 25618 41246 25630 41298
rect 32498 41246 32510 41298
rect 32562 41246 32574 41298
rect 21310 41234 21362 41246
rect 23774 41234 23826 41246
rect 34862 41234 34914 41246
rect 36990 41298 37042 41310
rect 36990 41234 37042 41246
rect 38558 41298 38610 41310
rect 43486 41298 43538 41310
rect 40114 41246 40126 41298
rect 40178 41246 40190 41298
rect 38558 41234 38610 41246
rect 43486 41234 43538 41246
rect 45166 41298 45218 41310
rect 52670 41298 52722 41310
rect 45490 41246 45502 41298
rect 45554 41246 45566 41298
rect 48626 41246 48638 41298
rect 48690 41246 48702 41298
rect 50530 41246 50542 41298
rect 50594 41246 50606 41298
rect 45166 41234 45218 41246
rect 52670 41234 52722 41246
rect 5518 41186 5570 41198
rect 12126 41186 12178 41198
rect 19854 41186 19906 41198
rect 25902 41186 25954 41198
rect 4050 41134 4062 41186
rect 4114 41134 4126 41186
rect 5170 41134 5182 41186
rect 5234 41134 5246 41186
rect 8642 41134 8654 41186
rect 8706 41134 8718 41186
rect 15810 41134 15822 41186
rect 15874 41134 15886 41186
rect 17378 41134 17390 41186
rect 17442 41134 17454 41186
rect 19058 41134 19070 41186
rect 19122 41134 19134 41186
rect 23314 41134 23326 41186
rect 23378 41134 23390 41186
rect 25218 41134 25230 41186
rect 25282 41134 25294 41186
rect 25442 41134 25454 41186
rect 25506 41134 25518 41186
rect 5518 41122 5570 41134
rect 12126 41122 12178 41134
rect 19854 41122 19906 41134
rect 25902 41122 25954 41134
rect 26574 41186 26626 41198
rect 26574 41122 26626 41134
rect 29038 41186 29090 41198
rect 34638 41186 34690 41198
rect 32050 41134 32062 41186
rect 32114 41134 32126 41186
rect 33170 41134 33182 41186
rect 33234 41134 33246 41186
rect 33506 41134 33518 41186
rect 33570 41134 33582 41186
rect 33954 41134 33966 41186
rect 34018 41134 34030 41186
rect 29038 41122 29090 41134
rect 34638 41122 34690 41134
rect 35534 41186 35586 41198
rect 35534 41122 35586 41134
rect 35758 41186 35810 41198
rect 37102 41186 37154 41198
rect 51662 41186 51714 41198
rect 36082 41134 36094 41186
rect 36146 41134 36158 41186
rect 37650 41134 37662 41186
rect 37714 41134 37726 41186
rect 43026 41134 43038 41186
rect 43090 41134 43102 41186
rect 50642 41134 50654 41186
rect 50706 41134 50718 41186
rect 35758 41122 35810 41134
rect 37102 41122 37154 41134
rect 51662 41122 51714 41134
rect 51886 41186 51938 41198
rect 51886 41122 51938 41134
rect 51998 41186 52050 41198
rect 51998 41122 52050 41134
rect 53118 41186 53170 41198
rect 55682 41134 55694 41186
rect 55746 41134 55758 41186
rect 57586 41134 57598 41186
rect 57650 41134 57662 41186
rect 53118 41122 53170 41134
rect 2830 41074 2882 41086
rect 2830 41010 2882 41022
rect 3054 41074 3106 41086
rect 5854 41074 5906 41086
rect 12350 41074 12402 41086
rect 3714 41022 3726 41074
rect 3778 41022 3790 41074
rect 9650 41022 9662 41074
rect 9714 41022 9726 41074
rect 3054 41010 3106 41022
rect 5854 41010 5906 41022
rect 12350 41010 12402 41022
rect 12462 41074 12514 41086
rect 12462 41010 12514 41022
rect 13470 41074 13522 41086
rect 13470 41010 13522 41022
rect 13918 41074 13970 41086
rect 20302 41074 20354 41086
rect 16370 41022 16382 41074
rect 16434 41022 16446 41074
rect 17490 41022 17502 41074
rect 17554 41022 17566 41074
rect 18834 41022 18846 41074
rect 18898 41022 18910 41074
rect 13918 41010 13970 41022
rect 20302 41010 20354 41022
rect 20526 41074 20578 41086
rect 20526 41010 20578 41022
rect 26462 41074 26514 41086
rect 26462 41010 26514 41022
rect 26686 41074 26738 41086
rect 26686 41010 26738 41022
rect 27918 41074 27970 41086
rect 27918 41010 27970 41022
rect 29374 41074 29426 41086
rect 29374 41010 29426 41022
rect 34750 41074 34802 41086
rect 44270 41074 44322 41086
rect 42242 41022 42254 41074
rect 42306 41022 42318 41074
rect 34750 41010 34802 41022
rect 44270 41010 44322 41022
rect 51550 41074 51602 41086
rect 55346 41022 55358 41074
rect 55410 41022 55422 41074
rect 57250 41022 57262 41074
rect 57314 41022 57326 41074
rect 51550 41010 51602 41022
rect 5742 40962 5794 40974
rect 13694 40962 13746 40974
rect 8306 40910 8318 40962
rect 8370 40910 8382 40962
rect 5742 40898 5794 40910
rect 13694 40898 13746 40910
rect 15150 40962 15202 40974
rect 15150 40898 15202 40910
rect 21870 40962 21922 40974
rect 21870 40898 21922 40910
rect 22318 40962 22370 40974
rect 22318 40898 22370 40910
rect 27470 40962 27522 40974
rect 27470 40898 27522 40910
rect 27694 40962 27746 40974
rect 27694 40898 27746 40910
rect 29262 40962 29314 40974
rect 29262 40898 29314 40910
rect 34974 40962 35026 40974
rect 34974 40898 35026 40910
rect 35086 40962 35138 40974
rect 35086 40898 35138 40910
rect 44158 40962 44210 40974
rect 44158 40898 44210 40910
rect 45390 40962 45442 40974
rect 45390 40898 45442 40910
rect 49086 40962 49138 40974
rect 49086 40898 49138 40910
rect 53566 40962 53618 40974
rect 56018 40910 56030 40962
rect 56082 40910 56094 40962
rect 53566 40898 53618 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 5070 40626 5122 40638
rect 14030 40626 14082 40638
rect 20414 40626 20466 40638
rect 2706 40574 2718 40626
rect 2770 40574 2782 40626
rect 8082 40574 8094 40626
rect 8146 40574 8158 40626
rect 19394 40574 19406 40626
rect 19458 40574 19470 40626
rect 5070 40562 5122 40574
rect 14030 40562 14082 40574
rect 20414 40562 20466 40574
rect 20974 40626 21026 40638
rect 20974 40562 21026 40574
rect 21422 40626 21474 40638
rect 21422 40562 21474 40574
rect 41134 40626 41186 40638
rect 41134 40562 41186 40574
rect 55694 40626 55746 40638
rect 55694 40562 55746 40574
rect 55918 40626 55970 40638
rect 55918 40562 55970 40574
rect 58158 40626 58210 40638
rect 58158 40562 58210 40574
rect 5294 40514 5346 40526
rect 17950 40514 18002 40526
rect 4274 40462 4286 40514
rect 4338 40462 4350 40514
rect 16706 40462 16718 40514
rect 16770 40462 16782 40514
rect 5294 40450 5346 40462
rect 17950 40450 18002 40462
rect 22878 40514 22930 40526
rect 38782 40514 38834 40526
rect 34850 40462 34862 40514
rect 34914 40462 34926 40514
rect 35634 40462 35646 40514
rect 35698 40462 35710 40514
rect 22878 40450 22930 40462
rect 38782 40450 38834 40462
rect 40238 40514 40290 40526
rect 40238 40450 40290 40462
rect 40350 40514 40402 40526
rect 44034 40462 44046 40514
rect 44098 40462 44110 40514
rect 45826 40462 45838 40514
rect 45890 40462 45902 40514
rect 56914 40462 56926 40514
rect 56978 40462 56990 40514
rect 40350 40450 40402 40462
rect 7758 40402 7810 40414
rect 17502 40402 17554 40414
rect 3042 40350 3054 40402
rect 3106 40350 3118 40402
rect 3938 40350 3950 40402
rect 4002 40350 4014 40402
rect 15026 40350 15038 40402
rect 15090 40350 15102 40402
rect 15810 40350 15822 40402
rect 15874 40350 15886 40402
rect 7758 40338 7810 40350
rect 17502 40338 17554 40350
rect 20302 40402 20354 40414
rect 23886 40402 23938 40414
rect 28926 40402 28978 40414
rect 23426 40350 23438 40402
rect 23490 40350 23502 40402
rect 27122 40350 27134 40402
rect 27186 40350 27198 40402
rect 27794 40350 27806 40402
rect 27858 40350 27870 40402
rect 20302 40338 20354 40350
rect 23886 40338 23938 40350
rect 28926 40338 28978 40350
rect 29262 40402 29314 40414
rect 40798 40402 40850 40414
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 34178 40350 34190 40402
rect 34242 40350 34254 40402
rect 35746 40350 35758 40402
rect 35810 40350 35822 40402
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 29262 40338 29314 40350
rect 40798 40338 40850 40350
rect 41246 40402 41298 40414
rect 41246 40338 41298 40350
rect 41358 40402 41410 40414
rect 56030 40402 56082 40414
rect 43810 40350 43822 40402
rect 43874 40350 43886 40402
rect 44594 40350 44606 40402
rect 44658 40350 44670 40402
rect 45042 40350 45054 40402
rect 45106 40350 45118 40402
rect 51650 40350 51662 40402
rect 51714 40350 51726 40402
rect 57026 40350 57038 40402
rect 57090 40350 57102 40402
rect 57474 40350 57486 40402
rect 57538 40350 57550 40402
rect 41358 40338 41410 40350
rect 56030 40338 56082 40350
rect 19182 40290 19234 40302
rect 31166 40290 31218 40302
rect 43598 40290 43650 40302
rect 50990 40290 51042 40302
rect 4946 40238 4958 40290
rect 5010 40238 5022 40290
rect 22978 40238 22990 40290
rect 23042 40238 23054 40290
rect 27570 40238 27582 40290
rect 27634 40238 27646 40290
rect 28018 40238 28030 40290
rect 28082 40238 28094 40290
rect 29474 40238 29486 40290
rect 29538 40238 29550 40290
rect 35858 40238 35870 40290
rect 35922 40238 35934 40290
rect 38098 40238 38110 40290
rect 38162 40238 38174 40290
rect 47954 40238 47966 40290
rect 48018 40238 48030 40290
rect 51762 40238 51774 40290
rect 51826 40238 51838 40290
rect 57250 40238 57262 40290
rect 57314 40238 57326 40290
rect 19182 40226 19234 40238
rect 31166 40226 31218 40238
rect 43598 40226 43650 40238
rect 50990 40226 51042 40238
rect 15150 40178 15202 40190
rect 20414 40178 20466 40190
rect 16482 40126 16494 40178
rect 16546 40126 16558 40178
rect 15150 40114 15202 40126
rect 20414 40114 20466 40126
rect 22654 40178 22706 40190
rect 22654 40114 22706 40126
rect 40238 40178 40290 40190
rect 40238 40114 40290 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 45838 39842 45890 39854
rect 14914 39790 14926 39842
rect 14978 39790 14990 39842
rect 26002 39790 26014 39842
rect 26066 39790 26078 39842
rect 45838 39778 45890 39790
rect 51326 39842 51378 39854
rect 51326 39778 51378 39790
rect 57486 39842 57538 39854
rect 57486 39778 57538 39790
rect 57822 39842 57874 39854
rect 57822 39778 57874 39790
rect 5070 39730 5122 39742
rect 2482 39678 2494 39730
rect 2546 39678 2558 39730
rect 4610 39678 4622 39730
rect 4674 39678 4686 39730
rect 5070 39666 5122 39678
rect 6862 39730 6914 39742
rect 6862 39666 6914 39678
rect 17726 39730 17778 39742
rect 17726 39666 17778 39678
rect 18846 39730 18898 39742
rect 18846 39666 18898 39678
rect 20750 39730 20802 39742
rect 32174 39730 32226 39742
rect 22194 39678 22206 39730
rect 22258 39678 22270 39730
rect 26114 39678 26126 39730
rect 26178 39678 26190 39730
rect 27906 39678 27918 39730
rect 27970 39678 27982 39730
rect 20750 39666 20802 39678
rect 32174 39666 32226 39678
rect 32510 39730 32562 39742
rect 32510 39666 32562 39678
rect 34638 39730 34690 39742
rect 47518 39730 47570 39742
rect 35186 39678 35198 39730
rect 35250 39678 35262 39730
rect 43362 39678 43374 39730
rect 43426 39678 43438 39730
rect 45266 39678 45278 39730
rect 45330 39678 45342 39730
rect 50978 39678 50990 39730
rect 51042 39678 51054 39730
rect 56466 39678 56478 39730
rect 56530 39678 56542 39730
rect 34638 39666 34690 39678
rect 47518 39666 47570 39678
rect 22654 39618 22706 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 11442 39566 11454 39618
rect 11506 39566 11518 39618
rect 12338 39566 12350 39618
rect 12402 39566 12414 39618
rect 14130 39566 14142 39618
rect 14194 39566 14206 39618
rect 14914 39566 14926 39618
rect 14978 39566 14990 39618
rect 15474 39566 15486 39618
rect 15538 39566 15550 39618
rect 17490 39566 17502 39618
rect 17554 39566 17566 39618
rect 18946 39566 18958 39618
rect 19010 39566 19022 39618
rect 19282 39566 19294 39618
rect 19346 39566 19358 39618
rect 22654 39554 22706 39566
rect 23774 39618 23826 39630
rect 31278 39618 31330 39630
rect 34862 39618 34914 39630
rect 25554 39566 25566 39618
rect 25618 39566 25630 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 26562 39566 26574 39618
rect 26626 39566 26638 39618
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 23774 39554 23826 39566
rect 31278 39554 31330 39566
rect 34862 39554 34914 39566
rect 41694 39618 41746 39630
rect 47406 39618 47458 39630
rect 43810 39566 43822 39618
rect 43874 39566 43886 39618
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 53666 39566 53678 39618
rect 53730 39566 53742 39618
rect 57026 39566 57038 39618
rect 57090 39566 57102 39618
rect 41694 39554 41746 39566
rect 47406 39554 47458 39566
rect 16494 39506 16546 39518
rect 12898 39454 12910 39506
rect 12962 39454 12974 39506
rect 16494 39442 16546 39454
rect 25006 39506 25058 39518
rect 25006 39442 25058 39454
rect 37550 39506 37602 39518
rect 37550 39442 37602 39454
rect 44270 39506 44322 39518
rect 44270 39442 44322 39454
rect 45054 39506 45106 39518
rect 45054 39442 45106 39454
rect 45726 39506 45778 39518
rect 45726 39442 45778 39454
rect 49310 39506 49362 39518
rect 57598 39506 57650 39518
rect 54338 39454 54350 39506
rect 54402 39454 54414 39506
rect 49310 39442 49362 39454
rect 57598 39442 57650 39454
rect 11678 39394 11730 39406
rect 17390 39394 17442 39406
rect 12562 39342 12574 39394
rect 12626 39342 12638 39394
rect 11678 39330 11730 39342
rect 17390 39330 17442 39342
rect 20190 39394 20242 39406
rect 20190 39330 20242 39342
rect 24110 39394 24162 39406
rect 24110 39330 24162 39342
rect 27470 39394 27522 39406
rect 27470 39330 27522 39342
rect 33070 39394 33122 39406
rect 33070 39330 33122 39342
rect 37886 39394 37938 39406
rect 37886 39330 37938 39342
rect 42254 39394 42306 39406
rect 42254 39330 42306 39342
rect 45838 39394 45890 39406
rect 45838 39330 45890 39342
rect 48974 39394 49026 39406
rect 48974 39330 49026 39342
rect 49758 39394 49810 39406
rect 49758 39330 49810 39342
rect 50654 39394 50706 39406
rect 50654 39330 50706 39342
rect 51102 39394 51154 39406
rect 56802 39342 56814 39394
rect 56866 39342 56878 39394
rect 51102 39330 51154 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 6190 39058 6242 39070
rect 6190 38994 6242 39006
rect 8206 39058 8258 39070
rect 27694 39058 27746 39070
rect 13010 39006 13022 39058
rect 13074 39006 13086 39058
rect 8206 38994 8258 39006
rect 27694 38994 27746 39006
rect 27918 39058 27970 39070
rect 27918 38994 27970 39006
rect 44718 39058 44770 39070
rect 44718 38994 44770 39006
rect 53566 39058 53618 39070
rect 53566 38994 53618 39006
rect 54126 39058 54178 39070
rect 54126 38994 54178 39006
rect 7870 38946 7922 38958
rect 7870 38882 7922 38894
rect 7982 38946 8034 38958
rect 7982 38882 8034 38894
rect 12014 38946 12066 38958
rect 12014 38882 12066 38894
rect 12238 38946 12290 38958
rect 20974 38946 21026 38958
rect 19842 38894 19854 38946
rect 19906 38894 19918 38946
rect 20402 38894 20414 38946
rect 20466 38894 20478 38946
rect 12238 38882 12290 38894
rect 20974 38882 21026 38894
rect 30382 38946 30434 38958
rect 36530 38894 36542 38946
rect 36594 38894 36606 38946
rect 38098 38894 38110 38946
rect 38162 38894 38174 38946
rect 38994 38894 39006 38946
rect 39058 38894 39070 38946
rect 50978 38894 50990 38946
rect 51042 38894 51054 38946
rect 57810 38894 57822 38946
rect 57874 38894 57886 38946
rect 30382 38882 30434 38894
rect 6414 38834 6466 38846
rect 6414 38770 6466 38782
rect 6638 38834 6690 38846
rect 11454 38834 11506 38846
rect 7074 38782 7086 38834
rect 7138 38782 7150 38834
rect 6638 38770 6690 38782
rect 11454 38770 11506 38782
rect 12462 38834 12514 38846
rect 12462 38770 12514 38782
rect 12574 38834 12626 38846
rect 18062 38834 18114 38846
rect 20750 38834 20802 38846
rect 15586 38782 15598 38834
rect 15650 38782 15662 38834
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 18498 38782 18510 38834
rect 18562 38782 18574 38834
rect 18834 38782 18846 38834
rect 18898 38782 18910 38834
rect 12574 38770 12626 38782
rect 18062 38770 18114 38782
rect 20750 38770 20802 38782
rect 23438 38834 23490 38846
rect 23438 38770 23490 38782
rect 23662 38834 23714 38846
rect 23662 38770 23714 38782
rect 23886 38834 23938 38846
rect 23886 38770 23938 38782
rect 24110 38834 24162 38846
rect 26350 38834 26402 38846
rect 28030 38834 28082 38846
rect 25666 38782 25678 38834
rect 25730 38782 25742 38834
rect 27010 38782 27022 38834
rect 27074 38782 27086 38834
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 24110 38770 24162 38782
rect 26350 38770 26402 38782
rect 28030 38770 28082 38782
rect 30046 38834 30098 38846
rect 30046 38770 30098 38782
rect 30606 38834 30658 38846
rect 30606 38770 30658 38782
rect 32510 38834 32562 38846
rect 48862 38834 48914 38846
rect 57598 38834 57650 38846
rect 34066 38782 34078 38834
rect 34130 38782 34142 38834
rect 34738 38782 34750 38834
rect 34802 38782 34814 38834
rect 36866 38782 36878 38834
rect 36930 38782 36942 38834
rect 37426 38782 37438 38834
rect 37490 38782 37502 38834
rect 39666 38782 39678 38834
rect 39730 38782 39742 38834
rect 40002 38782 40014 38834
rect 40066 38782 40078 38834
rect 50194 38782 50206 38834
rect 50258 38782 50270 38834
rect 58034 38782 58046 38834
rect 58098 38782 58110 38834
rect 32510 38770 32562 38782
rect 48862 38770 48914 38782
rect 57598 38770 57650 38782
rect 6526 38722 6578 38734
rect 6526 38658 6578 38670
rect 7534 38722 7586 38734
rect 7534 38658 7586 38670
rect 11678 38722 11730 38734
rect 29934 38722 29986 38734
rect 39230 38722 39282 38734
rect 15810 38670 15822 38722
rect 15874 38670 15886 38722
rect 18610 38670 18622 38722
rect 18674 38670 18686 38722
rect 25554 38670 25566 38722
rect 25618 38670 25630 38722
rect 32162 38670 32174 38722
rect 32226 38670 32238 38722
rect 34290 38670 34302 38722
rect 34354 38670 34366 38722
rect 34850 38670 34862 38722
rect 34914 38670 34926 38722
rect 11678 38658 11730 38670
rect 29934 38658 29986 38670
rect 39230 38658 39282 38670
rect 45950 38722 46002 38734
rect 45950 38658 46002 38670
rect 46174 38722 46226 38734
rect 46174 38658 46226 38670
rect 49422 38722 49474 38734
rect 53902 38722 53954 38734
rect 56702 38722 56754 38734
rect 53106 38670 53118 38722
rect 53170 38670 53182 38722
rect 54226 38670 54238 38722
rect 54290 38670 54302 38722
rect 49422 38658 49474 38670
rect 53902 38658 53954 38670
rect 56702 38658 56754 38670
rect 24222 38610 24274 38622
rect 30270 38610 30322 38622
rect 11106 38558 11118 38610
rect 11170 38558 11182 38610
rect 15362 38558 15374 38610
rect 15426 38558 15438 38610
rect 26786 38558 26798 38610
rect 26850 38558 26862 38610
rect 24222 38546 24274 38558
rect 30270 38546 30322 38558
rect 30830 38610 30882 38622
rect 31938 38558 31950 38610
rect 32002 38558 32014 38610
rect 46498 38558 46510 38610
rect 46562 38558 46574 38610
rect 30830 38546 30882 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 3950 38274 4002 38286
rect 3950 38210 4002 38222
rect 9886 38274 9938 38286
rect 9886 38210 9938 38222
rect 11790 38274 11842 38286
rect 12574 38274 12626 38286
rect 12226 38222 12238 38274
rect 12290 38222 12302 38274
rect 11790 38210 11842 38222
rect 12574 38210 12626 38222
rect 13694 38274 13746 38286
rect 13694 38210 13746 38222
rect 15374 38274 15426 38286
rect 24558 38274 24610 38286
rect 16706 38222 16718 38274
rect 16770 38222 16782 38274
rect 19058 38222 19070 38274
rect 19122 38222 19134 38274
rect 15374 38210 15426 38222
rect 24558 38210 24610 38222
rect 26014 38274 26066 38286
rect 26014 38210 26066 38222
rect 27358 38274 27410 38286
rect 27358 38210 27410 38222
rect 29262 38274 29314 38286
rect 29262 38210 29314 38222
rect 30494 38274 30546 38286
rect 30494 38210 30546 38222
rect 35534 38274 35586 38286
rect 35534 38210 35586 38222
rect 4510 38162 4562 38174
rect 4510 38098 4562 38110
rect 6750 38162 6802 38174
rect 6750 38098 6802 38110
rect 12798 38162 12850 38174
rect 16594 38110 16606 38162
rect 16658 38110 16670 38162
rect 18610 38110 18622 38162
rect 18674 38110 18686 38162
rect 27010 38110 27022 38162
rect 27074 38110 27086 38162
rect 28130 38110 28142 38162
rect 28194 38110 28206 38162
rect 38770 38110 38782 38162
rect 38834 38110 38846 38162
rect 46386 38110 46398 38162
rect 46450 38110 46462 38162
rect 58146 38110 58158 38162
rect 58210 38110 58222 38162
rect 12798 38098 12850 38110
rect 4062 38050 4114 38062
rect 4062 37986 4114 37998
rect 5854 38050 5906 38062
rect 5854 37986 5906 37998
rect 6190 38050 6242 38062
rect 6190 37986 6242 37998
rect 6414 38050 6466 38062
rect 9550 38050 9602 38062
rect 7186 37998 7198 38050
rect 7250 37998 7262 38050
rect 8866 37998 8878 38050
rect 8930 37998 8942 38050
rect 6414 37986 6466 37998
rect 9550 37986 9602 37998
rect 11454 38050 11506 38062
rect 11454 37986 11506 37998
rect 14030 38050 14082 38062
rect 24222 38050 24274 38062
rect 14802 37998 14814 38050
rect 14866 37998 14878 38050
rect 15362 37998 15374 38050
rect 15426 37998 15438 38050
rect 18498 37998 18510 38050
rect 18562 37998 18574 38050
rect 20738 37998 20750 38050
rect 20802 37998 20814 38050
rect 14030 37986 14082 37998
rect 24222 37986 24274 37998
rect 26126 38050 26178 38062
rect 41582 38050 41634 38062
rect 27122 37998 27134 38050
rect 27186 37998 27198 38050
rect 27458 37998 27470 38050
rect 27522 37998 27534 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 31266 37998 31278 38050
rect 31330 37998 31342 38050
rect 32946 37998 32958 38050
rect 33010 37998 33022 38050
rect 34402 37998 34414 38050
rect 34466 37998 34478 38050
rect 38098 37998 38110 38050
rect 38162 37998 38174 38050
rect 40226 37998 40238 38050
rect 40290 37998 40302 38050
rect 26126 37986 26178 37998
rect 41582 37986 41634 37998
rect 42142 38050 42194 38062
rect 42142 37986 42194 37998
rect 45390 38050 45442 38062
rect 45390 37986 45442 37998
rect 45838 38050 45890 38062
rect 54910 38050 54962 38062
rect 49298 37998 49310 38050
rect 49362 37998 49374 38050
rect 55346 37998 55358 38050
rect 55410 37998 55422 38050
rect 45838 37986 45890 37998
rect 54910 37986 54962 37998
rect 17054 37938 17106 37950
rect 23998 37938 24050 37950
rect 8754 37886 8766 37938
rect 8818 37886 8830 37938
rect 10658 37886 10670 37938
rect 10722 37886 10734 37938
rect 11218 37886 11230 37938
rect 11282 37886 11294 37938
rect 14690 37886 14702 37938
rect 14754 37886 14766 37938
rect 21298 37886 21310 37938
rect 21362 37886 21374 37938
rect 17054 37874 17106 37886
rect 23998 37874 24050 37886
rect 28142 37938 28194 37950
rect 28142 37874 28194 37886
rect 29262 37938 29314 37950
rect 29262 37874 29314 37886
rect 29374 37938 29426 37950
rect 29374 37874 29426 37886
rect 30606 37938 30658 37950
rect 35646 37938 35698 37950
rect 46062 37938 46114 37950
rect 31826 37886 31838 37938
rect 31890 37886 31902 37938
rect 35074 37886 35086 37938
rect 35138 37886 35150 37938
rect 37202 37886 37214 37938
rect 37266 37886 37278 37938
rect 37986 37886 37998 37938
rect 38050 37886 38062 37938
rect 38994 37886 39006 37938
rect 39058 37886 39070 37938
rect 48514 37886 48526 37938
rect 48578 37886 48590 37938
rect 56018 37886 56030 37938
rect 56082 37886 56094 37938
rect 30606 37874 30658 37886
rect 35646 37874 35698 37886
rect 46062 37874 46114 37886
rect 3950 37826 4002 37838
rect 3950 37762 4002 37774
rect 5966 37826 6018 37838
rect 5966 37762 6018 37774
rect 21646 37826 21698 37838
rect 21646 37762 21698 37774
rect 22206 37826 22258 37838
rect 22206 37762 22258 37774
rect 26014 37826 26066 37838
rect 26014 37762 26066 37774
rect 28366 37826 28418 37838
rect 28366 37762 28418 37774
rect 30158 37826 30210 37838
rect 30158 37762 30210 37774
rect 30494 37826 30546 37838
rect 30494 37762 30546 37774
rect 30830 37826 30882 37838
rect 30830 37762 30882 37774
rect 35534 37826 35586 37838
rect 45278 37826 45330 37838
rect 37426 37774 37438 37826
rect 37490 37774 37502 37826
rect 40786 37774 40798 37826
rect 40850 37774 40862 37826
rect 35534 37762 35586 37774
rect 45278 37762 45330 37774
rect 45950 37826 46002 37838
rect 45950 37762 46002 37774
rect 49758 37826 49810 37838
rect 49758 37762 49810 37774
rect 53566 37826 53618 37838
rect 53566 37762 53618 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 3614 37490 3666 37502
rect 15150 37490 15202 37502
rect 12674 37438 12686 37490
rect 12738 37438 12750 37490
rect 3614 37426 3666 37438
rect 15150 37426 15202 37438
rect 15486 37490 15538 37502
rect 15486 37426 15538 37438
rect 24558 37490 24610 37502
rect 24558 37426 24610 37438
rect 25342 37490 25394 37502
rect 39006 37490 39058 37502
rect 30706 37438 30718 37490
rect 30770 37438 30782 37490
rect 37090 37438 37102 37490
rect 37154 37438 37166 37490
rect 25342 37426 25394 37438
rect 39006 37426 39058 37438
rect 39902 37490 39954 37502
rect 39902 37426 39954 37438
rect 44270 37490 44322 37502
rect 44270 37426 44322 37438
rect 46622 37490 46674 37502
rect 46622 37426 46674 37438
rect 46734 37490 46786 37502
rect 46734 37426 46786 37438
rect 56702 37490 56754 37502
rect 56702 37426 56754 37438
rect 2718 37378 2770 37390
rect 2718 37314 2770 37326
rect 3054 37378 3106 37390
rect 8654 37378 8706 37390
rect 5282 37326 5294 37378
rect 5346 37326 5358 37378
rect 8530 37326 8542 37378
rect 8594 37326 8606 37378
rect 3054 37314 3106 37326
rect 8654 37314 8706 37326
rect 8766 37378 8818 37390
rect 8766 37314 8818 37326
rect 9886 37378 9938 37390
rect 9886 37314 9938 37326
rect 11342 37378 11394 37390
rect 14814 37378 14866 37390
rect 12002 37326 12014 37378
rect 12066 37326 12078 37378
rect 12450 37326 12462 37378
rect 12514 37326 12526 37378
rect 11342 37314 11394 37326
rect 14814 37314 14866 37326
rect 14926 37378 14978 37390
rect 23662 37378 23714 37390
rect 18274 37326 18286 37378
rect 18338 37326 18350 37378
rect 18946 37326 18958 37378
rect 19010 37326 19022 37378
rect 14926 37314 14978 37326
rect 23662 37314 23714 37326
rect 26014 37378 26066 37390
rect 26014 37314 26066 37326
rect 26126 37378 26178 37390
rect 35758 37378 35810 37390
rect 39566 37378 39618 37390
rect 26786 37326 26798 37378
rect 26850 37326 26862 37378
rect 37202 37326 37214 37378
rect 37266 37326 37278 37378
rect 37762 37326 37774 37378
rect 37826 37326 37838 37378
rect 26126 37314 26178 37326
rect 35758 37314 35810 37326
rect 39566 37314 39618 37326
rect 39678 37378 39730 37390
rect 39678 37314 39730 37326
rect 46510 37378 46562 37390
rect 46510 37314 46562 37326
rect 3166 37266 3218 37278
rect 3166 37202 3218 37214
rect 3726 37266 3778 37278
rect 3726 37202 3778 37214
rect 3838 37266 3890 37278
rect 3838 37202 3890 37214
rect 4286 37266 4338 37278
rect 7870 37266 7922 37278
rect 4610 37214 4622 37266
rect 4674 37214 4686 37266
rect 4286 37202 4338 37214
rect 7870 37202 7922 37214
rect 8990 37266 9042 37278
rect 8990 37202 9042 37214
rect 9438 37266 9490 37278
rect 9438 37202 9490 37214
rect 10222 37266 10274 37278
rect 15486 37266 15538 37278
rect 11890 37214 11902 37266
rect 11954 37214 11966 37266
rect 10222 37202 10274 37214
rect 15486 37202 15538 37214
rect 15598 37266 15650 37278
rect 27134 37266 27186 37278
rect 31278 37266 31330 37278
rect 16370 37214 16382 37266
rect 16434 37214 16446 37266
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 17938 37214 17950 37266
rect 18002 37214 18014 37266
rect 19618 37214 19630 37266
rect 19682 37214 19694 37266
rect 20402 37214 20414 37266
rect 20466 37214 20478 37266
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 24658 37214 24670 37266
rect 24722 37214 24734 37266
rect 26562 37214 26574 37266
rect 26626 37214 26638 37266
rect 27570 37214 27582 37266
rect 27634 37214 27646 37266
rect 29138 37214 29150 37266
rect 29202 37214 29214 37266
rect 15598 37202 15650 37214
rect 27134 37202 27186 37214
rect 31278 37202 31330 37214
rect 33518 37266 33570 37278
rect 33518 37202 33570 37214
rect 33854 37266 33906 37278
rect 35970 37214 35982 37266
rect 36034 37214 36046 37266
rect 37986 37214 37998 37266
rect 38050 37214 38062 37266
rect 39218 37214 39230 37266
rect 39282 37214 39294 37266
rect 43810 37214 43822 37266
rect 43874 37214 43886 37266
rect 33854 37202 33906 37214
rect 2830 37154 2882 37166
rect 15822 37154 15874 37166
rect 22878 37154 22930 37166
rect 7410 37102 7422 37154
rect 7474 37102 7486 37154
rect 8754 37102 8766 37154
rect 8818 37102 8830 37154
rect 16706 37102 16718 37154
rect 16770 37102 16782 37154
rect 18386 37102 18398 37154
rect 18450 37102 18462 37154
rect 19730 37102 19742 37154
rect 19794 37102 19806 37154
rect 20738 37102 20750 37154
rect 20802 37102 20814 37154
rect 2830 37090 2882 37102
rect 15822 37090 15874 37102
rect 22878 37090 22930 37102
rect 25230 37154 25282 37166
rect 34066 37102 34078 37154
rect 34130 37102 34142 37154
rect 40898 37102 40910 37154
rect 40962 37102 40974 37154
rect 43026 37102 43038 37154
rect 43090 37102 43102 37154
rect 25230 37090 25282 37102
rect 31054 37042 31106 37054
rect 11106 36990 11118 37042
rect 11170 36990 11182 37042
rect 27234 36990 27246 37042
rect 27298 36990 27310 37042
rect 31054 36978 31106 36990
rect 38894 37042 38946 37054
rect 38894 36978 38946 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 8878 36706 8930 36718
rect 23102 36706 23154 36718
rect 16146 36654 16158 36706
rect 16210 36654 16222 36706
rect 16930 36654 16942 36706
rect 16994 36654 17006 36706
rect 8878 36642 8930 36654
rect 23102 36642 23154 36654
rect 24558 36706 24610 36718
rect 35646 36706 35698 36718
rect 27346 36654 27358 36706
rect 27410 36654 27422 36706
rect 24558 36642 24610 36654
rect 35646 36642 35698 36654
rect 36878 36706 36930 36718
rect 36878 36642 36930 36654
rect 40910 36706 40962 36718
rect 40910 36642 40962 36654
rect 41246 36706 41298 36718
rect 41246 36642 41298 36654
rect 5182 36594 5234 36606
rect 2482 36542 2494 36594
rect 2546 36542 2558 36594
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 5182 36530 5234 36542
rect 9326 36594 9378 36606
rect 22542 36594 22594 36606
rect 12002 36542 12014 36594
rect 12066 36542 12078 36594
rect 15922 36542 15934 36594
rect 15986 36542 15998 36594
rect 16818 36542 16830 36594
rect 16882 36542 16894 36594
rect 18498 36542 18510 36594
rect 18562 36542 18574 36594
rect 9326 36530 9378 36542
rect 22542 36530 22594 36542
rect 24110 36594 24162 36606
rect 37886 36594 37938 36606
rect 52894 36594 52946 36606
rect 28242 36542 28254 36594
rect 28306 36542 28318 36594
rect 30706 36542 30718 36594
rect 30770 36542 30782 36594
rect 35522 36542 35534 36594
rect 35586 36542 35598 36594
rect 52098 36542 52110 36594
rect 52162 36542 52174 36594
rect 56130 36542 56142 36594
rect 56194 36542 56206 36594
rect 24110 36530 24162 36542
rect 37886 36530 37938 36542
rect 52894 36530 52946 36542
rect 11118 36482 11170 36494
rect 22766 36482 22818 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 11442 36430 11454 36482
rect 11506 36430 11518 36482
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 15698 36430 15710 36482
rect 15762 36430 15774 36482
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 17490 36430 17502 36482
rect 17554 36430 17566 36482
rect 18834 36430 18846 36482
rect 18898 36430 18910 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 11118 36418 11170 36430
rect 22766 36418 22818 36430
rect 23998 36482 24050 36494
rect 23998 36418 24050 36430
rect 24334 36482 24386 36494
rect 24334 36418 24386 36430
rect 24670 36482 24722 36494
rect 27246 36482 27298 36494
rect 33294 36482 33346 36494
rect 37102 36482 37154 36494
rect 26898 36430 26910 36482
rect 26962 36430 26974 36482
rect 31490 36430 31502 36482
rect 31554 36430 31566 36482
rect 35410 36430 35422 36482
rect 35474 36430 35486 36482
rect 36082 36430 36094 36482
rect 36146 36430 36158 36482
rect 24670 36418 24722 36430
rect 27246 36418 27298 36430
rect 33294 36418 33346 36430
rect 37102 36418 37154 36430
rect 37550 36482 37602 36494
rect 37550 36418 37602 36430
rect 37662 36482 37714 36494
rect 57038 36482 57090 36494
rect 38546 36430 38558 36482
rect 38610 36430 38622 36482
rect 49298 36430 49310 36482
rect 49362 36430 49374 36482
rect 53330 36430 53342 36482
rect 53394 36430 53406 36482
rect 37662 36418 37714 36430
rect 57038 36418 57090 36430
rect 57374 36482 57426 36494
rect 57374 36418 57426 36430
rect 8766 36370 8818 36382
rect 23662 36370 23714 36382
rect 11554 36318 11566 36370
rect 11618 36318 11630 36370
rect 19058 36318 19070 36370
rect 19122 36318 19134 36370
rect 8766 36306 8818 36318
rect 23662 36306 23714 36318
rect 32062 36370 32114 36382
rect 32062 36306 32114 36318
rect 38222 36370 38274 36382
rect 38222 36306 38274 36318
rect 44046 36370 44098 36382
rect 56702 36370 56754 36382
rect 49970 36318 49982 36370
rect 50034 36318 50046 36370
rect 54002 36318 54014 36370
rect 54066 36318 54078 36370
rect 44046 36306 44098 36318
rect 56702 36306 56754 36318
rect 8878 36258 8930 36270
rect 8878 36194 8930 36206
rect 9886 36258 9938 36270
rect 9886 36194 9938 36206
rect 10782 36258 10834 36270
rect 10782 36194 10834 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 12686 36258 12738 36270
rect 12686 36194 12738 36206
rect 21310 36258 21362 36270
rect 27806 36258 27858 36270
rect 21634 36206 21646 36258
rect 21698 36206 21710 36258
rect 21310 36194 21362 36206
rect 27806 36194 27858 36206
rect 31166 36258 31218 36270
rect 31166 36194 31218 36206
rect 32958 36258 33010 36270
rect 32958 36194 33010 36206
rect 41134 36258 41186 36270
rect 41134 36194 41186 36206
rect 41694 36258 41746 36270
rect 41694 36194 41746 36206
rect 43822 36258 43874 36270
rect 43822 36194 43874 36206
rect 43934 36258 43986 36270
rect 43934 36194 43986 36206
rect 57150 36258 57202 36270
rect 57150 36194 57202 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 11678 35922 11730 35934
rect 11678 35858 11730 35870
rect 15598 35922 15650 35934
rect 15598 35858 15650 35870
rect 18958 35922 19010 35934
rect 18958 35858 19010 35870
rect 23326 35922 23378 35934
rect 25230 35922 25282 35934
rect 24210 35870 24222 35922
rect 24274 35870 24286 35922
rect 23326 35858 23378 35870
rect 25230 35858 25282 35870
rect 27246 35922 27298 35934
rect 27246 35858 27298 35870
rect 28366 35922 28418 35934
rect 38222 35922 38274 35934
rect 31490 35870 31502 35922
rect 31554 35870 31566 35922
rect 37650 35870 37662 35922
rect 37714 35870 37726 35922
rect 28366 35858 28418 35870
rect 38222 35858 38274 35870
rect 39006 35922 39058 35934
rect 39006 35858 39058 35870
rect 39230 35922 39282 35934
rect 39230 35858 39282 35870
rect 50430 35922 50482 35934
rect 50430 35858 50482 35870
rect 51214 35922 51266 35934
rect 51214 35858 51266 35870
rect 55134 35922 55186 35934
rect 55134 35858 55186 35870
rect 56702 35922 56754 35934
rect 56702 35858 56754 35870
rect 57262 35922 57314 35934
rect 57262 35858 57314 35870
rect 57486 35922 57538 35934
rect 57486 35858 57538 35870
rect 57822 35922 57874 35934
rect 57822 35858 57874 35870
rect 58046 35922 58098 35934
rect 58046 35858 58098 35870
rect 17950 35810 18002 35822
rect 17950 35746 18002 35758
rect 27358 35810 27410 35822
rect 32398 35810 32450 35822
rect 30930 35758 30942 35810
rect 30994 35758 31006 35810
rect 27358 35746 27410 35758
rect 32398 35746 32450 35758
rect 34974 35810 35026 35822
rect 38334 35810 38386 35822
rect 51998 35810 52050 35822
rect 37202 35758 37214 35810
rect 37266 35758 37278 35810
rect 37426 35758 37438 35810
rect 37490 35758 37502 35810
rect 44818 35758 44830 35810
rect 44882 35758 44894 35810
rect 34974 35746 35026 35758
rect 38334 35746 38386 35758
rect 51998 35746 52050 35758
rect 11342 35698 11394 35710
rect 1810 35646 1822 35698
rect 1874 35646 1886 35698
rect 11342 35634 11394 35646
rect 11678 35698 11730 35710
rect 11678 35634 11730 35646
rect 12014 35698 12066 35710
rect 12014 35634 12066 35646
rect 16158 35698 16210 35710
rect 16158 35634 16210 35646
rect 18846 35698 18898 35710
rect 18846 35634 18898 35646
rect 20302 35698 20354 35710
rect 20302 35634 20354 35646
rect 22766 35698 22818 35710
rect 32510 35698 32562 35710
rect 23986 35646 23998 35698
rect 24050 35646 24062 35698
rect 30482 35646 30494 35698
rect 30546 35646 30558 35698
rect 31378 35646 31390 35698
rect 31442 35646 31454 35698
rect 22766 35634 22818 35646
rect 32510 35634 32562 35646
rect 35870 35698 35922 35710
rect 35870 35634 35922 35646
rect 37886 35698 37938 35710
rect 38894 35698 38946 35710
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 37886 35634 37938 35646
rect 38894 35634 38946 35646
rect 39342 35698 39394 35710
rect 39342 35634 39394 35646
rect 42478 35698 42530 35710
rect 52894 35698 52946 35710
rect 45490 35646 45502 35698
rect 45554 35646 45566 35698
rect 50642 35646 50654 35698
rect 50706 35646 50718 35698
rect 42478 35634 42530 35646
rect 52894 35634 52946 35646
rect 54910 35698 54962 35710
rect 54910 35634 54962 35646
rect 55358 35698 55410 35710
rect 55358 35634 55410 35646
rect 55582 35698 55634 35710
rect 55582 35634 55634 35646
rect 56478 35698 56530 35710
rect 56478 35634 56530 35646
rect 56814 35698 56866 35710
rect 56814 35634 56866 35646
rect 57150 35698 57202 35710
rect 57150 35634 57202 35646
rect 57710 35698 57762 35710
rect 57710 35634 57762 35646
rect 2270 35586 2322 35598
rect 2270 35522 2322 35534
rect 19182 35586 19234 35598
rect 21310 35586 21362 35598
rect 33630 35586 33682 35598
rect 20738 35534 20750 35586
rect 20802 35534 20814 35586
rect 25666 35534 25678 35586
rect 25730 35534 25742 35586
rect 19182 35522 19234 35534
rect 21310 35522 21362 35534
rect 33630 35522 33682 35534
rect 34190 35586 34242 35598
rect 42690 35534 42702 35586
rect 42754 35534 42766 35586
rect 51986 35534 51998 35586
rect 52050 35534 52062 35586
rect 34190 35522 34242 35534
rect 15934 35474 15986 35486
rect 15934 35410 15986 35422
rect 32398 35474 32450 35486
rect 32398 35410 32450 35422
rect 50318 35474 50370 35486
rect 51774 35474 51826 35486
rect 50866 35422 50878 35474
rect 50930 35471 50942 35474
rect 51202 35471 51214 35474
rect 50930 35425 51214 35471
rect 50930 35422 50942 35425
rect 51202 35422 51214 35425
rect 51266 35422 51278 35474
rect 50318 35410 50370 35422
rect 51774 35410 51826 35422
rect 53118 35474 53170 35486
rect 53118 35410 53170 35422
rect 53454 35474 53506 35486
rect 53454 35410 53506 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 12126 35138 12178 35150
rect 44942 35138 44994 35150
rect 10434 35086 10446 35138
rect 10498 35086 10510 35138
rect 14242 35086 14254 35138
rect 14306 35086 14318 35138
rect 17266 35086 17278 35138
rect 17330 35086 17342 35138
rect 12126 35074 12178 35086
rect 44942 35074 44994 35086
rect 1822 35026 1874 35038
rect 19070 35026 19122 35038
rect 20862 35026 20914 35038
rect 29710 35026 29762 35038
rect 35758 35026 35810 35038
rect 8642 34974 8654 35026
rect 8706 34974 8718 35026
rect 15810 34974 15822 35026
rect 15874 34974 15886 35026
rect 19506 34974 19518 35026
rect 19570 34974 19582 35026
rect 24210 34974 24222 35026
rect 24274 34974 24286 35026
rect 27906 34974 27918 35026
rect 27970 34974 27982 35026
rect 33730 34974 33742 35026
rect 33794 34974 33806 35026
rect 1822 34962 1874 34974
rect 19070 34962 19122 34974
rect 20862 34962 20914 34974
rect 29710 34962 29762 34974
rect 35758 34962 35810 34974
rect 37662 35026 37714 35038
rect 44046 35026 44098 35038
rect 38210 34974 38222 35026
rect 38274 34974 38286 35026
rect 37662 34962 37714 34974
rect 44046 34962 44098 34974
rect 45502 35026 45554 35038
rect 49982 35026 50034 35038
rect 46050 34974 46062 35026
rect 46114 34974 46126 35026
rect 45502 34962 45554 34974
rect 49982 34962 50034 34974
rect 7870 34914 7922 34926
rect 7870 34850 7922 34862
rect 8206 34914 8258 34926
rect 11454 34914 11506 34926
rect 8418 34862 8430 34914
rect 8482 34862 8494 34914
rect 9538 34862 9550 34914
rect 9602 34862 9614 34914
rect 9986 34862 9998 34914
rect 10050 34862 10062 34914
rect 10546 34862 10558 34914
rect 10610 34862 10622 34914
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 8206 34850 8258 34862
rect 11454 34850 11506 34862
rect 12574 34914 12626 34926
rect 16270 34914 16322 34926
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 12574 34850 12626 34862
rect 16270 34850 16322 34862
rect 16606 34914 16658 34926
rect 17838 34914 17890 34926
rect 29822 34914 29874 34926
rect 16818 34862 16830 34914
rect 16882 34862 16894 34914
rect 19954 34862 19966 34914
rect 20018 34862 20030 34914
rect 21298 34862 21310 34914
rect 21362 34862 21374 34914
rect 30146 34862 30158 34914
rect 30210 34862 30222 34914
rect 36194 34862 36206 34914
rect 36258 34862 36270 34914
rect 37202 34862 37214 34914
rect 37266 34862 37278 34914
rect 38322 34862 38334 34914
rect 38386 34862 38398 34914
rect 48850 34862 48862 34914
rect 48914 34862 48926 34914
rect 53218 34862 53230 34914
rect 53282 34862 53294 34914
rect 16606 34850 16658 34862
rect 17838 34850 17890 34862
rect 29822 34850 29874 34862
rect 12910 34802 12962 34814
rect 8754 34750 8766 34802
rect 8818 34750 8830 34802
rect 12910 34738 12962 34750
rect 13694 34802 13746 34814
rect 13694 34738 13746 34750
rect 13806 34802 13858 34814
rect 13806 34738 13858 34750
rect 17950 34802 18002 34814
rect 17950 34738 18002 34750
rect 18510 34802 18562 34814
rect 37998 34802 38050 34814
rect 22082 34750 22094 34802
rect 22146 34750 22158 34802
rect 18510 34738 18562 34750
rect 37998 34738 38050 34750
rect 43598 34802 43650 34814
rect 43598 34738 43650 34750
rect 43822 34802 43874 34814
rect 43822 34738 43874 34750
rect 44158 34802 44210 34814
rect 44158 34738 44210 34750
rect 44942 34802 44994 34814
rect 49422 34802 49474 34814
rect 44942 34738 44994 34750
rect 45054 34746 45106 34758
rect 48178 34750 48190 34802
rect 48242 34750 48254 34802
rect 7982 34690 8034 34702
rect 7982 34626 8034 34638
rect 11790 34690 11842 34702
rect 11790 34626 11842 34638
rect 12014 34690 12066 34702
rect 12014 34626 12066 34638
rect 12686 34690 12738 34702
rect 12686 34626 12738 34638
rect 28366 34690 28418 34702
rect 28366 34626 28418 34638
rect 29374 34690 29426 34702
rect 29374 34626 29426 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 38782 34690 38834 34702
rect 49422 34738 49474 34750
rect 49534 34802 49586 34814
rect 49534 34738 49586 34750
rect 56926 34802 56978 34814
rect 56926 34738 56978 34750
rect 57038 34802 57090 34814
rect 57038 34738 57090 34750
rect 45054 34682 45106 34694
rect 56702 34690 56754 34702
rect 53442 34638 53454 34690
rect 53506 34638 53518 34690
rect 38782 34626 38834 34638
rect 56702 34626 56754 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 9662 34354 9714 34366
rect 18622 34354 18674 34366
rect 11106 34302 11118 34354
rect 11170 34302 11182 34354
rect 9662 34290 9714 34302
rect 18622 34290 18674 34302
rect 29150 34354 29202 34366
rect 29150 34290 29202 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 30046 34354 30098 34366
rect 30046 34290 30098 34302
rect 34078 34354 34130 34366
rect 34078 34290 34130 34302
rect 41470 34354 41522 34366
rect 44270 34354 44322 34366
rect 42354 34302 42366 34354
rect 42418 34302 42430 34354
rect 41470 34290 41522 34302
rect 44270 34290 44322 34302
rect 44494 34354 44546 34366
rect 44494 34290 44546 34302
rect 54686 34354 54738 34366
rect 54686 34290 54738 34302
rect 30270 34242 30322 34254
rect 34638 34242 34690 34254
rect 10546 34190 10558 34242
rect 10610 34190 10622 34242
rect 10770 34190 10782 34242
rect 10834 34190 10846 34242
rect 14802 34190 14814 34242
rect 14866 34190 14878 34242
rect 30930 34190 30942 34242
rect 30994 34190 31006 34242
rect 31378 34190 31390 34242
rect 31442 34190 31454 34242
rect 30270 34178 30322 34190
rect 34638 34178 34690 34190
rect 35982 34242 36034 34254
rect 35982 34178 36034 34190
rect 37102 34242 37154 34254
rect 37102 34178 37154 34190
rect 47182 34242 47234 34254
rect 47182 34178 47234 34190
rect 54910 34242 54962 34254
rect 54910 34178 54962 34190
rect 56702 34242 56754 34254
rect 56702 34178 56754 34190
rect 11342 34130 11394 34142
rect 18286 34130 18338 34142
rect 8530 34078 8542 34130
rect 8594 34078 8606 34130
rect 9874 34078 9886 34130
rect 9938 34078 9950 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 12226 34078 12238 34130
rect 12290 34078 12302 34130
rect 13906 34078 13918 34130
rect 13970 34078 13982 34130
rect 17826 34078 17838 34130
rect 17890 34078 17902 34130
rect 11342 34066 11394 34078
rect 18286 34066 18338 34078
rect 19182 34130 19234 34142
rect 28702 34130 28754 34142
rect 23874 34078 23886 34130
rect 23938 34078 23950 34130
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 19182 34066 19234 34078
rect 28702 34066 28754 34078
rect 28926 34130 28978 34142
rect 28926 34066 28978 34078
rect 30382 34130 30434 34142
rect 34190 34130 34242 34142
rect 36766 34130 36818 34142
rect 30706 34078 30718 34130
rect 30770 34078 30782 34130
rect 31826 34078 31838 34130
rect 31890 34078 31902 34130
rect 36530 34078 36542 34130
rect 36594 34078 36606 34130
rect 30382 34066 30434 34078
rect 34190 34066 34242 34078
rect 36766 34066 36818 34078
rect 37438 34130 37490 34142
rect 37438 34066 37490 34078
rect 38782 34130 38834 34142
rect 40350 34130 40402 34142
rect 39218 34078 39230 34130
rect 39282 34078 39294 34130
rect 38782 34066 38834 34078
rect 40350 34066 40402 34078
rect 41022 34130 41074 34142
rect 41022 34066 41074 34078
rect 41694 34130 41746 34142
rect 41694 34066 41746 34078
rect 42030 34130 42082 34142
rect 42030 34066 42082 34078
rect 43934 34130 43986 34142
rect 43934 34066 43986 34078
rect 44606 34130 44658 34142
rect 44606 34066 44658 34078
rect 45726 34130 45778 34142
rect 55022 34130 55074 34142
rect 45938 34078 45950 34130
rect 46002 34078 46014 34130
rect 45726 34066 45778 34078
rect 55022 34066 55074 34078
rect 57038 34130 57090 34142
rect 57038 34066 57090 34078
rect 57262 34130 57314 34142
rect 57262 34066 57314 34078
rect 28814 34018 28866 34030
rect 33854 34018 33906 34030
rect 8866 33966 8878 34018
rect 8930 33966 8942 34018
rect 14466 33966 14478 34018
rect 14530 33966 14542 34018
rect 23538 33966 23550 34018
rect 23602 33966 23614 34018
rect 25442 33966 25454 34018
rect 25506 33966 25518 34018
rect 27570 33966 27582 34018
rect 27634 33966 27646 34018
rect 31602 33966 31614 34018
rect 31666 33966 31678 34018
rect 28814 33954 28866 33966
rect 33854 33954 33906 33966
rect 37326 34018 37378 34030
rect 39678 34018 39730 34030
rect 38322 33966 38334 34018
rect 38386 33966 38398 34018
rect 37326 33954 37378 33966
rect 39678 33954 39730 33966
rect 41582 34018 41634 34030
rect 41582 33954 41634 33966
rect 46622 34018 46674 34030
rect 46622 33954 46674 33966
rect 46958 34018 47010 34030
rect 47742 34018 47794 34030
rect 47282 33966 47294 34018
rect 47346 33966 47358 34018
rect 46958 33954 47010 33966
rect 47742 33954 47794 33966
rect 56814 34018 56866 34030
rect 56814 33954 56866 33966
rect 9550 33906 9602 33918
rect 9550 33842 9602 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 12798 33570 12850 33582
rect 12798 33506 12850 33518
rect 57038 33570 57090 33582
rect 57038 33506 57090 33518
rect 57598 33570 57650 33582
rect 57598 33506 57650 33518
rect 27918 33458 27970 33470
rect 13906 33406 13918 33458
rect 13970 33406 13982 33458
rect 18050 33406 18062 33458
rect 18114 33406 18126 33458
rect 24210 33406 24222 33458
rect 24274 33406 24286 33458
rect 51202 33406 51214 33458
rect 51266 33406 51278 33458
rect 55570 33406 55582 33458
rect 55634 33406 55646 33458
rect 27918 33394 27970 33406
rect 18846 33346 18898 33358
rect 11666 33294 11678 33346
rect 11730 33294 11742 33346
rect 12226 33294 12238 33346
rect 12290 33294 12302 33346
rect 12786 33294 12798 33346
rect 12850 33294 12862 33346
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 18846 33282 18898 33294
rect 19630 33346 19682 33358
rect 19630 33282 19682 33294
rect 20078 33346 20130 33358
rect 28142 33346 28194 33358
rect 21410 33294 21422 33346
rect 21474 33294 21486 33346
rect 22082 33294 22094 33346
rect 22146 33294 22158 33346
rect 20078 33282 20130 33294
rect 28142 33282 28194 33294
rect 28366 33346 28418 33358
rect 28366 33282 28418 33294
rect 31278 33346 31330 33358
rect 34302 33346 34354 33358
rect 39790 33346 39842 33358
rect 41694 33346 41746 33358
rect 31826 33294 31838 33346
rect 31890 33294 31902 33346
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 35074 33294 35086 33346
rect 35138 33294 35150 33346
rect 36978 33294 36990 33346
rect 37042 33294 37054 33346
rect 38434 33294 38446 33346
rect 38498 33294 38510 33346
rect 38882 33294 38894 33346
rect 38946 33294 38958 33346
rect 40226 33294 40238 33346
rect 40290 33294 40302 33346
rect 41234 33294 41246 33346
rect 41298 33294 41310 33346
rect 31278 33282 31330 33294
rect 34302 33282 34354 33294
rect 39790 33282 39842 33294
rect 41694 33282 41746 33294
rect 42030 33346 42082 33358
rect 42030 33282 42082 33294
rect 42366 33346 42418 33358
rect 51886 33346 51938 33358
rect 57486 33346 57538 33358
rect 43922 33294 43934 33346
rect 43986 33294 43998 33346
rect 48290 33294 48302 33346
rect 48354 33294 48366 33346
rect 52770 33294 52782 33346
rect 52834 33294 52846 33346
rect 42366 33282 42418 33294
rect 51886 33282 51938 33294
rect 57486 33282 57538 33294
rect 18510 33234 18562 33246
rect 15922 33182 15934 33234
rect 15986 33182 15998 33234
rect 18510 33170 18562 33182
rect 18622 33234 18674 33246
rect 18622 33170 18674 33182
rect 19070 33234 19122 33246
rect 27806 33234 27858 33246
rect 38110 33234 38162 33246
rect 51550 33234 51602 33246
rect 25778 33182 25790 33234
rect 25842 33182 25854 33234
rect 32386 33182 32398 33234
rect 32450 33182 32462 33234
rect 39106 33182 39118 33234
rect 39170 33182 39182 33234
rect 43698 33182 43710 33234
rect 43762 33182 43774 33234
rect 49074 33182 49086 33234
rect 49138 33182 49150 33234
rect 19070 33170 19122 33182
rect 27806 33170 27858 33182
rect 38110 33170 38162 33182
rect 51550 33170 51602 33182
rect 51998 33234 52050 33246
rect 51998 33170 52050 33182
rect 52110 33234 52162 33246
rect 57150 33234 57202 33246
rect 53442 33182 53454 33234
rect 53506 33182 53518 33234
rect 52110 33170 52162 33182
rect 57150 33170 57202 33182
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 14814 33122 14866 33134
rect 14814 33058 14866 33070
rect 19406 33122 19458 33134
rect 19406 33058 19458 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 20526 33122 20578 33134
rect 20526 33058 20578 33070
rect 24670 33122 24722 33134
rect 24670 33058 24722 33070
rect 25118 33122 25170 33134
rect 25118 33058 25170 33070
rect 25454 33122 25506 33134
rect 25454 33058 25506 33070
rect 27582 33122 27634 33134
rect 27582 33058 27634 33070
rect 29486 33122 29538 33134
rect 31502 33122 31554 33134
rect 30930 33070 30942 33122
rect 30994 33070 31006 33122
rect 29486 33058 29538 33070
rect 31502 33058 31554 33070
rect 36206 33122 36258 33134
rect 36206 33058 36258 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 42030 33122 42082 33134
rect 42030 33058 42082 33070
rect 56030 33122 56082 33134
rect 56030 33058 56082 33070
rect 57038 33122 57090 33134
rect 57038 33058 57090 33070
rect 57598 33122 57650 33134
rect 57598 33058 57650 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 13134 32786 13186 32798
rect 8978 32734 8990 32786
rect 9042 32734 9054 32786
rect 13134 32722 13186 32734
rect 18734 32786 18786 32798
rect 18734 32722 18786 32734
rect 24110 32786 24162 32798
rect 34078 32786 34130 32798
rect 24434 32734 24446 32786
rect 24498 32734 24510 32786
rect 32050 32734 32062 32786
rect 32114 32734 32126 32786
rect 24110 32722 24162 32734
rect 34078 32722 34130 32734
rect 38110 32786 38162 32798
rect 38110 32722 38162 32734
rect 39342 32786 39394 32798
rect 39342 32722 39394 32734
rect 43374 32786 43426 32798
rect 43374 32722 43426 32734
rect 49086 32786 49138 32798
rect 49086 32722 49138 32734
rect 51774 32786 51826 32798
rect 51774 32722 51826 32734
rect 53902 32786 53954 32798
rect 55122 32734 55134 32786
rect 55186 32734 55198 32786
rect 53902 32722 53954 32734
rect 11006 32674 11058 32686
rect 11006 32610 11058 32622
rect 13022 32674 13074 32686
rect 13022 32610 13074 32622
rect 50654 32674 50706 32686
rect 50654 32610 50706 32622
rect 51998 32674 52050 32686
rect 51998 32610 52050 32622
rect 52110 32674 52162 32686
rect 52110 32610 52162 32622
rect 52894 32674 52946 32686
rect 52894 32610 52946 32622
rect 53230 32674 53282 32686
rect 53230 32610 53282 32622
rect 54014 32674 54066 32686
rect 54014 32610 54066 32622
rect 54798 32674 54850 32686
rect 54798 32610 54850 32622
rect 9550 32562 9602 32574
rect 8754 32510 8766 32562
rect 8818 32510 8830 32562
rect 9550 32498 9602 32510
rect 10894 32562 10946 32574
rect 10894 32498 10946 32510
rect 11454 32562 11506 32574
rect 11454 32498 11506 32510
rect 12462 32562 12514 32574
rect 31726 32562 31778 32574
rect 34190 32562 34242 32574
rect 38446 32562 38498 32574
rect 12786 32510 12798 32562
rect 12850 32510 12862 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 33954 32510 33966 32562
rect 34018 32510 34030 32562
rect 34962 32510 34974 32562
rect 35026 32510 35038 32562
rect 37202 32510 37214 32562
rect 37266 32510 37278 32562
rect 12462 32498 12514 32510
rect 31726 32498 31778 32510
rect 34190 32498 34242 32510
rect 38446 32498 38498 32510
rect 39902 32562 39954 32574
rect 39902 32498 39954 32510
rect 43934 32562 43986 32574
rect 43934 32498 43986 32510
rect 44158 32562 44210 32574
rect 44942 32562 44994 32574
rect 47406 32562 47458 32574
rect 44482 32510 44494 32562
rect 44546 32510 44558 32562
rect 46722 32510 46734 32562
rect 46786 32510 46798 32562
rect 44158 32498 44210 32510
rect 44942 32498 44994 32510
rect 47406 32498 47458 32510
rect 48974 32562 49026 32574
rect 48974 32498 49026 32510
rect 49198 32562 49250 32574
rect 49198 32498 49250 32510
rect 49646 32562 49698 32574
rect 49646 32498 49698 32510
rect 50318 32562 50370 32574
rect 50318 32498 50370 32510
rect 50430 32562 50482 32574
rect 50430 32498 50482 32510
rect 50878 32562 50930 32574
rect 50878 32498 50930 32510
rect 18622 32450 18674 32462
rect 9874 32398 9886 32450
rect 9938 32398 9950 32450
rect 18622 32386 18674 32398
rect 19406 32450 19458 32462
rect 19406 32386 19458 32398
rect 20190 32450 20242 32462
rect 20190 32386 20242 32398
rect 28590 32450 28642 32462
rect 28590 32386 28642 32398
rect 31054 32450 31106 32462
rect 43598 32450 43650 32462
rect 31490 32398 31502 32450
rect 31554 32398 31566 32450
rect 34514 32398 34526 32450
rect 34578 32398 34590 32450
rect 36866 32398 36878 32450
rect 36930 32398 36942 32450
rect 37650 32398 37662 32450
rect 37714 32398 37726 32450
rect 38882 32398 38894 32450
rect 38946 32398 38958 32450
rect 31054 32386 31106 32398
rect 43598 32386 43650 32398
rect 44046 32450 44098 32462
rect 51438 32450 51490 32462
rect 46498 32398 46510 32450
rect 46562 32398 46574 32450
rect 44046 32386 44098 32398
rect 51438 32386 51490 32398
rect 58158 32450 58210 32462
rect 58158 32386 58210 32398
rect 43262 32338 43314 32350
rect 43262 32274 43314 32286
rect 53902 32338 53954 32350
rect 53902 32274 53954 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 9326 32002 9378 32014
rect 12238 32002 12290 32014
rect 10770 31950 10782 32002
rect 10834 31950 10846 32002
rect 9326 31938 9378 31950
rect 12238 31938 12290 31950
rect 35758 32002 35810 32014
rect 44046 32002 44098 32014
rect 43698 31950 43710 32002
rect 43762 31950 43774 32002
rect 49858 31950 49870 32002
rect 49922 31950 49934 32002
rect 35758 31938 35810 31950
rect 44046 31938 44098 31950
rect 8542 31890 8594 31902
rect 8542 31826 8594 31838
rect 10334 31890 10386 31902
rect 15038 31890 15090 31902
rect 31838 31890 31890 31902
rect 14242 31838 14254 31890
rect 14306 31838 14318 31890
rect 18274 31838 18286 31890
rect 18338 31838 18350 31890
rect 19058 31838 19070 31890
rect 19122 31838 19134 31890
rect 26786 31838 26798 31890
rect 26850 31838 26862 31890
rect 10334 31826 10386 31838
rect 15038 31826 15090 31838
rect 31838 31826 31890 31838
rect 34750 31890 34802 31902
rect 37886 31890 37938 31902
rect 42142 31890 42194 31902
rect 48750 31890 48802 31902
rect 37090 31838 37102 31890
rect 37154 31838 37166 31890
rect 39554 31838 39566 31890
rect 39618 31838 39630 31890
rect 41682 31838 41694 31890
rect 41746 31838 41758 31890
rect 45378 31838 45390 31890
rect 45442 31838 45454 31890
rect 56018 31838 56030 31890
rect 56082 31838 56094 31890
rect 58146 31838 58158 31890
rect 58210 31838 58222 31890
rect 34750 31826 34802 31838
rect 37886 31826 37938 31838
rect 42142 31826 42194 31838
rect 48750 31826 48802 31838
rect 8430 31778 8482 31790
rect 18622 31778 18674 31790
rect 34302 31778 34354 31790
rect 10434 31726 10446 31778
rect 10498 31726 10510 31778
rect 11330 31726 11342 31778
rect 11394 31726 11406 31778
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14018 31726 14030 31778
rect 14082 31726 14094 31778
rect 15362 31726 15374 31778
rect 15426 31726 15438 31778
rect 23874 31726 23886 31778
rect 23938 31726 23950 31778
rect 32050 31726 32062 31778
rect 32114 31726 32126 31778
rect 34178 31726 34190 31778
rect 34242 31726 34254 31778
rect 8430 31714 8482 31726
rect 18622 31714 18674 31726
rect 34302 31714 34354 31726
rect 35422 31778 35474 31790
rect 35422 31714 35474 31726
rect 37550 31778 37602 31790
rect 37550 31714 37602 31726
rect 37998 31778 38050 31790
rect 44270 31778 44322 31790
rect 49310 31778 49362 31790
rect 38882 31726 38894 31778
rect 38946 31726 38958 31778
rect 48290 31726 48302 31778
rect 48354 31726 48366 31778
rect 49522 31726 49534 31778
rect 49586 31726 49598 31778
rect 50082 31726 50094 31778
rect 50146 31726 50158 31778
rect 55234 31726 55246 31778
rect 55298 31726 55310 31778
rect 37998 31714 38050 31726
rect 44270 31714 44322 31726
rect 49310 31714 49362 31726
rect 8094 31666 8146 31678
rect 8094 31602 8146 31614
rect 8654 31666 8706 31678
rect 8654 31602 8706 31614
rect 8990 31666 9042 31678
rect 8990 31602 9042 31614
rect 12574 31666 12626 31678
rect 33070 31666 33122 31678
rect 14130 31614 14142 31666
rect 14194 31614 14206 31666
rect 16146 31614 16158 31666
rect 16210 31614 16222 31666
rect 24658 31614 24670 31666
rect 24722 31614 24734 31666
rect 12574 31602 12626 31614
rect 33070 31602 33122 31614
rect 35198 31666 35250 31678
rect 49422 31666 49474 31678
rect 47506 31614 47518 31666
rect 47570 31614 47582 31666
rect 35198 31602 35250 31614
rect 49422 31602 49474 31614
rect 9214 31554 9266 31566
rect 9214 31490 9266 31502
rect 12350 31554 12402 31566
rect 12350 31490 12402 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 32062 31554 32114 31566
rect 50766 31554 50818 31566
rect 50418 31502 50430 31554
rect 50482 31502 50494 31554
rect 32062 31490 32114 31502
rect 50766 31490 50818 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 22766 31218 22818 31230
rect 9874 31166 9886 31218
rect 9938 31166 9950 31218
rect 12450 31166 12462 31218
rect 12514 31166 12526 31218
rect 22766 31154 22818 31166
rect 23326 31218 23378 31230
rect 23326 31154 23378 31166
rect 24110 31218 24162 31230
rect 32062 31218 32114 31230
rect 31042 31166 31054 31218
rect 31106 31166 31118 31218
rect 24110 31154 24162 31166
rect 32062 31154 32114 31166
rect 34862 31218 34914 31230
rect 34862 31154 34914 31166
rect 35870 31218 35922 31230
rect 35870 31154 35922 31166
rect 49086 31218 49138 31230
rect 49086 31154 49138 31166
rect 56926 31218 56978 31230
rect 56926 31154 56978 31166
rect 13470 31106 13522 31118
rect 13470 31042 13522 31054
rect 21982 31106 22034 31118
rect 21982 31042 22034 31054
rect 22094 31106 22146 31118
rect 22094 31042 22146 31054
rect 22206 31106 22258 31118
rect 22206 31042 22258 31054
rect 35310 31106 35362 31118
rect 49982 31106 50034 31118
rect 43026 31054 43038 31106
rect 43090 31054 43102 31106
rect 35310 31042 35362 31054
rect 49982 31042 50034 31054
rect 55358 31106 55410 31118
rect 55358 31042 55410 31054
rect 57822 31106 57874 31118
rect 57822 31042 57874 31054
rect 58158 31106 58210 31118
rect 58158 31042 58210 31054
rect 7646 30994 7698 31006
rect 8878 30994 8930 31006
rect 22318 30994 22370 31006
rect 8530 30942 8542 30994
rect 8594 30942 8606 30994
rect 9874 30942 9886 30994
rect 9938 30942 9950 30994
rect 10210 30942 10222 30994
rect 10274 30942 10286 30994
rect 11442 30942 11454 30994
rect 11506 30942 11518 30994
rect 12898 30942 12910 30994
rect 12962 30942 12974 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 7646 30930 7698 30942
rect 8878 30930 8930 30942
rect 22318 30930 22370 30942
rect 22542 30994 22594 31006
rect 22542 30930 22594 30942
rect 22878 30994 22930 31006
rect 22878 30930 22930 30942
rect 23102 30994 23154 31006
rect 23102 30930 23154 30942
rect 23438 30994 23490 31006
rect 23438 30930 23490 30942
rect 23998 30994 24050 31006
rect 23998 30930 24050 30942
rect 24334 30994 24386 31006
rect 56590 30994 56642 31006
rect 28130 30942 28142 30994
rect 28194 30942 28206 30994
rect 42354 30942 42366 30994
rect 42418 30942 42430 30994
rect 55122 30942 55134 30994
rect 55186 30942 55198 30994
rect 24334 30930 24386 30942
rect 56590 30930 56642 30942
rect 56814 30994 56866 31006
rect 56814 30930 56866 30942
rect 57262 30994 57314 31006
rect 57262 30930 57314 30942
rect 8206 30882 8258 30894
rect 12686 30882 12738 30894
rect 9762 30830 9774 30882
rect 9826 30830 9838 30882
rect 11106 30830 11118 30882
rect 11170 30830 11182 30882
rect 8206 30818 8258 30830
rect 12686 30818 12738 30830
rect 21198 30882 21250 30894
rect 21198 30818 21250 30830
rect 25454 30882 25506 30894
rect 25454 30818 25506 30830
rect 27694 30882 27746 30894
rect 45614 30882 45666 30894
rect 50206 30882 50258 30894
rect 28802 30830 28814 30882
rect 28866 30830 28878 30882
rect 31602 30830 31614 30882
rect 31666 30830 31678 30882
rect 45154 30830 45166 30882
rect 45218 30830 45230 30882
rect 49858 30830 49870 30882
rect 49922 30830 49934 30882
rect 27694 30818 27746 30830
rect 45614 30818 45666 30830
rect 50206 30818 50258 30830
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 46510 30434 46562 30446
rect 46510 30370 46562 30382
rect 9214 30322 9266 30334
rect 9214 30258 9266 30270
rect 11118 30322 11170 30334
rect 19170 30270 19182 30322
rect 19234 30270 19246 30322
rect 21522 30270 21534 30322
rect 21586 30270 21598 30322
rect 24994 30270 25006 30322
rect 25058 30270 25070 30322
rect 28578 30270 28590 30322
rect 28642 30270 28654 30322
rect 29138 30270 29150 30322
rect 29202 30270 29214 30322
rect 39890 30270 39902 30322
rect 39954 30270 39966 30322
rect 46946 30270 46958 30322
rect 47010 30270 47022 30322
rect 56018 30270 56030 30322
rect 56082 30270 56094 30322
rect 58146 30270 58158 30322
rect 58210 30270 58222 30322
rect 11118 30258 11170 30270
rect 14814 30210 14866 30222
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 12898 30158 12910 30210
rect 12962 30158 12974 30210
rect 13570 30158 13582 30210
rect 13634 30158 13646 30210
rect 13794 30158 13806 30210
rect 13858 30158 13870 30210
rect 14130 30158 14142 30210
rect 14194 30158 14206 30210
rect 14814 30146 14866 30158
rect 19630 30210 19682 30222
rect 19630 30146 19682 30158
rect 22318 30210 22370 30222
rect 30158 30210 30210 30222
rect 25778 30158 25790 30210
rect 25842 30158 25854 30210
rect 22318 30146 22370 30158
rect 30158 30146 30210 30158
rect 34078 30210 34130 30222
rect 34078 30146 34130 30158
rect 34638 30210 34690 30222
rect 46622 30210 46674 30222
rect 50206 30210 50258 30222
rect 37090 30158 37102 30210
rect 37154 30158 37166 30210
rect 49858 30158 49870 30210
rect 49922 30158 49934 30210
rect 34638 30146 34690 30158
rect 46622 30146 46674 30158
rect 50206 30146 50258 30158
rect 50878 30210 50930 30222
rect 52670 30210 52722 30222
rect 51538 30158 51550 30210
rect 51602 30158 51614 30210
rect 55346 30158 55358 30210
rect 55410 30158 55422 30210
rect 50878 30146 50930 30158
rect 52670 30146 52722 30158
rect 7982 30098 8034 30110
rect 7982 30034 8034 30046
rect 9774 30098 9826 30110
rect 9774 30034 9826 30046
rect 11902 30098 11954 30110
rect 21982 30098 22034 30110
rect 21746 30046 21758 30098
rect 21810 30046 21822 30098
rect 11902 30034 11954 30046
rect 21982 30034 22034 30046
rect 22094 30098 22146 30110
rect 22094 30034 22146 30046
rect 24222 30098 24274 30110
rect 24222 30034 24274 30046
rect 24558 30098 24610 30110
rect 29598 30098 29650 30110
rect 24770 30046 24782 30098
rect 24834 30046 24846 30098
rect 26450 30046 26462 30098
rect 26514 30046 26526 30098
rect 29474 30046 29486 30098
rect 29538 30046 29550 30098
rect 24558 30034 24610 30046
rect 29598 30034 29650 30046
rect 30382 30098 30434 30110
rect 30382 30034 30434 30046
rect 30494 30098 30546 30110
rect 30494 30034 30546 30046
rect 31278 30098 31330 30110
rect 31278 30034 31330 30046
rect 35422 30098 35474 30110
rect 50318 30098 50370 30110
rect 37762 30046 37774 30098
rect 37826 30046 37838 30098
rect 49074 30046 49086 30098
rect 49138 30046 49150 30098
rect 35422 30034 35474 30046
rect 50318 30034 50370 30046
rect 51774 30098 51826 30110
rect 51774 30034 51826 30046
rect 12798 29986 12850 29998
rect 12798 29922 12850 29934
rect 15598 29986 15650 29998
rect 15598 29922 15650 29934
rect 22878 29986 22930 29998
rect 22878 29922 22930 29934
rect 24446 29986 24498 29998
rect 24446 29922 24498 29934
rect 29710 29986 29762 29998
rect 29710 29922 29762 29934
rect 29934 29986 29986 29998
rect 29934 29922 29986 29934
rect 31390 29986 31442 29998
rect 31390 29922 31442 29934
rect 31614 29986 31666 29998
rect 31614 29922 31666 29934
rect 35086 29986 35138 29998
rect 35086 29922 35138 29934
rect 35758 29986 35810 29998
rect 35758 29922 35810 29934
rect 40350 29986 40402 29998
rect 40350 29922 40402 29934
rect 46510 29986 46562 29998
rect 46510 29922 46562 29934
rect 50542 29986 50594 29998
rect 50542 29922 50594 29934
rect 53006 29986 53058 29998
rect 53006 29922 53058 29934
rect 54574 29986 54626 29998
rect 54898 29934 54910 29986
rect 54962 29934 54974 29986
rect 54574 29922 54626 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 16606 29650 16658 29662
rect 16606 29586 16658 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 18062 29650 18114 29662
rect 18062 29586 18114 29598
rect 21870 29650 21922 29662
rect 21870 29586 21922 29598
rect 22318 29650 22370 29662
rect 23214 29650 23266 29662
rect 25566 29650 25618 29662
rect 22866 29598 22878 29650
rect 22930 29598 22942 29650
rect 24322 29598 24334 29650
rect 24386 29598 24398 29650
rect 22318 29586 22370 29598
rect 23214 29586 23266 29598
rect 25566 29586 25618 29598
rect 26910 29650 26962 29662
rect 26910 29586 26962 29598
rect 27806 29650 27858 29662
rect 27806 29586 27858 29598
rect 28702 29650 28754 29662
rect 28702 29586 28754 29598
rect 30830 29650 30882 29662
rect 30830 29586 30882 29598
rect 31838 29650 31890 29662
rect 31838 29586 31890 29598
rect 37214 29650 37266 29662
rect 37214 29586 37266 29598
rect 42926 29650 42978 29662
rect 51102 29650 51154 29662
rect 43474 29598 43486 29650
rect 43538 29598 43550 29650
rect 42926 29586 42978 29598
rect 51102 29586 51154 29598
rect 53118 29650 53170 29662
rect 53118 29586 53170 29598
rect 56702 29650 56754 29662
rect 56702 29586 56754 29598
rect 56926 29650 56978 29662
rect 56926 29586 56978 29598
rect 57822 29650 57874 29662
rect 57822 29586 57874 29598
rect 14814 29538 14866 29550
rect 8978 29486 8990 29538
rect 9042 29486 9054 29538
rect 14814 29474 14866 29486
rect 16494 29538 16546 29550
rect 16494 29474 16546 29486
rect 17278 29538 17330 29550
rect 17278 29474 17330 29486
rect 21534 29538 21586 29550
rect 21534 29474 21586 29486
rect 21646 29538 21698 29550
rect 21646 29474 21698 29486
rect 22094 29538 22146 29550
rect 22094 29474 22146 29486
rect 22430 29538 22482 29550
rect 22430 29474 22482 29486
rect 23662 29538 23714 29550
rect 27694 29538 27746 29550
rect 25218 29486 25230 29538
rect 25282 29486 25294 29538
rect 27570 29486 27582 29538
rect 27634 29486 27646 29538
rect 23662 29474 23714 29486
rect 27694 29474 27746 29486
rect 28478 29538 28530 29550
rect 36990 29538 37042 29550
rect 31154 29486 31166 29538
rect 31218 29486 31230 29538
rect 28478 29474 28530 29486
rect 36990 29474 37042 29486
rect 51550 29538 51602 29550
rect 57038 29538 57090 29550
rect 53442 29486 53454 29538
rect 53506 29486 53518 29538
rect 51550 29474 51602 29486
rect 57038 29474 57090 29486
rect 8318 29426 8370 29438
rect 14590 29426 14642 29438
rect 16830 29426 16882 29438
rect 4386 29374 4398 29426
rect 4450 29374 4462 29426
rect 8754 29374 8766 29426
rect 8818 29374 8830 29426
rect 11218 29374 11230 29426
rect 11282 29374 11294 29426
rect 12002 29374 12014 29426
rect 12066 29374 12078 29426
rect 13010 29374 13022 29426
rect 13074 29374 13086 29426
rect 14242 29374 14254 29426
rect 14306 29374 14318 29426
rect 15026 29374 15038 29426
rect 15090 29374 15102 29426
rect 15362 29374 15374 29426
rect 15426 29374 15438 29426
rect 16034 29374 16046 29426
rect 16098 29374 16110 29426
rect 8318 29362 8370 29374
rect 14590 29362 14642 29374
rect 16830 29362 16882 29374
rect 17614 29426 17666 29438
rect 23998 29426 24050 29438
rect 28030 29426 28082 29438
rect 21074 29374 21086 29426
rect 21138 29374 21150 29426
rect 24546 29374 24558 29426
rect 24610 29374 24622 29426
rect 17614 29362 17666 29374
rect 23998 29362 24050 29374
rect 28030 29362 28082 29374
rect 28814 29426 28866 29438
rect 28814 29362 28866 29374
rect 30606 29426 30658 29438
rect 36878 29426 36930 29438
rect 31042 29374 31054 29426
rect 31106 29374 31118 29426
rect 35634 29374 35646 29426
rect 35698 29374 35710 29426
rect 30606 29362 30658 29374
rect 36878 29362 36930 29374
rect 37438 29426 37490 29438
rect 37438 29362 37490 29374
rect 50990 29426 51042 29438
rect 50990 29362 51042 29374
rect 51214 29426 51266 29438
rect 51214 29362 51266 29374
rect 14702 29314 14754 29326
rect 20750 29314 20802 29326
rect 29262 29314 29314 29326
rect 5058 29262 5070 29314
rect 5122 29262 5134 29314
rect 7186 29262 7198 29314
rect 7250 29262 7262 29314
rect 7858 29262 7870 29314
rect 7922 29262 7934 29314
rect 10434 29262 10446 29314
rect 10498 29262 10510 29314
rect 13906 29262 13918 29314
rect 13970 29262 13982 29314
rect 16482 29262 16494 29314
rect 16546 29262 16558 29314
rect 21522 29262 21534 29314
rect 21586 29262 21598 29314
rect 27682 29262 27694 29314
rect 27746 29262 27758 29314
rect 14702 29250 14754 29262
rect 20750 29250 20802 29262
rect 29262 29250 29314 29262
rect 29710 29314 29762 29326
rect 40238 29314 40290 29326
rect 31378 29262 31390 29314
rect 31442 29262 31454 29314
rect 35970 29262 35982 29314
rect 36034 29262 36046 29314
rect 29710 29250 29762 29262
rect 40238 29250 40290 29262
rect 44046 29314 44098 29326
rect 44046 29250 44098 29262
rect 53902 29314 53954 29326
rect 53902 29250 53954 29262
rect 58158 29314 58210 29326
rect 58158 29250 58210 29262
rect 40126 29202 40178 29214
rect 40126 29138 40178 29150
rect 42814 29202 42866 29214
rect 42814 29138 42866 29150
rect 43150 29202 43202 29214
rect 43150 29138 43202 29150
rect 43822 29202 43874 29214
rect 43822 29138 43874 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 12014 28866 12066 28878
rect 29026 28814 29038 28866
rect 29090 28863 29102 28866
rect 29362 28863 29374 28866
rect 29090 28817 29374 28863
rect 29090 28814 29102 28817
rect 29362 28814 29374 28817
rect 29426 28814 29438 28866
rect 12014 28802 12066 28814
rect 8094 28754 8146 28766
rect 15934 28754 15986 28766
rect 29374 28754 29426 28766
rect 36430 28754 36482 28766
rect 9986 28702 9998 28754
rect 10050 28702 10062 28754
rect 19618 28702 19630 28754
rect 19682 28702 19694 28754
rect 31938 28702 31950 28754
rect 32002 28702 32014 28754
rect 34066 28702 34078 28754
rect 34130 28702 34142 28754
rect 34850 28702 34862 28754
rect 34914 28702 34926 28754
rect 8094 28690 8146 28702
rect 15934 28690 15986 28702
rect 29374 28690 29426 28702
rect 36430 28690 36482 28702
rect 37886 28754 37938 28766
rect 41918 28754 41970 28766
rect 41458 28702 41470 28754
rect 41522 28702 41534 28754
rect 37886 28690 37938 28702
rect 41918 28690 41970 28702
rect 43486 28754 43538 28766
rect 43486 28690 43538 28702
rect 45278 28754 45330 28766
rect 49534 28754 49586 28766
rect 48514 28702 48526 28754
rect 48578 28702 48590 28754
rect 45278 28690 45330 28702
rect 49534 28690 49586 28702
rect 49758 28754 49810 28766
rect 49758 28690 49810 28702
rect 50654 28754 50706 28766
rect 56578 28702 56590 28754
rect 56642 28702 56654 28754
rect 50654 28690 50706 28702
rect 12350 28642 12402 28654
rect 7634 28590 7646 28642
rect 7698 28590 7710 28642
rect 9314 28590 9326 28642
rect 9378 28590 9390 28642
rect 10994 28590 11006 28642
rect 11058 28590 11070 28642
rect 12350 28578 12402 28590
rect 13918 28642 13970 28654
rect 15150 28642 15202 28654
rect 30270 28642 30322 28654
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 16818 28590 16830 28642
rect 16882 28590 16894 28642
rect 28130 28590 28142 28642
rect 28194 28590 28206 28642
rect 13918 28578 13970 28590
rect 15150 28578 15202 28590
rect 30270 28578 30322 28590
rect 30606 28642 30658 28654
rect 30606 28578 30658 28590
rect 30942 28642 30994 28654
rect 35310 28642 35362 28654
rect 31154 28590 31166 28642
rect 31218 28590 31230 28642
rect 30942 28578 30994 28590
rect 35310 28578 35362 28590
rect 35870 28642 35922 28654
rect 35870 28578 35922 28590
rect 37326 28642 37378 28654
rect 42702 28642 42754 28654
rect 38658 28590 38670 28642
rect 38722 28590 38734 28642
rect 37326 28578 37378 28590
rect 42702 28578 42754 28590
rect 42926 28642 42978 28654
rect 52670 28642 52722 28654
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 42926 28578 42978 28590
rect 52670 28578 52722 28590
rect 53230 28642 53282 28654
rect 54450 28590 54462 28642
rect 54514 28590 54526 28642
rect 53230 28578 53282 28590
rect 12574 28530 12626 28542
rect 10434 28478 10446 28530
rect 10498 28478 10510 28530
rect 12574 28466 12626 28478
rect 14142 28530 14194 28542
rect 14142 28466 14194 28478
rect 14254 28530 14306 28542
rect 14254 28466 14306 28478
rect 16158 28530 16210 28542
rect 16158 28466 16210 28478
rect 16270 28530 16322 28542
rect 30718 28530 30770 28542
rect 17490 28478 17502 28530
rect 17554 28478 17566 28530
rect 28354 28478 28366 28530
rect 28418 28478 28430 28530
rect 16270 28466 16322 28478
rect 30718 28466 30770 28478
rect 37774 28530 37826 28542
rect 53566 28530 53618 28542
rect 39330 28478 39342 28530
rect 39394 28478 39406 28530
rect 46386 28478 46398 28530
rect 46450 28478 46462 28530
rect 52994 28478 53006 28530
rect 53058 28478 53070 28530
rect 37774 28466 37826 28478
rect 53566 28466 53618 28478
rect 7198 28418 7250 28430
rect 7198 28354 7250 28366
rect 14030 28418 14082 28430
rect 14030 28354 14082 28366
rect 16494 28418 16546 28430
rect 16494 28354 16546 28366
rect 34414 28418 34466 28430
rect 34414 28354 34466 28366
rect 37102 28418 37154 28430
rect 37102 28354 37154 28366
rect 37998 28418 38050 28430
rect 37998 28354 38050 28366
rect 43374 28418 43426 28430
rect 43374 28354 43426 28366
rect 43598 28418 43650 28430
rect 53454 28418 53506 28430
rect 50082 28366 50094 28418
rect 50146 28366 50158 28418
rect 43598 28354 43650 28366
rect 53454 28354 53506 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 11454 28082 11506 28094
rect 11454 28018 11506 28030
rect 11790 28082 11842 28094
rect 11790 28018 11842 28030
rect 12798 28082 12850 28094
rect 12798 28018 12850 28030
rect 14142 28082 14194 28094
rect 14142 28018 14194 28030
rect 14926 28082 14978 28094
rect 14926 28018 14978 28030
rect 16382 28082 16434 28094
rect 16382 28018 16434 28030
rect 17390 28082 17442 28094
rect 17390 28018 17442 28030
rect 17502 28082 17554 28094
rect 19182 28082 19234 28094
rect 28926 28082 28978 28094
rect 18834 28030 18846 28082
rect 18898 28030 18910 28082
rect 28466 28030 28478 28082
rect 28530 28030 28542 28082
rect 17502 28018 17554 28030
rect 19182 28018 19234 28030
rect 28926 28018 28978 28030
rect 30830 28082 30882 28094
rect 30830 28018 30882 28030
rect 34526 28082 34578 28094
rect 38894 28082 38946 28094
rect 36082 28030 36094 28082
rect 36146 28030 36158 28082
rect 34526 28018 34578 28030
rect 38894 28018 38946 28030
rect 44382 28082 44434 28094
rect 44382 28018 44434 28030
rect 54686 28082 54738 28094
rect 54686 28018 54738 28030
rect 56590 28082 56642 28094
rect 56590 28018 56642 28030
rect 57374 28082 57426 28094
rect 57374 28018 57426 28030
rect 10446 27970 10498 27982
rect 5506 27918 5518 27970
rect 5570 27918 5582 27970
rect 10446 27906 10498 27918
rect 14366 27970 14418 27982
rect 14366 27906 14418 27918
rect 17614 27970 17666 27982
rect 17614 27906 17666 27918
rect 17726 27970 17778 27982
rect 31054 27970 31106 27982
rect 20290 27918 20302 27970
rect 20354 27918 20366 27970
rect 17726 27906 17778 27918
rect 31054 27906 31106 27918
rect 32062 27970 32114 27982
rect 32062 27906 32114 27918
rect 38110 27970 38162 27982
rect 38110 27906 38162 27918
rect 38222 27970 38274 27982
rect 38222 27906 38274 27918
rect 38446 27970 38498 27982
rect 38446 27906 38498 27918
rect 39006 27970 39058 27982
rect 57262 27970 57314 27982
rect 39106 27918 39118 27970
rect 39170 27918 39182 27970
rect 41794 27918 41806 27970
rect 41858 27918 41870 27970
rect 55458 27918 55470 27970
rect 55522 27918 55534 27970
rect 56914 27918 56926 27970
rect 56978 27918 56990 27970
rect 39006 27906 39058 27918
rect 57262 27906 57314 27918
rect 57934 27970 57986 27982
rect 57934 27906 57986 27918
rect 8094 27858 8146 27870
rect 4834 27806 4846 27858
rect 4898 27806 4910 27858
rect 8094 27794 8146 27806
rect 9550 27858 9602 27870
rect 11342 27858 11394 27870
rect 10882 27806 10894 27858
rect 10946 27806 10958 27858
rect 9550 27794 9602 27806
rect 11342 27794 11394 27806
rect 12686 27858 12738 27870
rect 14478 27858 14530 27870
rect 12898 27806 12910 27858
rect 12962 27806 12974 27858
rect 12686 27794 12738 27806
rect 14478 27794 14530 27806
rect 14814 27858 14866 27870
rect 22878 27858 22930 27870
rect 28142 27858 28194 27870
rect 32510 27858 32562 27870
rect 18162 27806 18174 27858
rect 18226 27806 18238 27858
rect 19618 27806 19630 27858
rect 19682 27806 19694 27858
rect 25778 27806 25790 27858
rect 25842 27806 25854 27858
rect 31266 27806 31278 27858
rect 31330 27806 31342 27858
rect 31490 27806 31502 27858
rect 31554 27806 31566 27858
rect 14814 27794 14866 27806
rect 22878 27794 22930 27806
rect 28142 27794 28194 27806
rect 32510 27794 32562 27806
rect 35758 27858 35810 27870
rect 35758 27794 35810 27806
rect 38670 27858 38722 27870
rect 55134 27858 55186 27870
rect 41122 27806 41134 27858
rect 41186 27806 41198 27858
rect 51426 27806 51438 27858
rect 51490 27806 51502 27858
rect 38670 27794 38722 27806
rect 55134 27794 55186 27806
rect 57822 27858 57874 27870
rect 57822 27794 57874 27806
rect 12350 27746 12402 27758
rect 37774 27746 37826 27758
rect 7634 27694 7646 27746
rect 7698 27694 7710 27746
rect 9986 27694 9998 27746
rect 10050 27694 10062 27746
rect 22418 27694 22430 27746
rect 22482 27694 22494 27746
rect 26338 27694 26350 27746
rect 26402 27694 26414 27746
rect 31602 27694 31614 27746
rect 31666 27694 31678 27746
rect 34962 27694 34974 27746
rect 35026 27694 35038 27746
rect 39442 27694 39454 27746
rect 39506 27694 39518 27746
rect 43922 27694 43934 27746
rect 43986 27694 43998 27746
rect 52098 27694 52110 27746
rect 52162 27694 52174 27746
rect 54226 27694 54238 27746
rect 54290 27694 54302 27746
rect 12350 27682 12402 27694
rect 37774 27682 37826 27694
rect 14926 27634 14978 27646
rect 14926 27570 14978 27582
rect 57374 27634 57426 27646
rect 57374 27570 57426 27582
rect 57934 27634 57986 27646
rect 57934 27570 57986 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 24558 27298 24610 27310
rect 24558 27234 24610 27246
rect 26686 27298 26738 27310
rect 26686 27234 26738 27246
rect 9662 27186 9714 27198
rect 18174 27186 18226 27198
rect 12450 27134 12462 27186
rect 12514 27134 12526 27186
rect 9662 27122 9714 27134
rect 18174 27122 18226 27134
rect 18622 27186 18674 27198
rect 18622 27122 18674 27134
rect 19518 27186 19570 27198
rect 52782 27186 52834 27198
rect 31714 27134 31726 27186
rect 31778 27134 31790 27186
rect 33842 27134 33854 27186
rect 33906 27134 33918 27186
rect 41906 27134 41918 27186
rect 41970 27134 41982 27186
rect 58146 27134 58158 27186
rect 58210 27134 58222 27186
rect 19518 27122 19570 27134
rect 52782 27122 52834 27134
rect 12910 27074 12962 27086
rect 12910 27010 12962 27022
rect 14142 27074 14194 27086
rect 14142 27010 14194 27022
rect 14926 27074 14978 27086
rect 14926 27010 14978 27022
rect 26014 27074 26066 27086
rect 26014 27010 26066 27022
rect 26238 27074 26290 27086
rect 26238 27010 26290 27022
rect 30606 27074 30658 27086
rect 40014 27074 40066 27086
rect 52558 27074 52610 27086
rect 30930 27022 30942 27074
rect 30994 27022 31006 27074
rect 37986 27022 37998 27074
rect 38050 27022 38062 27074
rect 40898 27022 40910 27074
rect 40962 27022 40974 27074
rect 30606 27010 30658 27022
rect 40014 27010 40066 27022
rect 52558 27010 52610 27022
rect 53230 27074 53282 27086
rect 53230 27010 53282 27022
rect 53790 27074 53842 27086
rect 55346 27022 55358 27074
rect 55410 27022 55422 27074
rect 53790 27010 53842 27022
rect 13470 26962 13522 26974
rect 9202 26910 9214 26962
rect 9266 26910 9278 26962
rect 13470 26898 13522 26910
rect 13806 26962 13858 26974
rect 13806 26898 13858 26910
rect 14254 26962 14306 26974
rect 14254 26898 14306 26910
rect 24670 26962 24722 26974
rect 24670 26898 24722 26910
rect 25790 26962 25842 26974
rect 25790 26898 25842 26910
rect 26574 26962 26626 26974
rect 26574 26898 26626 26910
rect 29374 26962 29426 26974
rect 38670 26962 38722 26974
rect 38210 26910 38222 26962
rect 38274 26910 38286 26962
rect 29374 26898 29426 26910
rect 38670 26898 38722 26910
rect 44270 26962 44322 26974
rect 44270 26898 44322 26910
rect 44830 26962 44882 26974
rect 44830 26898 44882 26910
rect 45166 26962 45218 26974
rect 45166 26898 45218 26910
rect 45390 26962 45442 26974
rect 45390 26898 45442 26910
rect 53006 26962 53058 26974
rect 53006 26898 53058 26910
rect 53454 26962 53506 26974
rect 56018 26910 56030 26962
rect 56082 26910 56094 26962
rect 53454 26898 53506 26910
rect 8878 26850 8930 26862
rect 8878 26786 8930 26798
rect 14478 26850 14530 26862
rect 14478 26786 14530 26798
rect 14590 26850 14642 26862
rect 14590 26786 14642 26798
rect 14814 26850 14866 26862
rect 14814 26786 14866 26798
rect 24558 26850 24610 26862
rect 24558 26786 24610 26798
rect 25566 26850 25618 26862
rect 25566 26786 25618 26798
rect 25678 26850 25730 26862
rect 25678 26786 25730 26798
rect 26686 26850 26738 26862
rect 26686 26786 26738 26798
rect 28590 26850 28642 26862
rect 28590 26786 28642 26798
rect 29822 26850 29874 26862
rect 29822 26786 29874 26798
rect 43934 26850 43986 26862
rect 43934 26786 43986 26798
rect 44158 26850 44210 26862
rect 44158 26786 44210 26798
rect 44942 26850 44994 26862
rect 44942 26786 44994 26798
rect 53678 26850 53730 26862
rect 53678 26786 53730 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 9774 26514 9826 26526
rect 9774 26450 9826 26462
rect 10670 26514 10722 26526
rect 22318 26514 22370 26526
rect 16482 26462 16494 26514
rect 16546 26462 16558 26514
rect 10670 26450 10722 26462
rect 22318 26450 22370 26462
rect 22654 26514 22706 26526
rect 22654 26450 22706 26462
rect 25342 26514 25394 26526
rect 25342 26450 25394 26462
rect 26462 26514 26514 26526
rect 26462 26450 26514 26462
rect 27358 26514 27410 26526
rect 27358 26450 27410 26462
rect 28478 26514 28530 26526
rect 28478 26450 28530 26462
rect 29038 26514 29090 26526
rect 29038 26450 29090 26462
rect 30270 26514 30322 26526
rect 30270 26450 30322 26462
rect 30830 26514 30882 26526
rect 30830 26450 30882 26462
rect 34414 26514 34466 26526
rect 34414 26450 34466 26462
rect 39230 26514 39282 26526
rect 39230 26450 39282 26462
rect 52334 26514 52386 26526
rect 52334 26450 52386 26462
rect 57038 26514 57090 26526
rect 57038 26450 57090 26462
rect 15934 26402 15986 26414
rect 18174 26402 18226 26414
rect 15586 26350 15598 26402
rect 15650 26350 15662 26402
rect 17378 26350 17390 26402
rect 17442 26350 17454 26402
rect 15934 26338 15986 26350
rect 18174 26338 18226 26350
rect 18622 26402 18674 26414
rect 18622 26338 18674 26350
rect 25118 26402 25170 26414
rect 25118 26338 25170 26350
rect 25454 26402 25506 26414
rect 25454 26338 25506 26350
rect 28814 26402 28866 26414
rect 28814 26338 28866 26350
rect 29598 26402 29650 26414
rect 29598 26338 29650 26350
rect 33966 26402 34018 26414
rect 41470 26402 41522 26414
rect 39778 26350 39790 26402
rect 39842 26350 39854 26402
rect 33966 26338 34018 26350
rect 41470 26338 41522 26350
rect 52558 26402 52610 26414
rect 52558 26338 52610 26350
rect 52670 26402 52722 26414
rect 52670 26338 52722 26350
rect 9550 26290 9602 26302
rect 6066 26238 6078 26290
rect 6130 26238 6142 26290
rect 9550 26226 9602 26238
rect 10222 26290 10274 26302
rect 10222 26226 10274 26238
rect 11790 26290 11842 26302
rect 16830 26290 16882 26302
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 11790 26226 11842 26238
rect 16830 26226 16882 26238
rect 17726 26290 17778 26302
rect 17726 26226 17778 26238
rect 18062 26290 18114 26302
rect 18062 26226 18114 26238
rect 19182 26290 19234 26302
rect 26350 26290 26402 26302
rect 23762 26238 23774 26290
rect 23826 26238 23838 26290
rect 24210 26238 24222 26290
rect 24274 26238 24286 26290
rect 19182 26226 19234 26238
rect 26350 26226 26402 26238
rect 26574 26290 26626 26302
rect 26574 26226 26626 26238
rect 27134 26290 27186 26302
rect 28254 26290 28306 26302
rect 27458 26238 27470 26290
rect 27522 26238 27534 26290
rect 27134 26226 27186 26238
rect 28254 26226 28306 26238
rect 28590 26290 28642 26302
rect 28590 26226 28642 26238
rect 29150 26290 29202 26302
rect 29150 26226 29202 26238
rect 30158 26290 30210 26302
rect 40126 26290 40178 26302
rect 39442 26238 39454 26290
rect 39506 26238 39518 26290
rect 30158 26226 30210 26238
rect 40126 26226 40178 26238
rect 41134 26290 41186 26302
rect 48190 26290 48242 26302
rect 42578 26238 42590 26290
rect 42642 26238 42654 26290
rect 47618 26238 47630 26290
rect 47682 26238 47694 26290
rect 41134 26226 41186 26238
rect 48190 26226 48242 26238
rect 56590 26290 56642 26302
rect 56590 26226 56642 26238
rect 56926 26290 56978 26302
rect 56926 26226 56978 26238
rect 57262 26290 57314 26302
rect 57262 26226 57314 26238
rect 9662 26178 9714 26190
rect 6738 26126 6750 26178
rect 6802 26126 6814 26178
rect 8866 26126 8878 26178
rect 8930 26126 8942 26178
rect 9662 26114 9714 26126
rect 11006 26178 11058 26190
rect 23214 26178 23266 26190
rect 12226 26126 12238 26178
rect 12290 26126 12302 26178
rect 13906 26126 13918 26178
rect 13970 26126 13982 26178
rect 11006 26114 11058 26126
rect 23214 26114 23266 26126
rect 24334 26178 24386 26190
rect 24334 26114 24386 26126
rect 26126 26178 26178 26190
rect 26126 26114 26178 26126
rect 27246 26178 27298 26190
rect 27246 26114 27298 26126
rect 36766 26178 36818 26190
rect 36766 26114 36818 26126
rect 37662 26178 37714 26190
rect 37662 26114 37714 26126
rect 41918 26178 41970 26190
rect 58158 26178 58210 26190
rect 43250 26126 43262 26178
rect 43314 26126 43326 26178
rect 45378 26126 45390 26178
rect 45442 26126 45454 26178
rect 41918 26114 41970 26126
rect 58158 26114 58210 26126
rect 18174 26066 18226 26078
rect 18174 26002 18226 26014
rect 25902 26066 25954 26078
rect 25902 26002 25954 26014
rect 27806 26066 27858 26078
rect 27806 26002 27858 26014
rect 29486 26066 29538 26078
rect 29486 26002 29538 26014
rect 30270 26066 30322 26078
rect 30270 26002 30322 26014
rect 33854 26066 33906 26078
rect 33854 26002 33906 26014
rect 39118 26066 39170 26078
rect 39118 26002 39170 26014
rect 41022 26066 41074 26078
rect 41022 26002 41074 26014
rect 41358 26066 41410 26078
rect 41358 26002 41410 26014
rect 47294 26066 47346 26078
rect 47294 26002 47346 26014
rect 47630 26066 47682 26078
rect 47630 26002 47682 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 24670 25730 24722 25742
rect 24670 25666 24722 25678
rect 27694 25730 27746 25742
rect 27694 25666 27746 25678
rect 39790 25730 39842 25742
rect 39790 25666 39842 25678
rect 39902 25730 39954 25742
rect 39902 25666 39954 25678
rect 40686 25730 40738 25742
rect 40686 25666 40738 25678
rect 43598 25730 43650 25742
rect 43598 25666 43650 25678
rect 43934 25730 43986 25742
rect 43934 25666 43986 25678
rect 44046 25730 44098 25742
rect 44046 25666 44098 25678
rect 8318 25618 8370 25630
rect 8318 25554 8370 25566
rect 9438 25618 9490 25630
rect 9438 25554 9490 25566
rect 15486 25618 15538 25630
rect 15486 25554 15538 25566
rect 15934 25618 15986 25630
rect 15934 25554 15986 25566
rect 19742 25618 19794 25630
rect 19742 25554 19794 25566
rect 23326 25618 23378 25630
rect 23326 25554 23378 25566
rect 26126 25618 26178 25630
rect 26126 25554 26178 25566
rect 27806 25618 27858 25630
rect 27806 25554 27858 25566
rect 28590 25618 28642 25630
rect 28590 25554 28642 25566
rect 33854 25618 33906 25630
rect 33854 25554 33906 25566
rect 34190 25618 34242 25630
rect 34190 25554 34242 25566
rect 36206 25618 36258 25630
rect 36206 25554 36258 25566
rect 38334 25618 38386 25630
rect 38334 25554 38386 25566
rect 39006 25618 39058 25630
rect 39006 25554 39058 25566
rect 39342 25618 39394 25630
rect 46622 25618 46674 25630
rect 50318 25618 50370 25630
rect 45042 25566 45054 25618
rect 45106 25566 45118 25618
rect 46946 25566 46958 25618
rect 47010 25566 47022 25618
rect 49074 25566 49086 25618
rect 49138 25566 49150 25618
rect 39342 25554 39394 25566
rect 46622 25554 46674 25566
rect 50318 25554 50370 25566
rect 8542 25506 8594 25518
rect 8542 25442 8594 25454
rect 8766 25506 8818 25518
rect 12798 25506 12850 25518
rect 12226 25454 12238 25506
rect 12290 25454 12302 25506
rect 8766 25442 8818 25454
rect 12798 25442 12850 25454
rect 16270 25506 16322 25518
rect 21422 25506 21474 25518
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 16270 25442 16322 25454
rect 21422 25442 21474 25454
rect 23886 25506 23938 25518
rect 23886 25442 23938 25454
rect 24222 25506 24274 25518
rect 24222 25442 24274 25454
rect 25566 25506 25618 25518
rect 26014 25506 26066 25518
rect 32398 25506 32450 25518
rect 25890 25454 25902 25506
rect 25954 25454 25966 25506
rect 26898 25454 26910 25506
rect 26962 25454 26974 25506
rect 29138 25454 29150 25506
rect 29202 25454 29214 25506
rect 25566 25442 25618 25454
rect 26014 25442 26066 25454
rect 32398 25442 32450 25454
rect 32734 25506 32786 25518
rect 32734 25442 32786 25454
rect 33294 25506 33346 25518
rect 33294 25442 33346 25454
rect 34974 25506 35026 25518
rect 34974 25442 35026 25454
rect 36990 25506 37042 25518
rect 36990 25442 37042 25454
rect 37214 25506 37266 25518
rect 37214 25442 37266 25454
rect 37550 25506 37602 25518
rect 37550 25442 37602 25454
rect 38446 25506 38498 25518
rect 38446 25442 38498 25454
rect 40126 25506 40178 25518
rect 43710 25506 43762 25518
rect 41906 25454 41918 25506
rect 41970 25454 41982 25506
rect 40126 25442 40178 25454
rect 43710 25442 43762 25454
rect 45726 25506 45778 25518
rect 52558 25506 52610 25518
rect 45938 25454 45950 25506
rect 46002 25454 46014 25506
rect 49858 25454 49870 25506
rect 49922 25454 49934 25506
rect 45726 25442 45778 25454
rect 52558 25442 52610 25454
rect 53006 25506 53058 25518
rect 53006 25442 53058 25454
rect 53118 25506 53170 25518
rect 53118 25442 53170 25454
rect 53454 25506 53506 25518
rect 53454 25442 53506 25454
rect 53790 25506 53842 25518
rect 53790 25442 53842 25454
rect 8206 25394 8258 25406
rect 14030 25394 14082 25406
rect 11554 25342 11566 25394
rect 11618 25342 11630 25394
rect 8206 25330 8258 25342
rect 14030 25330 14082 25342
rect 14254 25394 14306 25406
rect 21758 25394 21810 25406
rect 14466 25342 14478 25394
rect 14530 25342 14542 25394
rect 17602 25342 17614 25394
rect 17666 25342 17678 25394
rect 14254 25330 14306 25342
rect 21758 25330 21810 25342
rect 21982 25394 22034 25406
rect 21982 25330 22034 25342
rect 24110 25394 24162 25406
rect 24110 25330 24162 25342
rect 24558 25394 24610 25406
rect 32622 25394 32674 25406
rect 26674 25342 26686 25394
rect 26738 25342 26750 25394
rect 27346 25342 27358 25394
rect 27410 25342 27422 25394
rect 29474 25342 29486 25394
rect 29538 25342 29550 25394
rect 30930 25342 30942 25394
rect 30994 25342 31006 25394
rect 24558 25330 24610 25342
rect 32622 25330 32674 25342
rect 32958 25394 33010 25406
rect 39230 25394 39282 25406
rect 34626 25342 34638 25394
rect 34690 25342 34702 25394
rect 35410 25342 35422 25394
rect 35474 25342 35486 25394
rect 32958 25330 33010 25342
rect 39230 25330 39282 25342
rect 40238 25394 40290 25406
rect 40238 25330 40290 25342
rect 40574 25394 40626 25406
rect 40574 25330 40626 25342
rect 40686 25394 40738 25406
rect 40686 25330 40738 25342
rect 41470 25394 41522 25406
rect 41470 25330 41522 25342
rect 44830 25394 44882 25406
rect 44830 25330 44882 25342
rect 45054 25394 45106 25406
rect 45054 25330 45106 25342
rect 45278 25394 45330 25406
rect 45278 25330 45330 25342
rect 56590 25394 56642 25406
rect 56590 25330 56642 25342
rect 56702 25394 56754 25406
rect 56702 25330 56754 25342
rect 58158 25394 58210 25406
rect 58158 25330 58210 25342
rect 13918 25282 13970 25294
rect 13918 25218 13970 25230
rect 14142 25282 14194 25294
rect 14142 25218 14194 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 16606 25282 16658 25294
rect 16606 25218 16658 25230
rect 21534 25282 21586 25294
rect 21534 25218 21586 25230
rect 22542 25282 22594 25294
rect 22542 25218 22594 25230
rect 26238 25282 26290 25294
rect 31278 25282 31330 25294
rect 29698 25230 29710 25282
rect 29762 25230 29774 25282
rect 26238 25218 26290 25230
rect 31278 25218 31330 25230
rect 33182 25282 33234 25294
rect 33182 25218 33234 25230
rect 34078 25282 34130 25294
rect 34078 25218 34130 25230
rect 35758 25282 35810 25294
rect 35758 25218 35810 25230
rect 37102 25282 37154 25294
rect 37102 25218 37154 25230
rect 37998 25282 38050 25294
rect 37998 25218 38050 25230
rect 38222 25282 38274 25294
rect 42478 25282 42530 25294
rect 41682 25230 41694 25282
rect 41746 25230 41758 25282
rect 38222 25218 38274 25230
rect 42478 25218 42530 25230
rect 42926 25282 42978 25294
rect 42926 25218 42978 25230
rect 52782 25282 52834 25294
rect 52782 25218 52834 25230
rect 53678 25282 53730 25294
rect 53678 25218 53730 25230
rect 56366 25282 56418 25294
rect 56366 25218 56418 25230
rect 57598 25282 57650 25294
rect 57598 25218 57650 25230
rect 57822 25282 57874 25294
rect 57822 25218 57874 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 8990 24946 9042 24958
rect 8990 24882 9042 24894
rect 13358 24946 13410 24958
rect 13358 24882 13410 24894
rect 13918 24946 13970 24958
rect 13918 24882 13970 24894
rect 15150 24946 15202 24958
rect 15150 24882 15202 24894
rect 16046 24946 16098 24958
rect 16046 24882 16098 24894
rect 17390 24946 17442 24958
rect 17390 24882 17442 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 19070 24946 19122 24958
rect 19070 24882 19122 24894
rect 25566 24946 25618 24958
rect 25566 24882 25618 24894
rect 28142 24946 28194 24958
rect 28142 24882 28194 24894
rect 29934 24946 29986 24958
rect 29934 24882 29986 24894
rect 31390 24946 31442 24958
rect 31390 24882 31442 24894
rect 39230 24946 39282 24958
rect 39230 24882 39282 24894
rect 44382 24946 44434 24958
rect 44382 24882 44434 24894
rect 45838 24946 45890 24958
rect 45838 24882 45890 24894
rect 52558 24946 52610 24958
rect 56814 24946 56866 24958
rect 52558 24882 52610 24894
rect 53342 24890 53394 24902
rect 14142 24834 14194 24846
rect 16270 24834 16322 24846
rect 14466 24782 14478 24834
rect 14530 24782 14542 24834
rect 14142 24770 14194 24782
rect 16270 24770 16322 24782
rect 17614 24834 17666 24846
rect 17614 24770 17666 24782
rect 18622 24834 18674 24846
rect 25342 24834 25394 24846
rect 20514 24782 20526 24834
rect 20578 24782 20590 24834
rect 18622 24770 18674 24782
rect 25342 24770 25394 24782
rect 27694 24834 27746 24846
rect 27694 24770 27746 24782
rect 28926 24834 28978 24846
rect 40910 24834 40962 24846
rect 36082 24782 36094 24834
rect 36146 24782 36158 24834
rect 28926 24770 28978 24782
rect 40910 24770 40962 24782
rect 41134 24834 41186 24846
rect 41134 24770 41186 24782
rect 42142 24834 42194 24846
rect 52782 24834 52834 24846
rect 50194 24782 50206 24834
rect 50258 24782 50270 24834
rect 42142 24770 42194 24782
rect 52782 24770 52834 24782
rect 52894 24834 52946 24846
rect 56814 24882 56866 24894
rect 53342 24826 53394 24838
rect 53454 24834 53506 24846
rect 52894 24770 52946 24782
rect 53454 24770 53506 24782
rect 57822 24834 57874 24846
rect 57822 24770 57874 24782
rect 25230 24722 25282 24734
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 14354 24670 14366 24722
rect 14418 24670 14430 24722
rect 16482 24670 16494 24722
rect 16546 24670 16558 24722
rect 16706 24670 16718 24722
rect 16770 24670 16782 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 19730 24670 19742 24722
rect 19794 24670 19806 24722
rect 23426 24670 23438 24722
rect 23490 24670 23502 24722
rect 25230 24658 25282 24670
rect 27470 24722 27522 24734
rect 27470 24658 27522 24670
rect 28702 24722 28754 24734
rect 32958 24722 33010 24734
rect 29138 24670 29150 24722
rect 29202 24670 29214 24722
rect 29474 24670 29486 24722
rect 29538 24670 29550 24722
rect 28702 24658 28754 24670
rect 32958 24658 33010 24670
rect 33294 24722 33346 24734
rect 42702 24722 42754 24734
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 34178 24670 34190 24722
rect 34242 24670 34254 24722
rect 35410 24670 35422 24722
rect 35474 24670 35486 24722
rect 33294 24658 33346 24670
rect 42702 24658 42754 24670
rect 43038 24722 43090 24734
rect 56478 24722 56530 24734
rect 49522 24670 49534 24722
rect 49586 24670 49598 24722
rect 43038 24658 43090 24670
rect 56478 24658 56530 24670
rect 56926 24722 56978 24734
rect 56926 24658 56978 24670
rect 57150 24722 57202 24734
rect 57150 24658 57202 24670
rect 14030 24610 14082 24622
rect 10770 24558 10782 24610
rect 10834 24558 10846 24610
rect 12898 24558 12910 24610
rect 12962 24558 12974 24610
rect 14030 24546 14082 24558
rect 15598 24610 15650 24622
rect 15598 24546 15650 24558
rect 16158 24610 16210 24622
rect 22990 24610 23042 24622
rect 22642 24558 22654 24610
rect 22706 24558 22718 24610
rect 16158 24546 16210 24558
rect 22990 24546 23042 24558
rect 23998 24610 24050 24622
rect 38670 24610 38722 24622
rect 29026 24558 29038 24610
rect 29090 24558 29102 24610
rect 31826 24558 31838 24610
rect 31890 24558 31902 24610
rect 38210 24558 38222 24610
rect 38274 24558 38286 24610
rect 23998 24546 24050 24558
rect 38670 24546 38722 24558
rect 41022 24610 41074 24622
rect 41022 24546 41074 24558
rect 41806 24610 41858 24622
rect 44830 24610 44882 24622
rect 43474 24558 43486 24610
rect 43538 24558 43550 24610
rect 41806 24546 41858 24558
rect 44830 24546 44882 24558
rect 45278 24610 45330 24622
rect 53902 24610 53954 24622
rect 52322 24558 52334 24610
rect 52386 24558 52398 24610
rect 57474 24558 57486 24610
rect 57538 24558 57550 24610
rect 45278 24546 45330 24558
rect 53902 24546 53954 24558
rect 27134 24498 27186 24510
rect 27134 24434 27186 24446
rect 53342 24498 53394 24510
rect 53342 24434 53394 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 31502 24162 31554 24174
rect 31502 24098 31554 24110
rect 17838 24050 17890 24062
rect 17838 23986 17890 23998
rect 19406 24050 19458 24062
rect 19406 23986 19458 23998
rect 22318 24050 22370 24062
rect 22318 23986 22370 23998
rect 27694 24050 27746 24062
rect 27694 23986 27746 23998
rect 29150 24050 29202 24062
rect 29150 23986 29202 23998
rect 38446 24050 38498 24062
rect 38446 23986 38498 23998
rect 45166 24050 45218 24062
rect 55122 23998 55134 24050
rect 55186 23998 55198 24050
rect 57250 23998 57262 24050
rect 57314 23998 57326 24050
rect 45166 23986 45218 23998
rect 20302 23938 20354 23950
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 19842 23886 19854 23938
rect 19906 23886 19918 23938
rect 20302 23874 20354 23886
rect 22206 23938 22258 23950
rect 27918 23938 27970 23950
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 26898 23886 26910 23938
rect 26962 23886 26974 23938
rect 22206 23874 22258 23886
rect 27918 23874 27970 23886
rect 33742 23938 33794 23950
rect 45502 23938 45554 23950
rect 35746 23886 35758 23938
rect 35810 23886 35822 23938
rect 33742 23874 33794 23886
rect 45502 23874 45554 23886
rect 46062 23938 46114 23950
rect 46062 23874 46114 23886
rect 52782 23938 52834 23950
rect 52782 23874 52834 23886
rect 53006 23938 53058 23950
rect 53006 23874 53058 23886
rect 53342 23938 53394 23950
rect 53342 23874 53394 23886
rect 53790 23938 53842 23950
rect 58034 23886 58046 23938
rect 58098 23886 58110 23938
rect 53790 23874 53842 23886
rect 17278 23826 17330 23838
rect 17278 23762 17330 23774
rect 24334 23826 24386 23838
rect 24334 23762 24386 23774
rect 26350 23826 26402 23838
rect 31614 23826 31666 23838
rect 28242 23774 28254 23826
rect 28306 23774 28318 23826
rect 26350 23762 26402 23774
rect 31614 23762 31666 23774
rect 32062 23826 32114 23838
rect 35970 23774 35982 23826
rect 36034 23774 36046 23826
rect 32062 23762 32114 23774
rect 20750 23714 20802 23726
rect 20750 23650 20802 23662
rect 21982 23714 22034 23726
rect 21982 23650 22034 23662
rect 22430 23714 22482 23726
rect 22430 23650 22482 23662
rect 22654 23714 22706 23726
rect 29262 23714 29314 23726
rect 46510 23714 46562 23726
rect 26786 23662 26798 23714
rect 26850 23662 26862 23714
rect 33394 23662 33406 23714
rect 33458 23662 33470 23714
rect 45826 23662 45838 23714
rect 45890 23662 45902 23714
rect 22654 23650 22706 23662
rect 29262 23650 29314 23662
rect 46510 23650 46562 23662
rect 46622 23714 46674 23726
rect 46622 23650 46674 23662
rect 46734 23714 46786 23726
rect 46734 23650 46786 23662
rect 53006 23714 53058 23726
rect 53006 23650 53058 23662
rect 53454 23714 53506 23726
rect 53454 23650 53506 23662
rect 53678 23714 53730 23726
rect 53678 23650 53730 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 23438 23378 23490 23390
rect 23438 23314 23490 23326
rect 25342 23378 25394 23390
rect 25342 23314 25394 23326
rect 25566 23378 25618 23390
rect 25566 23314 25618 23326
rect 25790 23378 25842 23390
rect 25790 23314 25842 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 33630 23378 33682 23390
rect 33630 23314 33682 23326
rect 34078 23378 34130 23390
rect 34078 23314 34130 23326
rect 41022 23378 41074 23390
rect 41022 23314 41074 23326
rect 41806 23378 41858 23390
rect 41806 23314 41858 23326
rect 42030 23378 42082 23390
rect 42030 23314 42082 23326
rect 42478 23378 42530 23390
rect 42478 23314 42530 23326
rect 43374 23378 43426 23390
rect 43374 23314 43426 23326
rect 44158 23378 44210 23390
rect 44158 23314 44210 23326
rect 44606 23378 44658 23390
rect 44606 23314 44658 23326
rect 56702 23378 56754 23390
rect 56702 23314 56754 23326
rect 56926 23378 56978 23390
rect 56926 23314 56978 23326
rect 22766 23266 22818 23278
rect 16034 23214 16046 23266
rect 16098 23214 16110 23266
rect 22766 23202 22818 23214
rect 24334 23266 24386 23278
rect 24334 23202 24386 23214
rect 25230 23266 25282 23278
rect 39230 23266 39282 23278
rect 54126 23266 54178 23278
rect 30034 23214 30046 23266
rect 30098 23214 30110 23266
rect 44930 23214 44942 23266
rect 44994 23214 45006 23266
rect 51426 23214 51438 23266
rect 51490 23214 51502 23266
rect 25230 23202 25282 23214
rect 39230 23202 39282 23214
rect 54126 23202 54178 23214
rect 54350 23266 54402 23278
rect 54350 23202 54402 23214
rect 56590 23266 56642 23278
rect 56590 23202 56642 23214
rect 17502 23154 17554 23166
rect 16818 23102 16830 23154
rect 16882 23102 16894 23154
rect 17502 23090 17554 23102
rect 22318 23154 22370 23166
rect 22318 23090 22370 23102
rect 22990 23154 23042 23166
rect 22990 23090 23042 23102
rect 23662 23154 23714 23166
rect 23662 23090 23714 23102
rect 24110 23154 24162 23166
rect 24110 23090 24162 23102
rect 24222 23154 24274 23166
rect 24222 23090 24274 23102
rect 25902 23154 25954 23166
rect 38110 23154 38162 23166
rect 30706 23102 30718 23154
rect 30770 23102 30782 23154
rect 25902 23090 25954 23102
rect 38110 23090 38162 23102
rect 38446 23154 38498 23166
rect 38446 23090 38498 23102
rect 38782 23154 38834 23166
rect 38782 23090 38834 23102
rect 42254 23154 42306 23166
rect 54014 23154 54066 23166
rect 45266 23102 45278 23154
rect 45330 23102 45342 23154
rect 50754 23102 50766 23154
rect 50818 23102 50830 23154
rect 42254 23090 42306 23102
rect 54014 23090 54066 23102
rect 19742 23042 19794 23054
rect 13906 22990 13918 23042
rect 13970 22990 13982 23042
rect 19742 22978 19794 22990
rect 22542 23042 22594 23054
rect 33070 23042 33122 23054
rect 27906 22990 27918 23042
rect 27970 22990 27982 23042
rect 22542 22978 22594 22990
rect 33070 22978 33122 22990
rect 38334 23042 38386 23054
rect 38334 22978 38386 22990
rect 42142 23042 42194 23054
rect 54686 23042 54738 23054
rect 43698 22990 43710 23042
rect 43762 22990 43774 23042
rect 46050 22990 46062 23042
rect 46114 22990 46126 23042
rect 48178 22990 48190 23042
rect 48242 22990 48254 23042
rect 53554 22990 53566 23042
rect 53618 22990 53630 23042
rect 42142 22978 42194 22990
rect 54686 22978 54738 22990
rect 58158 23042 58210 23054
rect 58158 22978 58210 22990
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 33182 22482 33234 22494
rect 45054 22482 45106 22494
rect 36418 22430 36430 22482
rect 36482 22430 36494 22482
rect 40674 22430 40686 22482
rect 40738 22430 40750 22482
rect 44146 22430 44158 22482
rect 44210 22430 44222 22482
rect 33182 22418 33234 22430
rect 45054 22418 45106 22430
rect 45502 22482 45554 22494
rect 45502 22418 45554 22430
rect 45838 22482 45890 22494
rect 51214 22482 51266 22494
rect 47506 22430 47518 22482
rect 47570 22430 47582 22482
rect 50754 22430 50766 22482
rect 50818 22430 50830 22482
rect 45838 22418 45890 22430
rect 51214 22418 51266 22430
rect 24446 22370 24498 22382
rect 24446 22306 24498 22318
rect 26462 22370 26514 22382
rect 26462 22306 26514 22318
rect 26910 22370 26962 22382
rect 45614 22370 45666 22382
rect 33506 22318 33518 22370
rect 33570 22318 33582 22370
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 38546 22318 38558 22370
rect 38610 22318 38622 22370
rect 41234 22318 41246 22370
rect 41298 22318 41310 22370
rect 26910 22306 26962 22318
rect 45614 22306 45666 22318
rect 45950 22370 46002 22382
rect 45950 22306 46002 22318
rect 46286 22370 46338 22382
rect 46286 22306 46338 22318
rect 46734 22370 46786 22382
rect 54910 22370 54962 22382
rect 47954 22318 47966 22370
rect 48018 22318 48030 22370
rect 46734 22306 46786 22318
rect 54910 22306 54962 22318
rect 56814 22370 56866 22382
rect 56814 22306 56866 22318
rect 57374 22370 57426 22382
rect 57374 22306 57426 22318
rect 57934 22370 57986 22382
rect 57934 22306 57986 22318
rect 23886 22258 23938 22270
rect 23886 22194 23938 22206
rect 25342 22258 25394 22270
rect 25342 22194 25394 22206
rect 27918 22258 27970 22270
rect 37214 22258 37266 22270
rect 34290 22206 34302 22258
rect 34354 22206 34366 22258
rect 27918 22194 27970 22206
rect 37214 22194 37266 22206
rect 37326 22258 37378 22270
rect 37326 22194 37378 22206
rect 37438 22258 37490 22270
rect 47070 22258 47122 22270
rect 54574 22258 54626 22270
rect 42018 22206 42030 22258
rect 42082 22206 42094 22258
rect 47170 22206 47182 22258
rect 47234 22206 47246 22258
rect 48626 22206 48638 22258
rect 48690 22206 48702 22258
rect 37438 22194 37490 22206
rect 47070 22194 47122 22206
rect 54574 22194 54626 22206
rect 55134 22258 55186 22270
rect 55134 22194 55186 22206
rect 56702 22258 56754 22270
rect 56702 22194 56754 22206
rect 57038 22258 57090 22270
rect 57038 22194 57090 22206
rect 46958 22146 47010 22158
rect 28466 22094 28478 22146
rect 28530 22094 28542 22146
rect 46958 22082 47010 22094
rect 54686 22146 54738 22158
rect 54686 22082 54738 22094
rect 56478 22146 56530 22158
rect 56478 22082 56530 22094
rect 57262 22146 57314 22158
rect 57262 22082 57314 22094
rect 57598 22146 57650 22158
rect 57598 22082 57650 22094
rect 57822 22146 57874 22158
rect 57822 22082 57874 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 18622 21810 18674 21822
rect 18622 21746 18674 21758
rect 19294 21810 19346 21822
rect 19294 21746 19346 21758
rect 19966 21810 20018 21822
rect 33630 21810 33682 21822
rect 25330 21758 25342 21810
rect 25394 21758 25406 21810
rect 19966 21746 20018 21758
rect 33630 21746 33682 21758
rect 34414 21810 34466 21822
rect 34414 21746 34466 21758
rect 35534 21810 35586 21822
rect 35534 21746 35586 21758
rect 36766 21810 36818 21822
rect 36766 21746 36818 21758
rect 40350 21810 40402 21822
rect 40350 21746 40402 21758
rect 41470 21810 41522 21822
rect 41470 21746 41522 21758
rect 46398 21810 46450 21822
rect 46398 21746 46450 21758
rect 47070 21810 47122 21822
rect 47070 21746 47122 21758
rect 47294 21810 47346 21822
rect 47294 21746 47346 21758
rect 49646 21810 49698 21822
rect 49646 21746 49698 21758
rect 26350 21698 26402 21710
rect 18274 21646 18286 21698
rect 18338 21646 18350 21698
rect 18946 21646 18958 21698
rect 19010 21646 19022 21698
rect 19618 21646 19630 21698
rect 19682 21646 19694 21698
rect 22418 21646 22430 21698
rect 22482 21646 22494 21698
rect 26350 21634 26402 21646
rect 27806 21698 27858 21710
rect 38110 21698 38162 21710
rect 33954 21646 33966 21698
rect 34018 21646 34030 21698
rect 36082 21646 36094 21698
rect 36146 21646 36158 21698
rect 37090 21646 37102 21698
rect 37154 21646 37166 21698
rect 27806 21634 27858 21646
rect 38110 21634 38162 21646
rect 41806 21698 41858 21710
rect 41806 21634 41858 21646
rect 49758 21698 49810 21710
rect 56926 21698 56978 21710
rect 54338 21646 54350 21698
rect 54402 21646 54414 21698
rect 49758 21634 49810 21646
rect 56926 21634 56978 21646
rect 57150 21698 57202 21710
rect 57150 21634 57202 21646
rect 34190 21586 34242 21598
rect 21746 21534 21758 21586
rect 21810 21534 21822 21586
rect 26786 21534 26798 21586
rect 26850 21534 26862 21586
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 34190 21522 34242 21534
rect 34526 21586 34578 21598
rect 34526 21522 34578 21534
rect 34862 21586 34914 21598
rect 34862 21522 34914 21534
rect 35086 21586 35138 21598
rect 35086 21522 35138 21534
rect 35646 21586 35698 21598
rect 35646 21522 35698 21534
rect 35758 21586 35810 21598
rect 38334 21586 38386 21598
rect 41134 21586 41186 21598
rect 36306 21534 36318 21586
rect 36370 21534 36382 21586
rect 38994 21534 39006 21586
rect 39058 21534 39070 21586
rect 35758 21522 35810 21534
rect 38334 21522 38386 21534
rect 41134 21522 41186 21534
rect 41470 21586 41522 21598
rect 41470 21522 41522 21534
rect 47406 21586 47458 21598
rect 55582 21586 55634 21598
rect 55122 21534 55134 21586
rect 55186 21534 55198 21586
rect 47406 21522 47458 21534
rect 55582 21522 55634 21534
rect 56478 21586 56530 21598
rect 56478 21522 56530 21534
rect 37774 21474 37826 21486
rect 24546 21422 24558 21474
rect 24610 21422 24622 21474
rect 37774 21410 37826 21422
rect 45390 21474 45442 21486
rect 45390 21410 45442 21422
rect 47854 21474 47906 21486
rect 56702 21474 56754 21486
rect 52210 21422 52222 21474
rect 52274 21422 52286 21474
rect 47854 21410 47906 21422
rect 56702 21410 56754 21422
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 14702 20914 14754 20926
rect 19294 20914 19346 20926
rect 17938 20862 17950 20914
rect 18002 20862 18014 20914
rect 14702 20850 14754 20862
rect 19294 20850 19346 20862
rect 24894 20914 24946 20926
rect 24894 20850 24946 20862
rect 30158 20914 30210 20926
rect 33506 20862 33518 20914
rect 33570 20862 33582 20914
rect 56018 20862 56030 20914
rect 56082 20862 56094 20914
rect 58146 20862 58158 20914
rect 58210 20862 58222 20914
rect 30158 20850 30210 20862
rect 18286 20802 18338 20814
rect 15026 20750 15038 20802
rect 15090 20750 15102 20802
rect 18286 20738 18338 20750
rect 18622 20802 18674 20814
rect 18622 20738 18674 20750
rect 18734 20802 18786 20814
rect 18734 20738 18786 20750
rect 20078 20802 20130 20814
rect 20078 20738 20130 20750
rect 20526 20802 20578 20814
rect 20526 20738 20578 20750
rect 22542 20802 22594 20814
rect 22542 20738 22594 20750
rect 22878 20802 22930 20814
rect 29038 20802 29090 20814
rect 28018 20750 28030 20802
rect 28082 20750 28094 20802
rect 22878 20738 22930 20750
rect 29038 20738 29090 20750
rect 29374 20802 29426 20814
rect 33966 20802 34018 20814
rect 30706 20750 30718 20802
rect 30770 20750 30782 20802
rect 55234 20750 55246 20802
rect 55298 20750 55310 20802
rect 29374 20738 29426 20750
rect 33966 20738 34018 20750
rect 18398 20690 18450 20702
rect 15810 20638 15822 20690
rect 15874 20638 15886 20690
rect 18398 20626 18450 20638
rect 20750 20690 20802 20702
rect 20750 20626 20802 20638
rect 21982 20690 22034 20702
rect 21982 20626 22034 20638
rect 29710 20690 29762 20702
rect 31378 20638 31390 20690
rect 31442 20638 31454 20690
rect 29710 20626 29762 20638
rect 20302 20578 20354 20590
rect 20302 20514 20354 20526
rect 21870 20578 21922 20590
rect 21870 20514 21922 20526
rect 22094 20578 22146 20590
rect 29262 20578 29314 20590
rect 28242 20526 28254 20578
rect 28306 20526 28318 20578
rect 22094 20514 22146 20526
rect 29262 20514 29314 20526
rect 41582 20578 41634 20590
rect 41582 20514 41634 20526
rect 47294 20578 47346 20590
rect 47294 20514 47346 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 18510 20242 18562 20254
rect 18510 20178 18562 20190
rect 31278 20242 31330 20254
rect 31278 20178 31330 20190
rect 58158 20242 58210 20254
rect 58158 20178 58210 20190
rect 18062 20130 18114 20142
rect 18062 20066 18114 20078
rect 18398 20130 18450 20142
rect 31614 20130 31666 20142
rect 20178 20078 20190 20130
rect 20242 20078 20254 20130
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 27458 20078 27470 20130
rect 27522 20078 27534 20130
rect 18398 20066 18450 20078
rect 31614 20066 31666 20078
rect 32062 20130 32114 20142
rect 32062 20066 32114 20078
rect 32398 20130 32450 20142
rect 32398 20066 32450 20078
rect 40350 20130 40402 20142
rect 40350 20066 40402 20078
rect 41246 20130 41298 20142
rect 41246 20066 41298 20078
rect 46622 20130 46674 20142
rect 46622 20066 46674 20078
rect 47966 20130 48018 20142
rect 47966 20066 48018 20078
rect 18622 20018 18674 20030
rect 31054 20018 31106 20030
rect 18946 19966 18958 20018
rect 19010 19966 19022 20018
rect 19394 19966 19406 20018
rect 19458 19966 19470 20018
rect 26562 19966 26574 20018
rect 26626 19966 26638 20018
rect 27234 19966 27246 20018
rect 27298 19966 27310 20018
rect 27906 19966 27918 20018
rect 27970 19966 27982 20018
rect 28578 19966 28590 20018
rect 28642 19966 28654 20018
rect 18622 19954 18674 19966
rect 31054 19954 31106 19966
rect 31390 20018 31442 20030
rect 31390 19954 31442 19966
rect 31950 20018 32002 20030
rect 31950 19954 32002 19966
rect 32174 20018 32226 20030
rect 32174 19954 32226 19966
rect 40910 20018 40962 20030
rect 40910 19954 40962 19966
rect 41470 20018 41522 20030
rect 46846 20018 46898 20030
rect 41794 19966 41806 20018
rect 41858 19966 41870 20018
rect 41470 19954 41522 19966
rect 46846 19954 46898 19966
rect 47070 20018 47122 20030
rect 47070 19954 47122 19966
rect 47518 20018 47570 20030
rect 47518 19954 47570 19966
rect 47742 20018 47794 20030
rect 47742 19954 47794 19966
rect 37774 19906 37826 19918
rect 22306 19854 22318 19906
rect 22370 19854 22382 19906
rect 30706 19854 30718 19906
rect 30770 19854 30782 19906
rect 37774 19842 37826 19854
rect 41022 19906 41074 19918
rect 46286 19906 46338 19918
rect 42578 19854 42590 19906
rect 42642 19854 42654 19906
rect 44706 19854 44718 19906
rect 44770 19854 44782 19906
rect 41022 19842 41074 19854
rect 46286 19842 46338 19854
rect 46734 19906 46786 19918
rect 46734 19842 46786 19854
rect 47630 19906 47682 19918
rect 47630 19842 47682 19854
rect 50318 19906 50370 19918
rect 50318 19842 50370 19854
rect 51214 19906 51266 19918
rect 51214 19842 51266 19854
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 17838 19346 17890 19358
rect 17266 19294 17278 19346
rect 17330 19294 17342 19346
rect 17838 19282 17890 19294
rect 26238 19346 26290 19358
rect 26238 19282 26290 19294
rect 30046 19346 30098 19358
rect 30046 19282 30098 19294
rect 39790 19346 39842 19358
rect 39790 19282 39842 19294
rect 42142 19346 42194 19358
rect 47842 19294 47854 19346
rect 47906 19294 47918 19346
rect 49970 19294 49982 19346
rect 50034 19294 50046 19346
rect 42142 19282 42194 19294
rect 18286 19234 18338 19246
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 18286 19170 18338 19182
rect 18958 19234 19010 19246
rect 18958 19170 19010 19182
rect 23662 19234 23714 19246
rect 23662 19170 23714 19182
rect 24334 19234 24386 19246
rect 24334 19170 24386 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 26798 19234 26850 19246
rect 26798 19170 26850 19182
rect 33742 19234 33794 19246
rect 33742 19170 33794 19182
rect 34302 19234 34354 19246
rect 34302 19170 34354 19182
rect 36990 19234 37042 19246
rect 36990 19170 37042 19182
rect 37214 19234 37266 19246
rect 37214 19170 37266 19182
rect 37550 19234 37602 19246
rect 37550 19170 37602 19182
rect 37998 19234 38050 19246
rect 37998 19170 38050 19182
rect 38782 19234 38834 19246
rect 38782 19170 38834 19182
rect 39118 19234 39170 19246
rect 39118 19170 39170 19182
rect 42254 19234 42306 19246
rect 42254 19170 42306 19182
rect 45614 19234 45666 19246
rect 45614 19170 45666 19182
rect 46174 19234 46226 19246
rect 50766 19234 50818 19246
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 46174 19170 46226 19182
rect 50766 19170 50818 19182
rect 50990 19234 51042 19246
rect 50990 19170 51042 19182
rect 27134 19122 27186 19134
rect 15138 19070 15150 19122
rect 15202 19070 15214 19122
rect 27134 19058 27186 19070
rect 35422 19122 35474 19134
rect 35422 19058 35474 19070
rect 39342 19122 39394 19134
rect 39342 19058 39394 19070
rect 45950 19122 46002 19134
rect 45950 19058 46002 19070
rect 50542 19122 50594 19134
rect 50542 19058 50594 19070
rect 51886 19122 51938 19134
rect 51886 19058 51938 19070
rect 18398 19010 18450 19022
rect 18398 18946 18450 18958
rect 18510 19010 18562 19022
rect 18510 18946 18562 18958
rect 23998 19010 24050 19022
rect 23998 18946 24050 18958
rect 26686 19010 26738 19022
rect 26686 18946 26738 18958
rect 29934 19010 29986 19022
rect 29934 18946 29986 18958
rect 30158 19010 30210 19022
rect 30158 18946 30210 18958
rect 30382 19010 30434 19022
rect 30382 18946 30434 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 34638 19010 34690 19022
rect 35982 19010 36034 19022
rect 34962 18958 34974 19010
rect 35026 18958 35038 19010
rect 34638 18946 34690 18958
rect 35982 18946 36034 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 37886 19010 37938 19022
rect 37886 18946 37938 18958
rect 38110 19010 38162 19022
rect 38110 18946 38162 18958
rect 38334 19010 38386 19022
rect 38334 18946 38386 18958
rect 38894 19010 38946 19022
rect 38894 18946 38946 18958
rect 41806 19010 41858 19022
rect 41806 18946 41858 18958
rect 42030 19010 42082 19022
rect 42030 18946 42082 18958
rect 45278 19010 45330 19022
rect 45278 18946 45330 18958
rect 45838 19010 45890 19022
rect 45838 18946 45890 18958
rect 50766 19010 50818 19022
rect 50766 18946 50818 18958
rect 51438 19010 51490 19022
rect 51438 18946 51490 18958
rect 51550 19010 51602 19022
rect 51550 18946 51602 18958
rect 51662 19010 51714 19022
rect 51662 18946 51714 18958
rect 52782 19010 52834 19022
rect 52782 18946 52834 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 21758 18674 21810 18686
rect 21758 18610 21810 18622
rect 28478 18674 28530 18686
rect 39566 18674 39618 18686
rect 33842 18622 33854 18674
rect 33906 18622 33918 18674
rect 28478 18610 28530 18622
rect 39566 18610 39618 18622
rect 39678 18674 39730 18686
rect 39678 18610 39730 18622
rect 41246 18674 41298 18686
rect 51314 18622 51326 18674
rect 51378 18622 51390 18674
rect 41246 18610 41298 18622
rect 18510 18562 18562 18574
rect 28702 18562 28754 18574
rect 24434 18510 24446 18562
rect 24498 18510 24510 18562
rect 26002 18510 26014 18562
rect 26066 18510 26078 18562
rect 18510 18498 18562 18510
rect 28702 18498 28754 18510
rect 39790 18562 39842 18574
rect 52670 18562 52722 18574
rect 45826 18510 45838 18562
rect 45890 18510 45902 18562
rect 50866 18510 50878 18562
rect 50930 18510 50942 18562
rect 39790 18498 39842 18510
rect 52670 18498 52722 18510
rect 17950 18450 18002 18462
rect 17950 18386 18002 18398
rect 18062 18450 18114 18462
rect 18062 18386 18114 18398
rect 18286 18450 18338 18462
rect 18286 18386 18338 18398
rect 19070 18450 19122 18462
rect 19070 18386 19122 18398
rect 21982 18450 22034 18462
rect 22990 18450 23042 18462
rect 22306 18398 22318 18450
rect 22370 18398 22382 18450
rect 21982 18386 22034 18398
rect 22990 18386 23042 18398
rect 23214 18450 23266 18462
rect 28590 18450 28642 18462
rect 34190 18450 34242 18462
rect 24210 18398 24222 18450
rect 24274 18398 24286 18450
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 29026 18398 29038 18450
rect 29090 18398 29102 18450
rect 33618 18398 33630 18450
rect 33682 18398 33694 18450
rect 23214 18386 23266 18398
rect 28590 18386 28642 18398
rect 34190 18386 34242 18398
rect 34750 18450 34802 18462
rect 40238 18450 40290 18462
rect 35298 18398 35310 18450
rect 35362 18398 35374 18450
rect 35970 18398 35982 18450
rect 36034 18398 36046 18450
rect 34750 18386 34802 18398
rect 40238 18386 40290 18398
rect 41358 18450 41410 18462
rect 41358 18386 41410 18398
rect 41470 18450 41522 18462
rect 42030 18450 42082 18462
rect 41794 18398 41806 18450
rect 41858 18398 41870 18450
rect 41470 18386 41522 18398
rect 42030 18386 42082 18398
rect 42366 18450 42418 18462
rect 42366 18386 42418 18398
rect 42590 18450 42642 18462
rect 42590 18386 42642 18398
rect 43150 18450 43202 18462
rect 43150 18386 43202 18398
rect 43934 18450 43986 18462
rect 43934 18386 43986 18398
rect 44494 18450 44546 18462
rect 52222 18450 52274 18462
rect 53118 18450 53170 18462
rect 45042 18398 45054 18450
rect 45106 18398 45118 18450
rect 50418 18398 50430 18450
rect 50482 18398 50494 18450
rect 51314 18398 51326 18450
rect 51378 18398 51390 18450
rect 52882 18398 52894 18450
rect 52946 18398 52958 18450
rect 44494 18386 44546 18398
rect 52222 18386 52274 18398
rect 53118 18386 53170 18398
rect 53790 18450 53842 18462
rect 53790 18386 53842 18398
rect 21870 18338 21922 18350
rect 23774 18338 23826 18350
rect 31390 18338 31442 18350
rect 38558 18338 38610 18350
rect 22306 18286 22318 18338
rect 22370 18335 22382 18338
rect 22754 18335 22766 18338
rect 22370 18289 22766 18335
rect 22370 18286 22382 18289
rect 22754 18286 22766 18289
rect 22818 18286 22830 18338
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 38098 18286 38110 18338
rect 38162 18286 38174 18338
rect 21870 18274 21922 18286
rect 23774 18274 23826 18286
rect 31390 18274 31442 18286
rect 38558 18274 38610 18286
rect 42254 18338 42306 18350
rect 42254 18274 42306 18286
rect 43598 18338 43650 18350
rect 53566 18338 53618 18350
rect 47954 18286 47966 18338
rect 48018 18286 48030 18338
rect 53218 18286 53230 18338
rect 53282 18286 53294 18338
rect 43598 18274 43650 18286
rect 53566 18274 53618 18286
rect 54462 18338 54514 18350
rect 54462 18274 54514 18286
rect 55134 18338 55186 18350
rect 55134 18274 55186 18286
rect 52334 18226 52386 18238
rect 54574 18226 54626 18238
rect 54114 18174 54126 18226
rect 54178 18174 54190 18226
rect 52334 18162 52386 18174
rect 54574 18162 54626 18174
rect 55246 18226 55298 18238
rect 55246 18162 55298 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 51550 17890 51602 17902
rect 52782 17890 52834 17902
rect 51874 17838 51886 17890
rect 51938 17838 51950 17890
rect 51550 17826 51602 17838
rect 52782 17826 52834 17838
rect 22318 17778 22370 17790
rect 47070 17778 47122 17790
rect 40674 17726 40686 17778
rect 40738 17726 40750 17778
rect 42130 17726 42142 17778
rect 42194 17726 42206 17778
rect 44258 17726 44270 17778
rect 44322 17726 44334 17778
rect 54338 17726 54350 17778
rect 54402 17726 54414 17778
rect 56466 17726 56478 17778
rect 56530 17726 56542 17778
rect 22318 17714 22370 17726
rect 47070 17714 47122 17726
rect 17390 17666 17442 17678
rect 17390 17602 17442 17614
rect 17950 17666 18002 17678
rect 17950 17602 18002 17614
rect 18398 17666 18450 17678
rect 18398 17602 18450 17614
rect 18958 17666 19010 17678
rect 18958 17602 19010 17614
rect 19182 17666 19234 17678
rect 19182 17602 19234 17614
rect 19854 17666 19906 17678
rect 19854 17602 19906 17614
rect 21198 17666 21250 17678
rect 21198 17602 21250 17614
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 23102 17666 23154 17678
rect 23102 17602 23154 17614
rect 30494 17666 30546 17678
rect 30494 17602 30546 17614
rect 30942 17666 30994 17678
rect 30942 17602 30994 17614
rect 31166 17666 31218 17678
rect 31166 17602 31218 17614
rect 31502 17666 31554 17678
rect 31502 17602 31554 17614
rect 31614 17666 31666 17678
rect 31614 17602 31666 17614
rect 32174 17666 32226 17678
rect 35534 17666 35586 17678
rect 44942 17666 44994 17678
rect 35074 17614 35086 17666
rect 35138 17614 35150 17666
rect 37762 17614 37774 17666
rect 37826 17614 37838 17666
rect 38546 17614 38558 17666
rect 38610 17614 38622 17666
rect 41458 17614 41470 17666
rect 41522 17614 41534 17666
rect 32174 17602 32226 17614
rect 35534 17602 35586 17614
rect 44942 17602 44994 17614
rect 46958 17666 47010 17678
rect 46958 17602 47010 17614
rect 47182 17666 47234 17678
rect 47182 17602 47234 17614
rect 50318 17666 50370 17678
rect 50318 17602 50370 17614
rect 50654 17666 50706 17678
rect 50654 17602 50706 17614
rect 50990 17666 51042 17678
rect 50990 17602 51042 17614
rect 52670 17666 52722 17678
rect 57138 17614 57150 17666
rect 57202 17614 57214 17666
rect 17726 17554 17778 17566
rect 51314 17558 51326 17610
rect 51378 17558 51390 17610
rect 52670 17602 52722 17614
rect 53330 17558 53342 17610
rect 53394 17558 53406 17610
rect 53566 17554 53618 17566
rect 58158 17554 58210 17566
rect 22754 17502 22766 17554
rect 22818 17502 22830 17554
rect 57810 17502 57822 17554
rect 57874 17502 57886 17554
rect 17726 17490 17778 17502
rect 53566 17490 53618 17502
rect 58158 17490 58210 17502
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 18286 17442 18338 17454
rect 18286 17378 18338 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 19294 17442 19346 17454
rect 19294 17378 19346 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 21422 17442 21474 17454
rect 21422 17378 21474 17390
rect 28366 17442 28418 17454
rect 28366 17378 28418 17390
rect 30718 17442 30770 17454
rect 30718 17378 30770 17390
rect 31726 17442 31778 17454
rect 31726 17378 31778 17390
rect 35982 17442 36034 17454
rect 35982 17378 36034 17390
rect 46622 17442 46674 17454
rect 46622 17378 46674 17390
rect 47406 17442 47458 17454
rect 47406 17378 47458 17390
rect 50654 17442 50706 17454
rect 50654 17378 50706 17390
rect 53118 17442 53170 17454
rect 53118 17378 53170 17390
rect 53454 17442 53506 17454
rect 53454 17378 53506 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 18286 17106 18338 17118
rect 18286 17042 18338 17054
rect 27582 17106 27634 17118
rect 27582 17042 27634 17054
rect 28030 17106 28082 17118
rect 28030 17042 28082 17054
rect 33182 17106 33234 17118
rect 33182 17042 33234 17054
rect 51214 17106 51266 17118
rect 51214 17042 51266 17054
rect 51662 17106 51714 17118
rect 51662 17042 51714 17054
rect 51886 17106 51938 17118
rect 51886 17042 51938 17054
rect 52110 17106 52162 17118
rect 52110 17042 52162 17054
rect 57486 17106 57538 17118
rect 57486 17042 57538 17054
rect 58270 17106 58322 17118
rect 58270 17042 58322 17054
rect 18622 16994 18674 17006
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 18622 16930 18674 16942
rect 18846 16994 18898 17006
rect 18846 16930 18898 16942
rect 19070 16994 19122 17006
rect 28142 16994 28194 17006
rect 20626 16942 20638 16994
rect 20690 16942 20702 16994
rect 19070 16930 19122 16942
rect 28142 16930 28194 16942
rect 28702 16994 28754 17006
rect 48974 16994 49026 17006
rect 30370 16942 30382 16994
rect 30434 16942 30446 16994
rect 28702 16930 28754 16942
rect 48974 16930 49026 16942
rect 17614 16882 17666 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 17614 16818 17666 16830
rect 18398 16882 18450 16894
rect 18398 16818 18450 16830
rect 19630 16882 19682 16894
rect 27694 16882 27746 16894
rect 19842 16830 19854 16882
rect 19906 16830 19918 16882
rect 19630 16818 19682 16830
rect 27694 16818 27746 16830
rect 28254 16882 28306 16894
rect 28254 16818 28306 16830
rect 28926 16882 28978 16894
rect 28926 16818 28978 16830
rect 29374 16882 29426 16894
rect 49310 16882 49362 16894
rect 29698 16830 29710 16882
rect 29762 16830 29774 16882
rect 29374 16818 29426 16830
rect 49310 16818 49362 16830
rect 52670 16882 52722 16894
rect 52670 16818 52722 16830
rect 52894 16882 52946 16894
rect 52894 16818 52946 16830
rect 53566 16882 53618 16894
rect 53566 16818 53618 16830
rect 28814 16770 28866 16782
rect 33630 16770 33682 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 22754 16718 22766 16770
rect 22818 16718 22830 16770
rect 32498 16718 32510 16770
rect 32562 16718 32574 16770
rect 28814 16706 28866 16718
rect 33630 16706 33682 16718
rect 41022 16770 41074 16782
rect 41022 16706 41074 16718
rect 41470 16770 41522 16782
rect 41470 16706 41522 16718
rect 51998 16770 52050 16782
rect 51998 16706 52050 16718
rect 53342 16770 53394 16782
rect 53342 16706 53394 16718
rect 53790 16770 53842 16782
rect 53790 16706 53842 16718
rect 54014 16770 54066 16782
rect 54014 16706 54066 16718
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 36082 16270 36094 16322
rect 36146 16319 36158 16322
rect 36418 16319 36430 16322
rect 36146 16273 36430 16319
rect 36146 16270 36158 16273
rect 36418 16270 36430 16273
rect 36482 16270 36494 16322
rect 37762 16270 37774 16322
rect 37826 16319 37838 16322
rect 38322 16319 38334 16322
rect 37826 16273 38334 16319
rect 37826 16270 37838 16273
rect 38322 16270 38334 16273
rect 38386 16270 38398 16322
rect 19742 16210 19794 16222
rect 16594 16158 16606 16210
rect 16658 16158 16670 16210
rect 18722 16158 18734 16210
rect 18786 16158 18798 16210
rect 19742 16146 19794 16158
rect 22430 16210 22482 16222
rect 36094 16210 36146 16222
rect 32162 16158 32174 16210
rect 32226 16158 32238 16210
rect 35634 16158 35646 16210
rect 35698 16158 35710 16210
rect 22430 16146 22482 16158
rect 36094 16146 36146 16158
rect 38334 16210 38386 16222
rect 38334 16146 38386 16158
rect 41470 16210 41522 16222
rect 54910 16210 54962 16222
rect 49298 16158 49310 16210
rect 49362 16158 49374 16210
rect 55234 16158 55246 16210
rect 55298 16158 55310 16210
rect 57362 16158 57374 16210
rect 57426 16158 57438 16210
rect 41470 16146 41522 16158
rect 54910 16146 54962 16158
rect 22766 16098 22818 16110
rect 15810 16046 15822 16098
rect 15874 16046 15886 16098
rect 22766 16034 22818 16046
rect 22990 16098 23042 16110
rect 22990 16034 23042 16046
rect 27694 16098 27746 16110
rect 27694 16034 27746 16046
rect 29262 16098 29314 16110
rect 29262 16034 29314 16046
rect 32510 16098 32562 16110
rect 32510 16034 32562 16046
rect 32734 16098 32786 16110
rect 32734 16034 32786 16046
rect 33630 16098 33682 16110
rect 33630 16034 33682 16046
rect 33966 16098 34018 16110
rect 33966 16034 34018 16046
rect 49534 16098 49586 16110
rect 51650 16046 51662 16098
rect 51714 16046 51726 16098
rect 58034 16046 58046 16098
rect 58098 16046 58110 16098
rect 49534 16034 49586 16046
rect 19294 15986 19346 15998
rect 19294 15922 19346 15934
rect 23326 15986 23378 15998
rect 23326 15922 23378 15934
rect 24446 15986 24498 15998
rect 24446 15922 24498 15934
rect 27470 15986 27522 15998
rect 27470 15922 27522 15934
rect 28142 15986 28194 15998
rect 28142 15922 28194 15934
rect 28366 15986 28418 15998
rect 28366 15922 28418 15934
rect 29374 15986 29426 15998
rect 29374 15922 29426 15934
rect 29710 15986 29762 15998
rect 29710 15922 29762 15934
rect 34302 15986 34354 15998
rect 34302 15922 34354 15934
rect 35310 15986 35362 15998
rect 35310 15922 35362 15934
rect 35534 15986 35586 15998
rect 50542 15986 50594 15998
rect 47842 15934 47854 15986
rect 47906 15934 47918 15986
rect 35534 15922 35586 15934
rect 50542 15922 50594 15934
rect 22990 15874 23042 15886
rect 22990 15810 23042 15822
rect 24558 15874 24610 15886
rect 24558 15810 24610 15822
rect 24670 15874 24722 15886
rect 24670 15810 24722 15822
rect 25230 15874 25282 15886
rect 25230 15810 25282 15822
rect 27918 15874 27970 15886
rect 27918 15810 27970 15822
rect 29486 15874 29538 15886
rect 29486 15810 29538 15822
rect 33182 15874 33234 15886
rect 33182 15810 33234 15822
rect 33966 15874 34018 15886
rect 33966 15810 34018 15822
rect 37998 15874 38050 15886
rect 45726 15874 45778 15886
rect 45378 15822 45390 15874
rect 45442 15822 45454 15874
rect 37998 15810 38050 15822
rect 45726 15810 45778 15822
rect 52110 15874 52162 15886
rect 52110 15810 52162 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 47742 15538 47794 15550
rect 21858 15486 21870 15538
rect 21922 15486 21934 15538
rect 38210 15486 38222 15538
rect 38274 15486 38286 15538
rect 47742 15474 47794 15486
rect 52110 15538 52162 15550
rect 52110 15474 52162 15486
rect 52334 15538 52386 15550
rect 52334 15474 52386 15486
rect 24222 15426 24274 15438
rect 34638 15426 34690 15438
rect 45054 15426 45106 15438
rect 27346 15374 27358 15426
rect 27410 15374 27422 15426
rect 35746 15374 35758 15426
rect 35810 15374 35822 15426
rect 39218 15374 39230 15426
rect 39282 15374 39294 15426
rect 24222 15362 24274 15374
rect 34638 15362 34690 15374
rect 45054 15362 45106 15374
rect 49086 15426 49138 15438
rect 49086 15362 49138 15374
rect 49422 15426 49474 15438
rect 49422 15362 49474 15374
rect 31502 15314 31554 15326
rect 38558 15314 38610 15326
rect 40910 15314 40962 15326
rect 23762 15262 23774 15314
rect 23826 15262 23838 15314
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 34066 15262 34078 15314
rect 34130 15262 34142 15314
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 39666 15262 39678 15314
rect 39730 15262 39742 15314
rect 40226 15262 40238 15314
rect 40290 15262 40302 15314
rect 31502 15250 31554 15262
rect 38558 15250 38610 15262
rect 40910 15250 40962 15262
rect 41134 15314 41186 15326
rect 45278 15314 45330 15326
rect 41906 15262 41918 15314
rect 41970 15262 41982 15314
rect 41134 15250 41186 15262
rect 45278 15250 45330 15262
rect 45614 15314 45666 15326
rect 45614 15250 45666 15262
rect 46846 15314 46898 15326
rect 46846 15250 46898 15262
rect 47294 15314 47346 15326
rect 47294 15250 47346 15262
rect 48974 15314 49026 15326
rect 48974 15250 49026 15262
rect 49982 15314 50034 15326
rect 49982 15250 50034 15262
rect 50318 15314 50370 15326
rect 50318 15250 50370 15262
rect 50654 15314 50706 15326
rect 50654 15250 50706 15262
rect 51662 15314 51714 15326
rect 51662 15250 51714 15262
rect 52558 15314 52610 15326
rect 52558 15250 52610 15262
rect 22430 15202 22482 15214
rect 29934 15202 29986 15214
rect 23650 15150 23662 15202
rect 23714 15150 23726 15202
rect 29474 15150 29486 15202
rect 29538 15150 29550 15202
rect 22430 15138 22482 15150
rect 29934 15138 29986 15150
rect 31726 15202 31778 15214
rect 38782 15202 38834 15214
rect 45166 15202 45218 15214
rect 33954 15150 33966 15202
rect 34018 15150 34030 15202
rect 37874 15150 37886 15202
rect 37938 15150 37950 15202
rect 39778 15150 39790 15202
rect 39842 15150 39854 15202
rect 42578 15150 42590 15202
rect 42642 15150 42654 15202
rect 44706 15150 44718 15202
rect 44770 15150 44782 15202
rect 31726 15138 31778 15150
rect 38782 15138 38834 15150
rect 45166 15138 45218 15150
rect 46622 15202 46674 15214
rect 46622 15138 46674 15150
rect 47070 15202 47122 15214
rect 47070 15138 47122 15150
rect 49310 15202 49362 15214
rect 49310 15138 49362 15150
rect 50206 15202 50258 15214
rect 50206 15138 50258 15150
rect 51438 15202 51490 15214
rect 51438 15138 51490 15150
rect 52446 15202 52498 15214
rect 52446 15138 52498 15150
rect 54126 15202 54178 15214
rect 54126 15138 54178 15150
rect 22206 15090 22258 15102
rect 54238 15090 54290 15102
rect 32050 15038 32062 15090
rect 32114 15038 32126 15090
rect 41458 15038 41470 15090
rect 41522 15038 41534 15090
rect 51090 15038 51102 15090
rect 51154 15038 51166 15090
rect 22206 15026 22258 15038
rect 54238 15026 54290 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 50542 14754 50594 14766
rect 50542 14690 50594 14702
rect 52670 14754 52722 14766
rect 52670 14690 52722 14702
rect 18286 14642 18338 14654
rect 18286 14578 18338 14590
rect 22654 14642 22706 14654
rect 27582 14642 27634 14654
rect 43710 14642 43762 14654
rect 24322 14590 24334 14642
rect 24386 14590 24398 14642
rect 26450 14590 26462 14642
rect 26514 14590 26526 14642
rect 38322 14590 38334 14642
rect 38386 14590 38398 14642
rect 41458 14590 41470 14642
rect 41522 14590 41534 14642
rect 22654 14578 22706 14590
rect 27582 14578 27634 14590
rect 43710 14578 43762 14590
rect 47854 14642 47906 14654
rect 47854 14578 47906 14590
rect 50766 14642 50818 14654
rect 50766 14578 50818 14590
rect 52782 14642 52834 14654
rect 57710 14642 57762 14654
rect 53666 14590 53678 14642
rect 53730 14590 53742 14642
rect 54338 14590 54350 14642
rect 54402 14590 54414 14642
rect 56466 14590 56478 14642
rect 56530 14590 56542 14642
rect 52782 14578 52834 14590
rect 57710 14578 57762 14590
rect 18510 14530 18562 14542
rect 26798 14530 26850 14542
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 18510 14466 18562 14478
rect 26798 14466 26850 14478
rect 37550 14530 37602 14542
rect 42590 14530 42642 14542
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 41682 14478 41694 14530
rect 41746 14478 41758 14530
rect 41906 14478 41918 14530
rect 41970 14478 41982 14530
rect 37550 14466 37602 14478
rect 42590 14466 42642 14478
rect 42814 14530 42866 14542
rect 42814 14466 42866 14478
rect 45054 14530 45106 14542
rect 45054 14466 45106 14478
rect 46734 14530 46786 14542
rect 46734 14466 46786 14478
rect 46846 14530 46898 14542
rect 46846 14466 46898 14478
rect 48078 14530 48130 14542
rect 51102 14530 51154 14542
rect 50194 14478 50206 14530
rect 50258 14478 50270 14530
rect 48078 14466 48130 14478
rect 51102 14466 51154 14478
rect 51214 14530 51266 14542
rect 53566 14530 53618 14542
rect 52098 14478 52110 14530
rect 52162 14478 52174 14530
rect 57250 14478 57262 14530
rect 57314 14478 57326 14530
rect 51214 14466 51266 14478
rect 53566 14466 53618 14478
rect 40910 14418 40962 14430
rect 39106 14366 39118 14418
rect 39170 14366 39182 14418
rect 39554 14366 39566 14418
rect 39618 14366 39630 14418
rect 40910 14354 40962 14366
rect 43038 14418 43090 14430
rect 43038 14354 43090 14366
rect 44718 14418 44770 14430
rect 44718 14354 44770 14366
rect 47182 14418 47234 14430
rect 51762 14366 51774 14418
rect 51826 14366 51838 14418
rect 53330 14366 53342 14418
rect 53394 14366 53406 14418
rect 47182 14354 47234 14366
rect 22094 14306 22146 14318
rect 18834 14254 18846 14306
rect 18898 14254 18910 14306
rect 22094 14242 22146 14254
rect 23214 14306 23266 14318
rect 33742 14306 33794 14318
rect 37886 14306 37938 14318
rect 42702 14306 42754 14318
rect 27122 14254 27134 14306
rect 27186 14254 27198 14306
rect 37202 14254 37214 14306
rect 37266 14254 37278 14306
rect 38994 14254 39006 14306
rect 39058 14254 39070 14306
rect 23214 14242 23266 14254
rect 33742 14242 33794 14254
rect 37886 14242 37938 14254
rect 42702 14242 42754 14254
rect 44942 14306 44994 14318
rect 44942 14242 44994 14254
rect 47070 14306 47122 14318
rect 51550 14306 51602 14318
rect 47506 14254 47518 14306
rect 47570 14254 47582 14306
rect 47070 14242 47122 14254
rect 51550 14242 51602 14254
rect 51886 14306 51938 14318
rect 51886 14242 51938 14254
rect 53118 14306 53170 14318
rect 53118 14242 53170 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 20750 13970 20802 13982
rect 20750 13906 20802 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 24334 13970 24386 13982
rect 24334 13906 24386 13918
rect 34190 13970 34242 13982
rect 34190 13906 34242 13918
rect 40014 13970 40066 13982
rect 40014 13906 40066 13918
rect 42478 13970 42530 13982
rect 42478 13906 42530 13918
rect 43262 13970 43314 13982
rect 43262 13906 43314 13918
rect 44158 13970 44210 13982
rect 44158 13906 44210 13918
rect 47630 13970 47682 13982
rect 47630 13906 47682 13918
rect 47854 13970 47906 13982
rect 47854 13906 47906 13918
rect 50654 13970 50706 13982
rect 50654 13906 50706 13918
rect 50766 13970 50818 13982
rect 50766 13906 50818 13918
rect 56702 13970 56754 13982
rect 56702 13906 56754 13918
rect 18734 13858 18786 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 18734 13794 18786 13806
rect 22654 13858 22706 13870
rect 34302 13858 34354 13870
rect 27906 13806 27918 13858
rect 27970 13806 27982 13858
rect 22654 13794 22706 13806
rect 34302 13794 34354 13806
rect 35310 13858 35362 13870
rect 35310 13794 35362 13806
rect 35758 13858 35810 13870
rect 35758 13794 35810 13806
rect 37550 13858 37602 13870
rect 37550 13794 37602 13806
rect 38446 13858 38498 13870
rect 38446 13794 38498 13806
rect 41470 13858 41522 13870
rect 41470 13794 41522 13806
rect 42814 13858 42866 13870
rect 42814 13794 42866 13806
rect 44046 13858 44098 13870
rect 44046 13794 44098 13806
rect 44942 13858 44994 13870
rect 44942 13794 44994 13806
rect 45166 13858 45218 13870
rect 45166 13794 45218 13806
rect 47406 13858 47458 13870
rect 47406 13794 47458 13806
rect 18286 13746 18338 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 18286 13682 18338 13694
rect 18846 13746 18898 13758
rect 18846 13682 18898 13694
rect 18958 13746 19010 13758
rect 20862 13746 20914 13758
rect 19842 13694 19854 13746
rect 19906 13694 19918 13746
rect 20178 13694 20190 13746
rect 20242 13694 20254 13746
rect 18958 13682 19010 13694
rect 20862 13682 20914 13694
rect 21086 13746 21138 13758
rect 21086 13682 21138 13694
rect 21310 13746 21362 13758
rect 21310 13682 21362 13694
rect 21422 13746 21474 13758
rect 22430 13746 22482 13758
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 21422 13682 21474 13694
rect 22430 13682 22482 13694
rect 22766 13746 22818 13758
rect 22766 13682 22818 13694
rect 22990 13746 23042 13758
rect 22990 13682 23042 13694
rect 23326 13746 23378 13758
rect 33854 13746 33906 13758
rect 23650 13694 23662 13746
rect 23714 13694 23726 13746
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 33058 13694 33070 13746
rect 33122 13694 33134 13746
rect 23326 13682 23378 13694
rect 33854 13682 33906 13694
rect 34526 13746 34578 13758
rect 34526 13682 34578 13694
rect 34750 13746 34802 13758
rect 39342 13746 39394 13758
rect 41918 13746 41970 13758
rect 35074 13694 35086 13746
rect 35138 13694 35150 13746
rect 39554 13694 39566 13746
rect 39618 13694 39630 13746
rect 41682 13694 41694 13746
rect 41746 13694 41758 13746
rect 34750 13682 34802 13694
rect 39342 13682 39394 13694
rect 41918 13682 41970 13694
rect 42366 13746 42418 13758
rect 42366 13682 42418 13694
rect 42702 13746 42754 13758
rect 42702 13682 42754 13694
rect 44382 13746 44434 13758
rect 44382 13682 44434 13694
rect 50206 13746 50258 13758
rect 50206 13682 50258 13694
rect 50878 13746 50930 13758
rect 50878 13682 50930 13694
rect 52670 13746 52722 13758
rect 56018 13694 56030 13746
rect 56082 13694 56094 13746
rect 52670 13682 52722 13694
rect 17502 13634 17554 13646
rect 22206 13634 22258 13646
rect 30494 13634 30546 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 19394 13582 19406 13634
rect 19458 13582 19470 13634
rect 23762 13582 23774 13634
rect 23826 13582 23838 13634
rect 30034 13582 30046 13634
rect 30098 13582 30110 13634
rect 17502 13570 17554 13582
rect 22206 13570 22258 13582
rect 30494 13570 30546 13582
rect 32062 13634 32114 13646
rect 32062 13570 32114 13582
rect 32398 13634 32450 13646
rect 32398 13570 32450 13582
rect 38110 13634 38162 13646
rect 38110 13570 38162 13582
rect 42142 13634 42194 13646
rect 42142 13570 42194 13582
rect 43710 13634 43762 13646
rect 47742 13634 47794 13646
rect 44930 13582 44942 13634
rect 44994 13582 45006 13634
rect 43710 13570 43762 13582
rect 47742 13570 47794 13582
rect 52782 13634 52834 13646
rect 53106 13582 53118 13634
rect 53170 13582 53182 13634
rect 55234 13582 55246 13634
rect 55298 13582 55310 13634
rect 52782 13570 52834 13582
rect 32510 13522 32562 13534
rect 20402 13470 20414 13522
rect 20466 13470 20478 13522
rect 21970 13470 21982 13522
rect 22034 13519 22046 13522
rect 22194 13519 22206 13522
rect 22034 13473 22206 13519
rect 22034 13470 22046 13473
rect 22194 13470 22206 13473
rect 22258 13470 22270 13522
rect 32510 13458 32562 13470
rect 33070 13522 33122 13534
rect 33070 13458 33122 13470
rect 33406 13522 33458 13534
rect 33406 13458 33458 13470
rect 34974 13522 35026 13534
rect 39006 13522 39058 13534
rect 37650 13470 37662 13522
rect 37714 13519 37726 13522
rect 38098 13519 38110 13522
rect 37714 13473 38110 13519
rect 37714 13470 37726 13473
rect 38098 13470 38110 13473
rect 38162 13470 38174 13522
rect 34974 13458 35026 13470
rect 39006 13458 39058 13470
rect 39118 13522 39170 13534
rect 39118 13458 39170 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 17838 13186 17890 13198
rect 17838 13122 17890 13134
rect 19966 13186 20018 13198
rect 19966 13122 20018 13134
rect 20526 13186 20578 13198
rect 20526 13122 20578 13134
rect 21310 13186 21362 13198
rect 21310 13122 21362 13134
rect 23550 13186 23602 13198
rect 23550 13122 23602 13134
rect 23774 13186 23826 13198
rect 23774 13122 23826 13134
rect 34638 13186 34690 13198
rect 34638 13122 34690 13134
rect 34750 13186 34802 13198
rect 34750 13122 34802 13134
rect 44830 13186 44882 13198
rect 44830 13122 44882 13134
rect 44942 13186 44994 13198
rect 44942 13122 44994 13134
rect 48190 13186 48242 13198
rect 48190 13122 48242 13134
rect 20414 13074 20466 13086
rect 19506 13022 19518 13074
rect 19570 13022 19582 13074
rect 20414 13010 20466 13022
rect 21422 13074 21474 13086
rect 34974 13074 35026 13086
rect 32386 13022 32398 13074
rect 32450 13022 32462 13074
rect 33618 13022 33630 13074
rect 33682 13022 33694 13074
rect 21422 13010 21474 13022
rect 34974 13010 35026 13022
rect 36430 13074 36482 13086
rect 36430 13010 36482 13022
rect 37102 13074 37154 13086
rect 42814 13074 42866 13086
rect 41010 13022 41022 13074
rect 41074 13022 41086 13074
rect 37102 13010 37154 13022
rect 42814 13010 42866 13022
rect 43374 13074 43426 13086
rect 43374 13010 43426 13022
rect 48078 13074 48130 13086
rect 48078 13010 48130 13022
rect 18398 12962 18450 12974
rect 18398 12898 18450 12910
rect 18622 12962 18674 12974
rect 18622 12898 18674 12910
rect 19854 12962 19906 12974
rect 22542 12962 22594 12974
rect 24222 12962 24274 12974
rect 21634 12910 21646 12962
rect 21698 12910 21710 12962
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 19854 12898 19906 12910
rect 22542 12898 22594 12910
rect 24222 12898 24274 12910
rect 24446 12962 24498 12974
rect 24446 12898 24498 12910
rect 24782 12962 24834 12974
rect 24782 12898 24834 12910
rect 25230 12962 25282 12974
rect 33518 12962 33570 12974
rect 29474 12910 29486 12962
rect 29538 12910 29550 12962
rect 33282 12910 33294 12962
rect 33346 12910 33358 12962
rect 25230 12898 25282 12910
rect 33518 12898 33570 12910
rect 35646 12962 35698 12974
rect 35646 12898 35698 12910
rect 38782 12962 38834 12974
rect 42366 12962 42418 12974
rect 39666 12910 39678 12962
rect 39730 12910 39742 12962
rect 38782 12898 38834 12910
rect 42366 12898 42418 12910
rect 43710 12962 43762 12974
rect 52894 12962 52946 12974
rect 45826 12910 45838 12962
rect 45890 12910 45902 12962
rect 47170 12910 47182 12962
rect 47234 12910 47246 12962
rect 43710 12898 43762 12910
rect 52894 12898 52946 12910
rect 17950 12850 18002 12862
rect 17950 12786 18002 12798
rect 18734 12850 18786 12862
rect 18734 12786 18786 12798
rect 18846 12850 18898 12862
rect 18846 12786 18898 12798
rect 19182 12850 19234 12862
rect 19182 12786 19234 12798
rect 22094 12850 22146 12862
rect 22094 12786 22146 12798
rect 22430 12850 22482 12862
rect 22430 12786 22482 12798
rect 22766 12850 22818 12862
rect 22766 12786 22818 12798
rect 22990 12850 23042 12862
rect 35422 12850 35474 12862
rect 30258 12798 30270 12850
rect 30322 12798 30334 12850
rect 22990 12786 23042 12798
rect 35422 12786 35474 12798
rect 35982 12850 36034 12862
rect 45278 12850 45330 12862
rect 47854 12850 47906 12862
rect 42018 12798 42030 12850
rect 42082 12798 42094 12850
rect 44034 12798 44046 12850
rect 44098 12798 44110 12850
rect 45490 12798 45502 12850
rect 45554 12798 45566 12850
rect 47506 12798 47518 12850
rect 47570 12798 47582 12850
rect 35982 12786 36034 12798
rect 45278 12786 45330 12798
rect 47854 12786 47906 12798
rect 17838 12738 17890 12750
rect 17838 12674 17890 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19966 12738 20018 12750
rect 19966 12674 20018 12686
rect 23438 12738 23490 12750
rect 23438 12674 23490 12686
rect 24334 12738 24386 12750
rect 24334 12674 24386 12686
rect 27470 12738 27522 12750
rect 34638 12738 34690 12750
rect 33954 12686 33966 12738
rect 34018 12686 34030 12738
rect 27470 12674 27522 12686
rect 34638 12674 34690 12686
rect 35646 12738 35698 12750
rect 35646 12674 35698 12686
rect 45614 12738 45666 12750
rect 45614 12674 45666 12686
rect 47406 12738 47458 12750
rect 47406 12674 47458 12686
rect 51102 12738 51154 12750
rect 51102 12674 51154 12686
rect 51438 12738 51490 12750
rect 51438 12674 51490 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 20862 12402 20914 12414
rect 20862 12338 20914 12350
rect 23326 12402 23378 12414
rect 23326 12338 23378 12350
rect 24222 12402 24274 12414
rect 24222 12338 24274 12350
rect 27022 12402 27074 12414
rect 27022 12338 27074 12350
rect 33070 12402 33122 12414
rect 33070 12338 33122 12350
rect 33518 12402 33570 12414
rect 33518 12338 33570 12350
rect 34526 12402 34578 12414
rect 34526 12338 34578 12350
rect 39006 12402 39058 12414
rect 39006 12338 39058 12350
rect 39902 12402 39954 12414
rect 39902 12338 39954 12350
rect 41134 12402 41186 12414
rect 41134 12338 41186 12350
rect 42590 12402 42642 12414
rect 42590 12338 42642 12350
rect 49758 12402 49810 12414
rect 49758 12338 49810 12350
rect 50654 12402 50706 12414
rect 52110 12402 52162 12414
rect 51650 12350 51662 12402
rect 51714 12350 51726 12402
rect 50654 12338 50706 12350
rect 52110 12338 52162 12350
rect 24558 12290 24610 12302
rect 24558 12226 24610 12238
rect 26686 12290 26738 12302
rect 26686 12226 26738 12238
rect 27694 12290 27746 12302
rect 40910 12290 40962 12302
rect 35970 12238 35982 12290
rect 36034 12238 36046 12290
rect 27694 12226 27746 12238
rect 40910 12226 40962 12238
rect 44718 12290 44770 12302
rect 44718 12226 44770 12238
rect 47742 12290 47794 12302
rect 52222 12290 52274 12302
rect 50978 12238 50990 12290
rect 51042 12238 51054 12290
rect 47742 12226 47794 12238
rect 52222 12226 52274 12238
rect 52670 12290 52722 12302
rect 52670 12226 52722 12238
rect 27022 12178 27074 12190
rect 18274 12126 18286 12178
rect 18338 12126 18350 12178
rect 27022 12114 27074 12126
rect 27246 12178 27298 12190
rect 27246 12114 27298 12126
rect 27470 12178 27522 12190
rect 27470 12114 27522 12126
rect 27806 12178 27858 12190
rect 33294 12178 33346 12190
rect 30146 12126 30158 12178
rect 30210 12126 30222 12178
rect 27806 12114 27858 12126
rect 33294 12114 33346 12126
rect 34302 12178 34354 12190
rect 34302 12114 34354 12126
rect 34638 12178 34690 12190
rect 34638 12114 34690 12126
rect 34750 12178 34802 12190
rect 38782 12178 38834 12190
rect 35298 12126 35310 12178
rect 35362 12126 35374 12178
rect 34750 12114 34802 12126
rect 38782 12114 38834 12126
rect 39118 12178 39170 12190
rect 39118 12114 39170 12126
rect 39230 12178 39282 12190
rect 39230 12114 39282 12126
rect 39566 12178 39618 12190
rect 39566 12114 39618 12126
rect 39902 12178 39954 12190
rect 39902 12114 39954 12126
rect 40238 12178 40290 12190
rect 40238 12114 40290 12126
rect 50318 12178 50370 12190
rect 50318 12114 50370 12126
rect 51326 12178 51378 12190
rect 51326 12114 51378 12126
rect 51886 12178 51938 12190
rect 53218 12126 53230 12178
rect 53282 12126 53294 12178
rect 51886 12114 51938 12126
rect 21198 12066 21250 12078
rect 18834 12014 18846 12066
rect 18898 12014 18910 12066
rect 21198 12002 21250 12014
rect 28254 12066 28306 12078
rect 33182 12066 33234 12078
rect 41694 12066 41746 12078
rect 30930 12014 30942 12066
rect 30994 12014 31006 12066
rect 38098 12014 38110 12066
rect 38162 12014 38174 12066
rect 41234 12014 41246 12066
rect 41298 12014 41310 12066
rect 28254 12002 28306 12014
rect 33182 12002 33234 12014
rect 41694 12002 41746 12014
rect 42142 12066 42194 12078
rect 55346 12014 55358 12066
rect 55410 12014 55422 12066
rect 42142 12002 42194 12014
rect 44606 11954 44658 11966
rect 44606 11890 44658 11902
rect 47854 11954 47906 11966
rect 47854 11890 47906 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 19518 11618 19570 11630
rect 19518 11554 19570 11566
rect 19630 11618 19682 11630
rect 57262 11618 57314 11630
rect 32722 11566 32734 11618
rect 32786 11615 32798 11618
rect 33170 11615 33182 11618
rect 32786 11569 33182 11615
rect 32786 11566 32798 11569
rect 33170 11566 33182 11569
rect 33234 11566 33246 11618
rect 19630 11554 19682 11566
rect 57262 11554 57314 11566
rect 29262 11506 29314 11518
rect 17266 11454 17278 11506
rect 17330 11454 17342 11506
rect 24658 11454 24670 11506
rect 24722 11454 24734 11506
rect 26786 11454 26798 11506
rect 26850 11454 26862 11506
rect 29262 11442 29314 11454
rect 29710 11506 29762 11518
rect 29710 11442 29762 11454
rect 31838 11506 31890 11518
rect 31838 11442 31890 11454
rect 33070 11506 33122 11518
rect 33070 11442 33122 11454
rect 33518 11506 33570 11518
rect 33518 11442 33570 11454
rect 35086 11506 35138 11518
rect 35086 11442 35138 11454
rect 37886 11506 37938 11518
rect 37886 11442 37938 11454
rect 38334 11506 38386 11518
rect 42366 11506 42418 11518
rect 40226 11454 40238 11506
rect 40290 11454 40302 11506
rect 38334 11442 38386 11454
rect 42366 11442 42418 11454
rect 43038 11506 43090 11518
rect 50094 11506 50146 11518
rect 46722 11454 46734 11506
rect 46786 11454 46798 11506
rect 48850 11454 48862 11506
rect 48914 11454 48926 11506
rect 43038 11442 43090 11454
rect 50094 11442 50146 11454
rect 50654 11506 50706 11518
rect 56030 11506 56082 11518
rect 52658 11454 52670 11506
rect 52722 11454 52734 11506
rect 50654 11442 50706 11454
rect 56030 11442 56082 11454
rect 24334 11394 24386 11406
rect 28254 11394 28306 11406
rect 14354 11342 14366 11394
rect 14418 11342 14430 11394
rect 21522 11342 21534 11394
rect 21586 11342 21598 11394
rect 27458 11342 27470 11394
rect 27522 11342 27534 11394
rect 24334 11330 24386 11342
rect 28254 11330 28306 11342
rect 31614 11394 31666 11406
rect 31614 11330 31666 11342
rect 32062 11394 32114 11406
rect 32622 11394 32674 11406
rect 32274 11342 32286 11394
rect 32338 11342 32350 11394
rect 32062 11330 32114 11342
rect 32622 11330 32674 11342
rect 38670 11394 38722 11406
rect 50990 11394 51042 11406
rect 39442 11342 39454 11394
rect 39506 11342 39518 11394
rect 49634 11342 49646 11394
rect 49698 11342 49710 11394
rect 38670 11330 38722 11342
rect 50990 11330 51042 11342
rect 51886 11394 51938 11406
rect 51886 11330 51938 11342
rect 52110 11394 52162 11406
rect 55570 11342 55582 11394
rect 55634 11342 55646 11394
rect 52110 11330 52162 11342
rect 18734 11282 18786 11294
rect 21310 11282 21362 11294
rect 15138 11230 15150 11282
rect 15202 11230 15214 11282
rect 18946 11230 18958 11282
rect 19010 11230 19022 11282
rect 18734 11218 18786 11230
rect 21310 11218 21362 11230
rect 33966 11282 34018 11294
rect 33966 11218 34018 11230
rect 51326 11282 51378 11294
rect 51326 11218 51378 11230
rect 51550 11282 51602 11294
rect 57374 11282 57426 11294
rect 54786 11230 54798 11282
rect 54850 11230 54862 11282
rect 51550 11218 51602 11230
rect 57374 11218 57426 11230
rect 57822 11282 57874 11294
rect 57822 11218 57874 11230
rect 58158 11282 58210 11294
rect 58158 11218 58210 11230
rect 17726 11170 17778 11182
rect 17726 11106 17778 11118
rect 18846 11170 18898 11182
rect 18846 11106 18898 11118
rect 19182 11170 19234 11182
rect 19182 11106 19234 11118
rect 20190 11170 20242 11182
rect 30606 11170 30658 11182
rect 23986 11118 23998 11170
rect 24050 11118 24062 11170
rect 27906 11118 27918 11170
rect 27970 11118 27982 11170
rect 20190 11106 20242 11118
rect 30606 11106 30658 11118
rect 31502 11170 31554 11182
rect 31502 11106 31554 11118
rect 39006 11170 39058 11182
rect 39006 11106 39058 11118
rect 51102 11170 51154 11182
rect 51102 11106 51154 11118
rect 51774 11170 51826 11182
rect 51774 11106 51826 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 15822 10834 15874 10846
rect 15822 10770 15874 10782
rect 18174 10834 18226 10846
rect 18174 10770 18226 10782
rect 26686 10834 26738 10846
rect 26686 10770 26738 10782
rect 27246 10834 27298 10846
rect 27246 10770 27298 10782
rect 31166 10834 31218 10846
rect 31166 10770 31218 10782
rect 31726 10834 31778 10846
rect 31726 10770 31778 10782
rect 41694 10834 41746 10846
rect 41694 10770 41746 10782
rect 42814 10834 42866 10846
rect 51998 10834 52050 10846
rect 47170 10782 47182 10834
rect 47234 10782 47246 10834
rect 42814 10770 42866 10782
rect 51998 10770 52050 10782
rect 15934 10722 15986 10734
rect 15934 10658 15986 10670
rect 18062 10722 18114 10734
rect 18062 10658 18114 10670
rect 18398 10722 18450 10734
rect 18398 10658 18450 10670
rect 18734 10722 18786 10734
rect 27022 10722 27074 10734
rect 51326 10722 51378 10734
rect 23762 10670 23774 10722
rect 23826 10670 23838 10722
rect 43922 10670 43934 10722
rect 43986 10670 43998 10722
rect 50194 10670 50206 10722
rect 50258 10670 50270 10722
rect 18734 10658 18786 10670
rect 27022 10658 27074 10670
rect 51326 10658 51378 10670
rect 51438 10722 51490 10734
rect 51438 10658 51490 10670
rect 17838 10610 17890 10622
rect 25342 10610 25394 10622
rect 24546 10558 24558 10610
rect 24610 10558 24622 10610
rect 17838 10546 17890 10558
rect 25342 10546 25394 10558
rect 26910 10610 26962 10622
rect 30942 10610 30994 10622
rect 30258 10558 30270 10610
rect 30322 10558 30334 10610
rect 26910 10546 26962 10558
rect 30942 10546 30994 10558
rect 31278 10610 31330 10622
rect 31278 10546 31330 10558
rect 42254 10610 42306 10622
rect 46846 10610 46898 10622
rect 43138 10558 43150 10610
rect 43202 10558 43214 10610
rect 42254 10546 42306 10558
rect 46846 10546 46898 10558
rect 49870 10610 49922 10622
rect 49870 10546 49922 10558
rect 51662 10610 51714 10622
rect 51662 10546 51714 10558
rect 58158 10610 58210 10622
rect 58158 10546 58210 10558
rect 49534 10498 49586 10510
rect 21634 10446 21646 10498
rect 21698 10446 21710 10498
rect 27458 10446 27470 10498
rect 27522 10446 27534 10498
rect 29586 10446 29598 10498
rect 29650 10446 29662 10498
rect 46050 10446 46062 10498
rect 46114 10446 46126 10498
rect 49534 10434 49586 10446
rect 50654 10498 50706 10510
rect 50654 10434 50706 10446
rect 18958 10386 19010 10398
rect 18958 10322 19010 10334
rect 19182 10386 19234 10398
rect 19182 10322 19234 10334
rect 19406 10386 19458 10398
rect 19406 10322 19458 10334
rect 19854 10386 19906 10398
rect 19854 10322 19906 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 17950 10050 18002 10062
rect 17950 9986 18002 9998
rect 15934 9938 15986 9950
rect 19966 9938 20018 9950
rect 17602 9886 17614 9938
rect 17666 9886 17678 9938
rect 18610 9886 18622 9938
rect 18674 9886 18686 9938
rect 15934 9874 15986 9886
rect 19966 9874 20018 9886
rect 22206 9938 22258 9950
rect 30494 9938 30546 9950
rect 26674 9886 26686 9938
rect 26738 9886 26750 9938
rect 22206 9874 22258 9886
rect 30494 9874 30546 9886
rect 32286 9938 32338 9950
rect 32286 9874 32338 9886
rect 35422 9938 35474 9950
rect 35422 9874 35474 9886
rect 42590 9938 42642 9950
rect 42590 9874 42642 9886
rect 43486 9938 43538 9950
rect 43486 9874 43538 9886
rect 52110 9938 52162 9950
rect 52110 9874 52162 9886
rect 18174 9826 18226 9838
rect 19406 9826 19458 9838
rect 18834 9774 18846 9826
rect 18898 9774 18910 9826
rect 18174 9762 18226 9774
rect 19406 9762 19458 9774
rect 19518 9826 19570 9838
rect 19518 9762 19570 9774
rect 21758 9826 21810 9838
rect 31838 9826 31890 9838
rect 24882 9774 24894 9826
rect 24946 9774 24958 9826
rect 25330 9774 25342 9826
rect 25394 9774 25406 9826
rect 27570 9774 27582 9826
rect 27634 9774 27646 9826
rect 28018 9774 28030 9826
rect 28082 9774 28094 9826
rect 31154 9774 31166 9826
rect 31218 9774 31230 9826
rect 21758 9762 21810 9774
rect 31838 9762 31890 9774
rect 32958 9826 33010 9838
rect 32958 9762 33010 9774
rect 33294 9826 33346 9838
rect 33294 9762 33346 9774
rect 33518 9826 33570 9838
rect 33518 9762 33570 9774
rect 33854 9826 33906 9838
rect 33854 9762 33906 9774
rect 35646 9826 35698 9838
rect 35646 9762 35698 9774
rect 35870 9826 35922 9838
rect 35870 9762 35922 9774
rect 36094 9826 36146 9838
rect 42926 9826 42978 9838
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 36094 9762 36146 9774
rect 42926 9762 42978 9774
rect 43822 9826 43874 9838
rect 43822 9762 43874 9774
rect 50766 9826 50818 9838
rect 50766 9762 50818 9774
rect 52558 9826 52610 9838
rect 52558 9762 52610 9774
rect 52894 9826 52946 9838
rect 52894 9762 52946 9774
rect 53230 9826 53282 9838
rect 53230 9762 53282 9774
rect 18622 9714 18674 9726
rect 26462 9714 26514 9726
rect 29934 9714 29986 9726
rect 23426 9662 23438 9714
rect 23490 9662 23502 9714
rect 28578 9662 28590 9714
rect 28642 9662 28654 9714
rect 18622 9650 18674 9662
rect 26462 9650 26514 9662
rect 29934 9650 29986 9662
rect 30718 9714 30770 9726
rect 32846 9714 32898 9726
rect 31490 9662 31502 9714
rect 31554 9662 31566 9714
rect 30718 9650 30770 9662
rect 32846 9650 32898 9662
rect 34190 9714 34242 9726
rect 34190 9650 34242 9662
rect 34526 9714 34578 9726
rect 34526 9650 34578 9662
rect 36542 9714 36594 9726
rect 40350 9714 40402 9726
rect 37762 9662 37774 9714
rect 37826 9662 37838 9714
rect 39554 9662 39566 9714
rect 39618 9662 39630 9714
rect 36542 9650 36594 9662
rect 40350 9650 40402 9662
rect 50878 9714 50930 9726
rect 50878 9650 50930 9662
rect 51102 9714 51154 9726
rect 51102 9650 51154 9662
rect 51438 9714 51490 9726
rect 51438 9650 51490 9662
rect 15822 9602 15874 9614
rect 15822 9538 15874 9550
rect 19070 9602 19122 9614
rect 30046 9602 30098 9614
rect 21410 9550 21422 9602
rect 21474 9550 21486 9602
rect 27570 9550 27582 9602
rect 27634 9550 27646 9602
rect 19070 9538 19122 9550
rect 30046 9538 30098 9550
rect 30382 9602 30434 9614
rect 30382 9538 30434 9550
rect 30606 9602 30658 9614
rect 30606 9538 30658 9550
rect 32622 9602 32674 9614
rect 32622 9538 32674 9550
rect 33518 9602 33570 9614
rect 50430 9602 50482 9614
rect 44146 9550 44158 9602
rect 44210 9550 44222 9602
rect 33518 9538 33570 9550
rect 50430 9538 50482 9550
rect 52894 9602 52946 9614
rect 52894 9538 52946 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 17502 9266 17554 9278
rect 17502 9202 17554 9214
rect 18734 9266 18786 9278
rect 18734 9202 18786 9214
rect 18846 9266 18898 9278
rect 31390 9266 31442 9278
rect 22082 9214 22094 9266
rect 22146 9214 22158 9266
rect 18846 9202 18898 9214
rect 31390 9202 31442 9214
rect 33294 9266 33346 9278
rect 33294 9202 33346 9214
rect 33854 9266 33906 9278
rect 33854 9202 33906 9214
rect 39230 9266 39282 9278
rect 39230 9202 39282 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 41918 9266 41970 9278
rect 41918 9202 41970 9214
rect 42478 9266 42530 9278
rect 42478 9202 42530 9214
rect 42814 9266 42866 9278
rect 42814 9202 42866 9214
rect 43486 9266 43538 9278
rect 43486 9202 43538 9214
rect 44382 9266 44434 9278
rect 44382 9202 44434 9214
rect 50206 9266 50258 9278
rect 50206 9202 50258 9214
rect 55694 9266 55746 9278
rect 55694 9202 55746 9214
rect 18958 9154 19010 9166
rect 33518 9154 33570 9166
rect 14690 9102 14702 9154
rect 14754 9102 14766 9154
rect 31042 9102 31054 9154
rect 31106 9102 31118 9154
rect 18958 9090 19010 9102
rect 33518 9090 33570 9102
rect 33630 9154 33682 9166
rect 33630 9090 33682 9102
rect 35534 9154 35586 9166
rect 35534 9090 35586 9102
rect 37102 9154 37154 9166
rect 37102 9090 37154 9102
rect 37326 9154 37378 9166
rect 37326 9090 37378 9102
rect 37662 9154 37714 9166
rect 37662 9090 37714 9102
rect 39566 9154 39618 9166
rect 39890 9102 39902 9154
rect 39954 9102 39966 9154
rect 42130 9102 42142 9154
rect 42194 9102 42206 9154
rect 43138 9102 43150 9154
rect 43202 9102 43214 9154
rect 43810 9102 43822 9154
rect 43874 9102 43886 9154
rect 54450 9102 54462 9154
rect 54514 9102 54526 9154
rect 39566 9090 39618 9102
rect 22430 9042 22482 9054
rect 14018 8990 14030 9042
rect 14082 8990 14094 9042
rect 19282 8990 19294 9042
rect 19346 8990 19358 9042
rect 22430 8978 22482 8990
rect 35086 9042 35138 9054
rect 35086 8978 35138 8990
rect 35310 9042 35362 9054
rect 49758 9042 49810 9054
rect 44706 8990 44718 9042
rect 44770 8990 44782 9042
rect 35310 8978 35362 8990
rect 49758 8978 49810 8990
rect 50430 9042 50482 9054
rect 55234 8990 55246 9042
rect 55298 8990 55310 9042
rect 50430 8978 50482 8990
rect 35422 8930 35474 8942
rect 16818 8878 16830 8930
rect 16882 8878 16894 8930
rect 35422 8866 35474 8878
rect 37550 8930 37602 8942
rect 50318 8930 50370 8942
rect 45490 8878 45502 8930
rect 45554 8878 45566 8930
rect 47618 8878 47630 8930
rect 47682 8878 47694 8930
rect 52322 8878 52334 8930
rect 52386 8878 52398 8930
rect 37550 8866 37602 8878
rect 50318 8866 50370 8878
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 35310 8482 35362 8494
rect 35310 8418 35362 8430
rect 33630 8370 33682 8382
rect 33630 8306 33682 8318
rect 47518 8370 47570 8382
rect 51102 8370 51154 8382
rect 50194 8318 50206 8370
rect 50258 8318 50270 8370
rect 47518 8306 47570 8318
rect 51102 8306 51154 8318
rect 26910 8258 26962 8270
rect 26910 8194 26962 8206
rect 27358 8258 27410 8270
rect 27358 8194 27410 8206
rect 30942 8258 30994 8270
rect 30942 8194 30994 8206
rect 31502 8258 31554 8270
rect 31502 8194 31554 8206
rect 32174 8258 32226 8270
rect 35534 8258 35586 8270
rect 33954 8206 33966 8258
rect 34018 8206 34030 8258
rect 32174 8194 32226 8206
rect 35534 8194 35586 8206
rect 35870 8258 35922 8270
rect 35870 8194 35922 8206
rect 44942 8258 44994 8270
rect 44942 8194 44994 8206
rect 45166 8258 45218 8270
rect 45166 8194 45218 8206
rect 45614 8258 45666 8270
rect 45614 8194 45666 8206
rect 45838 8258 45890 8270
rect 45838 8194 45890 8206
rect 46286 8258 46338 8270
rect 46286 8194 46338 8206
rect 46398 8258 46450 8270
rect 46398 8194 46450 8206
rect 47294 8258 47346 8270
rect 47294 8194 47346 8206
rect 47630 8258 47682 8270
rect 47630 8194 47682 8206
rect 48526 8258 48578 8270
rect 48526 8194 48578 8206
rect 48750 8258 48802 8270
rect 48750 8194 48802 8206
rect 48974 8258 49026 8270
rect 51326 8258 51378 8270
rect 49634 8206 49646 8258
rect 49698 8206 49710 8258
rect 50754 8206 50766 8258
rect 50818 8206 50830 8258
rect 48974 8194 49026 8206
rect 51326 8194 51378 8206
rect 30606 8146 30658 8158
rect 30606 8082 30658 8094
rect 31166 8146 31218 8158
rect 31166 8082 31218 8094
rect 36318 8146 36370 8158
rect 36318 8082 36370 8094
rect 39006 8146 39058 8158
rect 39006 8082 39058 8094
rect 39678 8146 39730 8158
rect 39678 8082 39730 8094
rect 47966 8146 48018 8158
rect 47966 8082 48018 8094
rect 48302 8146 48354 8158
rect 49970 8094 49982 8146
rect 50034 8094 50046 8146
rect 48302 8082 48354 8094
rect 26686 8034 26738 8046
rect 26686 7970 26738 7982
rect 26798 8034 26850 8046
rect 26798 7970 26850 7982
rect 30718 8034 30770 8046
rect 30718 7970 30770 7982
rect 31614 8034 31666 8046
rect 31614 7970 31666 7982
rect 31726 8034 31778 8046
rect 31726 7970 31778 7982
rect 32510 8034 32562 8046
rect 32510 7970 32562 7982
rect 33742 8034 33794 8046
rect 35982 8034 36034 8046
rect 34962 7982 34974 8034
rect 35026 7982 35038 8034
rect 33742 7970 33794 7982
rect 35982 7970 36034 7982
rect 36094 8034 36146 8046
rect 45502 8034 45554 8046
rect 39330 7982 39342 8034
rect 39394 7982 39406 8034
rect 36094 7970 36146 7982
rect 45502 7970 45554 7982
rect 46174 8034 46226 8046
rect 46174 7970 46226 7982
rect 46622 8034 46674 8046
rect 46622 7970 46674 7982
rect 49422 8034 49474 8046
rect 51650 7982 51662 8034
rect 51714 7982 51726 8034
rect 49422 7970 49474 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 19070 7698 19122 7710
rect 19070 7634 19122 7646
rect 24782 7698 24834 7710
rect 24782 7634 24834 7646
rect 31502 7698 31554 7710
rect 31502 7634 31554 7646
rect 38446 7698 38498 7710
rect 38446 7634 38498 7646
rect 38894 7698 38946 7710
rect 38894 7634 38946 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 41246 7698 41298 7710
rect 41246 7634 41298 7646
rect 41470 7698 41522 7710
rect 41470 7634 41522 7646
rect 43598 7698 43650 7710
rect 43598 7634 43650 7646
rect 45838 7698 45890 7710
rect 45838 7634 45890 7646
rect 50094 7698 50146 7710
rect 50094 7634 50146 7646
rect 18734 7586 18786 7598
rect 18734 7522 18786 7534
rect 19294 7586 19346 7598
rect 19294 7522 19346 7534
rect 26798 7586 26850 7598
rect 33966 7586 34018 7598
rect 29810 7534 29822 7586
rect 29874 7534 29886 7586
rect 26798 7522 26850 7534
rect 33966 7522 34018 7534
rect 35646 7586 35698 7598
rect 39790 7586 39842 7598
rect 36418 7534 36430 7586
rect 36482 7534 36494 7586
rect 35646 7522 35698 7534
rect 39790 7522 39842 7534
rect 40126 7586 40178 7598
rect 50878 7586 50930 7598
rect 43250 7534 43262 7586
rect 43314 7534 43326 7586
rect 51202 7534 51214 7586
rect 51266 7534 51278 7586
rect 40126 7522 40178 7534
rect 50878 7522 50930 7534
rect 18958 7474 19010 7486
rect 23326 7474 23378 7486
rect 19618 7422 19630 7474
rect 19682 7422 19694 7474
rect 18958 7410 19010 7422
rect 23326 7410 23378 7422
rect 24334 7474 24386 7486
rect 24334 7410 24386 7422
rect 26350 7474 26402 7486
rect 26350 7410 26402 7422
rect 26574 7474 26626 7486
rect 26574 7410 26626 7422
rect 27022 7474 27074 7486
rect 27022 7410 27074 7422
rect 27246 7474 27298 7486
rect 33630 7474 33682 7486
rect 30482 7422 30494 7474
rect 30546 7422 30558 7474
rect 27246 7410 27298 7422
rect 33630 7410 33682 7422
rect 33742 7474 33794 7486
rect 34414 7474 34466 7486
rect 35310 7474 35362 7486
rect 36094 7474 36146 7486
rect 34290 7422 34302 7474
rect 34354 7422 34366 7474
rect 34626 7422 34638 7474
rect 34690 7422 34702 7474
rect 35074 7422 35086 7474
rect 35138 7422 35150 7474
rect 35410 7422 35422 7474
rect 35474 7422 35486 7474
rect 33742 7410 33794 7422
rect 34414 7410 34466 7422
rect 35310 7410 35362 7422
rect 36094 7410 36146 7422
rect 36766 7474 36818 7486
rect 36766 7410 36818 7422
rect 37886 7474 37938 7486
rect 37886 7410 37938 7422
rect 38110 7474 38162 7486
rect 38110 7410 38162 7422
rect 38670 7474 38722 7486
rect 38670 7410 38722 7422
rect 40350 7474 40402 7486
rect 40350 7410 40402 7422
rect 40798 7474 40850 7486
rect 40798 7410 40850 7422
rect 42926 7474 42978 7486
rect 42926 7410 42978 7422
rect 43822 7474 43874 7486
rect 49646 7474 49698 7486
rect 44146 7422 44158 7474
rect 44210 7422 44222 7474
rect 43822 7410 43874 7422
rect 49646 7410 49698 7422
rect 49870 7474 49922 7486
rect 49870 7410 49922 7422
rect 50542 7474 50594 7486
rect 50542 7410 50594 7422
rect 50654 7474 50706 7486
rect 50654 7410 50706 7422
rect 51438 7474 51490 7486
rect 51438 7410 51490 7422
rect 20190 7362 20242 7374
rect 20190 7298 20242 7310
rect 21086 7362 21138 7374
rect 21086 7298 21138 7310
rect 21310 7362 21362 7374
rect 21310 7298 21362 7310
rect 23662 7362 23714 7374
rect 31838 7362 31890 7374
rect 25778 7310 25790 7362
rect 25842 7310 25854 7362
rect 27682 7310 27694 7362
rect 27746 7310 27758 7362
rect 23662 7298 23714 7310
rect 31838 7298 31890 7310
rect 38558 7362 38610 7374
rect 38558 7298 38610 7310
rect 41358 7362 41410 7374
rect 41358 7298 41410 7310
rect 42590 7362 42642 7374
rect 42590 7298 42642 7310
rect 43710 7362 43762 7374
rect 44606 7362 44658 7374
rect 44146 7310 44158 7362
rect 44210 7359 44222 7362
rect 44210 7313 44319 7359
rect 44210 7310 44222 7313
rect 43710 7298 43762 7310
rect 19966 7250 20018 7262
rect 23102 7250 23154 7262
rect 20738 7198 20750 7250
rect 20802 7198 20814 7250
rect 22754 7198 22766 7250
rect 22818 7198 22830 7250
rect 19966 7186 20018 7198
rect 23102 7186 23154 7198
rect 23886 7250 23938 7262
rect 23886 7186 23938 7198
rect 24110 7250 24162 7262
rect 24110 7186 24162 7198
rect 26126 7250 26178 7262
rect 26126 7186 26178 7198
rect 35982 7250 36034 7262
rect 37538 7198 37550 7250
rect 37602 7198 37614 7250
rect 44273 7247 44319 7313
rect 44606 7298 44658 7310
rect 49758 7362 49810 7374
rect 52446 7362 52498 7374
rect 51538 7310 51550 7362
rect 51602 7310 51614 7362
rect 49758 7298 49810 7310
rect 52446 7298 52498 7310
rect 52558 7250 52610 7262
rect 44594 7247 44606 7250
rect 44273 7201 44606 7247
rect 44594 7198 44606 7201
rect 44658 7198 44670 7250
rect 35982 7186 36034 7198
rect 52558 7186 52610 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 19518 6914 19570 6926
rect 19518 6850 19570 6862
rect 21422 6914 21474 6926
rect 21422 6850 21474 6862
rect 23550 6914 23602 6926
rect 23550 6850 23602 6862
rect 26798 6914 26850 6926
rect 26798 6850 26850 6862
rect 26910 6914 26962 6926
rect 38782 6914 38834 6926
rect 32274 6911 32286 6914
rect 26910 6850 26962 6862
rect 31953 6865 32286 6911
rect 31953 6802 31999 6865
rect 32274 6862 32286 6865
rect 32338 6862 32350 6914
rect 38782 6850 38834 6862
rect 38894 6914 38946 6926
rect 38894 6850 38946 6862
rect 40798 6914 40850 6926
rect 40798 6850 40850 6862
rect 40910 6914 40962 6926
rect 40910 6850 40962 6862
rect 41582 6914 41634 6926
rect 41582 6850 41634 6862
rect 50318 6914 50370 6926
rect 50318 6850 50370 6862
rect 32286 6802 32338 6814
rect 18274 6750 18286 6802
rect 18338 6750 18350 6802
rect 18610 6750 18622 6802
rect 18674 6750 18686 6802
rect 22194 6750 22206 6802
rect 22258 6750 22270 6802
rect 24322 6750 24334 6802
rect 24386 6750 24398 6802
rect 31938 6750 31950 6802
rect 32002 6750 32014 6802
rect 32286 6738 32338 6750
rect 36206 6802 36258 6814
rect 36206 6738 36258 6750
rect 46398 6802 46450 6814
rect 46398 6738 46450 6750
rect 48750 6802 48802 6814
rect 48750 6738 48802 6750
rect 49758 6802 49810 6814
rect 49758 6738 49810 6750
rect 50430 6802 50482 6814
rect 52658 6750 52670 6802
rect 52722 6750 52734 6802
rect 50430 6738 50482 6750
rect 18734 6690 18786 6702
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 18734 6626 18786 6638
rect 19630 6690 19682 6702
rect 19630 6626 19682 6638
rect 20526 6690 20578 6702
rect 20526 6626 20578 6638
rect 20638 6690 20690 6702
rect 20638 6626 20690 6638
rect 21310 6690 21362 6702
rect 23438 6690 23490 6702
rect 25454 6690 25506 6702
rect 27582 6690 27634 6702
rect 22306 6638 22318 6690
rect 22370 6638 22382 6690
rect 24434 6638 24446 6690
rect 24498 6638 24510 6690
rect 25890 6638 25902 6690
rect 25954 6638 25966 6690
rect 21310 6626 21362 6638
rect 23438 6626 23490 6638
rect 25454 6626 25506 6638
rect 27582 6626 27634 6638
rect 28030 6690 28082 6702
rect 28030 6626 28082 6638
rect 30942 6690 30994 6702
rect 30942 6626 30994 6638
rect 31278 6690 31330 6702
rect 31278 6626 31330 6638
rect 31950 6690 32002 6702
rect 41806 6690 41858 6702
rect 37874 6638 37886 6690
rect 37938 6638 37950 6690
rect 38210 6638 38222 6690
rect 38274 6638 38286 6690
rect 41234 6638 41246 6690
rect 41298 6638 41310 6690
rect 31950 6626 32002 6638
rect 41806 6626 41858 6638
rect 43486 6690 43538 6702
rect 43486 6626 43538 6638
rect 43934 6690 43986 6702
rect 43934 6626 43986 6638
rect 46846 6690 46898 6702
rect 46846 6626 46898 6638
rect 48414 6690 48466 6702
rect 48414 6626 48466 6638
rect 49982 6690 50034 6702
rect 56030 6690 56082 6702
rect 50978 6638 50990 6690
rect 51042 6638 51054 6690
rect 54786 6638 54798 6690
rect 54850 6638 54862 6690
rect 55458 6638 55470 6690
rect 55522 6638 55534 6690
rect 49982 6626 50034 6638
rect 56030 6626 56082 6638
rect 19294 6578 19346 6590
rect 24782 6578 24834 6590
rect 16146 6526 16158 6578
rect 16210 6526 16222 6578
rect 18946 6526 18958 6578
rect 19010 6526 19022 6578
rect 21970 6526 21982 6578
rect 22034 6526 22046 6578
rect 24098 6526 24110 6578
rect 24162 6526 24174 6578
rect 19294 6514 19346 6526
rect 24782 6514 24834 6526
rect 25006 6578 25058 6590
rect 31502 6578 31554 6590
rect 26226 6526 26238 6578
rect 26290 6526 26302 6578
rect 27234 6526 27246 6578
rect 27298 6526 27310 6578
rect 25006 6514 25058 6526
rect 31502 6514 31554 6526
rect 38558 6578 38610 6590
rect 38558 6514 38610 6526
rect 40014 6578 40066 6590
rect 40462 6578 40514 6590
rect 40226 6526 40238 6578
rect 40290 6526 40302 6578
rect 40014 6514 40066 6526
rect 40462 6514 40514 6526
rect 42926 6578 42978 6590
rect 42926 6514 42978 6526
rect 43262 6578 43314 6590
rect 43262 6514 43314 6526
rect 48526 6578 48578 6590
rect 48526 6514 48578 6526
rect 48862 6578 48914 6590
rect 50766 6578 50818 6590
rect 49410 6526 49422 6578
rect 49474 6526 49486 6578
rect 48862 6514 48914 6526
rect 50766 6514 50818 6526
rect 51214 6578 51266 6590
rect 51214 6514 51266 6526
rect 20302 6466 20354 6478
rect 20302 6402 20354 6414
rect 20750 6466 20802 6478
rect 20750 6402 20802 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 23886 6466 23938 6478
rect 23886 6402 23938 6414
rect 25118 6466 25170 6478
rect 25118 6402 25170 6414
rect 26126 6466 26178 6478
rect 26126 6402 26178 6414
rect 26462 6466 26514 6478
rect 26462 6402 26514 6414
rect 30158 6466 30210 6478
rect 30158 6402 30210 6414
rect 30494 6466 30546 6478
rect 30494 6402 30546 6414
rect 30718 6466 30770 6478
rect 30718 6402 30770 6414
rect 30830 6466 30882 6478
rect 30830 6402 30882 6414
rect 31390 6466 31442 6478
rect 31390 6402 31442 6414
rect 38110 6466 38162 6478
rect 38110 6402 38162 6414
rect 40126 6466 40178 6478
rect 40126 6402 40178 6414
rect 43150 6466 43202 6478
rect 43150 6402 43202 6414
rect 51102 6466 51154 6478
rect 51102 6402 51154 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 17390 6130 17442 6142
rect 17390 6066 17442 6078
rect 18510 6130 18562 6142
rect 18510 6066 18562 6078
rect 18846 6130 18898 6142
rect 18846 6066 18898 6078
rect 21646 6130 21698 6142
rect 21646 6066 21698 6078
rect 23662 6130 23714 6142
rect 23662 6066 23714 6078
rect 23774 6130 23826 6142
rect 23774 6066 23826 6078
rect 23998 6130 24050 6142
rect 31278 6130 31330 6142
rect 30818 6127 30830 6130
rect 23998 6066 24050 6078
rect 30721 6081 30830 6127
rect 17502 6018 17554 6030
rect 17502 5954 17554 5966
rect 19070 6018 19122 6030
rect 19070 5954 19122 5966
rect 21534 6018 21586 6030
rect 21534 5954 21586 5966
rect 22094 6018 22146 6030
rect 22094 5954 22146 5966
rect 21758 5906 21810 5918
rect 19394 5854 19406 5906
rect 19458 5854 19470 5906
rect 21758 5842 21810 5854
rect 23550 5906 23602 5918
rect 30370 5854 30382 5906
rect 30434 5854 30446 5906
rect 23550 5842 23602 5854
rect 18958 5794 19010 5806
rect 30721 5794 30767 6081
rect 30818 6078 30830 6081
rect 30882 6078 30894 6130
rect 31278 6066 31330 6078
rect 32174 6130 32226 6142
rect 32174 6066 32226 6078
rect 32510 6130 32562 6142
rect 32510 6066 32562 6078
rect 46286 6130 46338 6142
rect 46286 6066 46338 6078
rect 31614 6018 31666 6030
rect 31614 5954 31666 5966
rect 33854 6018 33906 6030
rect 33854 5954 33906 5966
rect 35422 6018 35474 6030
rect 46174 6018 46226 6030
rect 43698 5966 43710 6018
rect 43762 5966 43774 6018
rect 35422 5954 35474 5966
rect 46174 5954 46226 5966
rect 46510 6018 46562 6030
rect 46510 5954 46562 5966
rect 46958 6018 47010 6030
rect 46958 5954 47010 5966
rect 47070 6018 47122 6030
rect 47170 5966 47182 6018
rect 47234 5966 47246 6018
rect 47070 5954 47122 5966
rect 30942 5906 30994 5918
rect 30942 5842 30994 5854
rect 31390 5906 31442 5918
rect 45054 5906 45106 5918
rect 44370 5854 44382 5906
rect 44434 5854 44446 5906
rect 31390 5842 31442 5854
rect 45054 5842 45106 5854
rect 45278 5906 45330 5918
rect 45278 5842 45330 5854
rect 45614 5906 45666 5918
rect 45614 5842 45666 5854
rect 46734 5906 46786 5918
rect 46734 5842 46786 5854
rect 41246 5794 41298 5806
rect 45166 5794 45218 5806
rect 27570 5742 27582 5794
rect 27634 5742 27646 5794
rect 29698 5742 29710 5794
rect 29762 5742 29774 5794
rect 30706 5742 30718 5794
rect 30770 5742 30782 5794
rect 41570 5742 41582 5794
rect 41634 5742 41646 5794
rect 47506 5742 47518 5794
rect 47570 5742 47582 5794
rect 18958 5730 19010 5742
rect 41246 5730 41298 5742
rect 45166 5730 45218 5742
rect 33742 5682 33794 5694
rect 33742 5618 33794 5630
rect 35534 5682 35586 5694
rect 35534 5618 35586 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 20190 5234 20242 5246
rect 20190 5170 20242 5182
rect 21422 5234 21474 5246
rect 21422 5170 21474 5182
rect 23214 5234 23266 5246
rect 23214 5170 23266 5182
rect 26126 5234 26178 5246
rect 26126 5170 26178 5182
rect 31054 5234 31106 5246
rect 31054 5170 31106 5182
rect 31614 5234 31666 5246
rect 31614 5170 31666 5182
rect 32062 5234 32114 5246
rect 40350 5234 40402 5246
rect 33506 5182 33518 5234
rect 33570 5182 33582 5234
rect 35634 5182 35646 5234
rect 35698 5182 35710 5234
rect 36978 5182 36990 5234
rect 37042 5182 37054 5234
rect 32062 5170 32114 5182
rect 40350 5170 40402 5182
rect 40686 5234 40738 5246
rect 40686 5170 40738 5182
rect 44046 5234 44098 5246
rect 44046 5170 44098 5182
rect 44942 5234 44994 5246
rect 51214 5234 51266 5246
rect 47730 5182 47742 5234
rect 47794 5182 47806 5234
rect 49858 5182 49870 5234
rect 49922 5182 49934 5234
rect 44942 5170 44994 5182
rect 51214 5170 51266 5182
rect 30718 5122 30770 5134
rect 30718 5058 30770 5070
rect 30942 5122 30994 5134
rect 30942 5058 30994 5070
rect 31166 5122 31218 5134
rect 45502 5122 45554 5134
rect 32722 5070 32734 5122
rect 32786 5070 32798 5122
rect 39106 5070 39118 5122
rect 39170 5070 39182 5122
rect 39778 5070 39790 5122
rect 39842 5070 39854 5122
rect 31166 5058 31218 5070
rect 45502 5058 45554 5070
rect 45838 5122 45890 5134
rect 50318 5122 50370 5134
rect 46386 5070 46398 5122
rect 46450 5070 46462 5122
rect 47058 5070 47070 5122
rect 47122 5070 47134 5122
rect 45838 5058 45890 5070
rect 50318 5058 50370 5070
rect 20078 4898 20130 4910
rect 20078 4834 20130 4846
rect 23102 4898 23154 4910
rect 23102 4834 23154 4846
rect 26014 4898 26066 4910
rect 26014 4834 26066 4846
rect 40798 4898 40850 4910
rect 40798 4834 40850 4846
rect 45950 4898 46002 4910
rect 45950 4834 46002 4846
rect 46062 4898 46114 4910
rect 46062 4834 46114 4846
rect 51326 4898 51378 4910
rect 51326 4834 51378 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 28590 4562 28642 4574
rect 28590 4498 28642 4510
rect 33182 4562 33234 4574
rect 33182 4498 33234 4510
rect 37662 4562 37714 4574
rect 37662 4498 37714 4510
rect 38222 4562 38274 4574
rect 38222 4498 38274 4510
rect 48750 4562 48802 4574
rect 48750 4498 48802 4510
rect 53902 4562 53954 4574
rect 53902 4498 53954 4510
rect 38110 4450 38162 4462
rect 48862 4450 48914 4462
rect 19170 4398 19182 4450
rect 19234 4398 19246 4450
rect 22418 4398 22430 4450
rect 22482 4398 22494 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 31490 4398 31502 4450
rect 31554 4398 31566 4450
rect 36418 4398 36430 4450
rect 36482 4398 36494 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 44930 4398 44942 4450
rect 44994 4398 45006 4450
rect 52658 4398 52670 4450
rect 52722 4398 52734 4450
rect 38110 4386 38162 4398
rect 48862 4386 48914 4398
rect 57598 4338 57650 4350
rect 18498 4286 18510 4338
rect 18562 4286 18574 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 32274 4286 32286 4338
rect 32338 4286 32350 4338
rect 37202 4286 37214 4338
rect 37266 4286 37278 4338
rect 40898 4286 40910 4338
rect 40962 4286 40974 4338
rect 44146 4286 44158 4338
rect 44210 4286 44222 4338
rect 53330 4286 53342 4338
rect 53394 4286 53406 4338
rect 57598 4274 57650 4286
rect 58158 4338 58210 4350
rect 58158 4274 58210 4286
rect 57374 4226 57426 4238
rect 21298 4174 21310 4226
rect 21362 4174 21374 4226
rect 24546 4174 24558 4226
rect 24610 4174 24622 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 29362 4174 29374 4226
rect 29426 4174 29438 4226
rect 34290 4174 34302 4226
rect 34354 4174 34366 4226
rect 43810 4174 43822 4226
rect 43874 4174 43886 4226
rect 47058 4174 47070 4226
rect 47122 4174 47134 4226
rect 50530 4174 50542 4226
rect 50594 4174 50606 4226
rect 57374 4162 57426 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 21646 3666 21698 3678
rect 21646 3602 21698 3614
rect 43934 3666 43986 3678
rect 43934 3602 43986 3614
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 8766 66782 8818 66834
rect 9326 66782 9378 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 26126 66446 26178 66498
rect 40798 66446 40850 66498
rect 43822 66446 43874 66498
rect 48414 66446 48466 66498
rect 52222 66446 52274 66498
rect 56030 66446 56082 66498
rect 18846 66334 18898 66386
rect 22878 66334 22930 66386
rect 36990 66334 37042 66386
rect 17614 66222 17666 66274
rect 23550 66222 23602 66274
rect 25118 66222 25170 66274
rect 39230 66222 39282 66274
rect 39790 66222 39842 66274
rect 46174 66222 46226 66274
rect 47406 66222 47458 66274
rect 51214 66222 51266 66274
rect 55022 66222 55074 66274
rect 2942 66110 2994 66162
rect 5518 66110 5570 66162
rect 6974 66110 7026 66162
rect 9326 66110 9378 66162
rect 11006 66110 11058 66162
rect 13134 66110 13186 66162
rect 15038 66110 15090 66162
rect 17054 66110 17106 66162
rect 29150 66110 29202 66162
rect 31166 66110 31218 66162
rect 33182 66110 33234 66162
rect 35198 66110 35250 66162
rect 43038 66110 43090 66162
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 34862 65550 34914 65602
rect 57822 65550 57874 65602
rect 20190 65438 20242 65490
rect 21870 65438 21922 65490
rect 29710 65438 29762 65490
rect 35534 65438 35586 65490
rect 36654 65438 36706 65490
rect 44382 65438 44434 65490
rect 44830 65438 44882 65490
rect 48862 65438 48914 65490
rect 54910 65438 54962 65490
rect 57598 65438 57650 65490
rect 58158 65438 58210 65490
rect 12574 65326 12626 65378
rect 13246 65326 13298 65378
rect 17390 65326 17442 65378
rect 19518 65326 19570 65378
rect 20862 65326 20914 65378
rect 22542 65326 22594 65378
rect 24670 65326 24722 65378
rect 25454 65326 25506 65378
rect 27358 65326 27410 65378
rect 30270 65326 30322 65378
rect 34974 65326 35026 65378
rect 37438 65326 37490 65378
rect 39566 65326 39618 65378
rect 40126 65326 40178 65378
rect 41134 65326 41186 65378
rect 41582 65326 41634 65378
rect 43710 65326 43762 65378
rect 45614 65326 45666 65378
rect 47742 65326 47794 65378
rect 49534 65326 49586 65378
rect 51662 65326 51714 65378
rect 51998 65326 52050 65378
rect 54126 65326 54178 65378
rect 55470 65326 55522 65378
rect 35086 65214 35138 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 23550 64878 23602 64930
rect 42702 64878 42754 64930
rect 47518 64878 47570 64930
rect 50206 64878 50258 64930
rect 51774 64878 51826 64930
rect 8542 64766 8594 64818
rect 10110 64766 10162 64818
rect 12238 64766 12290 64818
rect 12798 64766 12850 64818
rect 16382 64766 16434 64818
rect 20750 64766 20802 64818
rect 26910 64766 26962 64818
rect 33518 64766 33570 64818
rect 35646 64766 35698 64818
rect 41358 64766 41410 64818
rect 44942 64766 44994 64818
rect 45390 64766 45442 64818
rect 54910 64766 54962 64818
rect 55246 64766 55298 64818
rect 5742 64654 5794 64706
rect 8878 64654 8930 64706
rect 9438 64654 9490 64706
rect 13582 64654 13634 64706
rect 16830 64654 16882 64706
rect 17950 64654 18002 64706
rect 23998 64654 24050 64706
rect 27918 64654 27970 64706
rect 29038 64654 29090 64706
rect 29486 64654 29538 64706
rect 30382 64654 30434 64706
rect 36430 64654 36482 64706
rect 37102 64654 37154 64706
rect 38558 64654 38610 64706
rect 41694 64654 41746 64706
rect 49422 64654 49474 64706
rect 58158 64654 58210 64706
rect 6414 64542 6466 64594
rect 12574 64542 12626 64594
rect 14254 64542 14306 64594
rect 18622 64542 18674 64594
rect 23662 64542 23714 64594
rect 24782 64542 24834 64594
rect 30942 64542 30994 64594
rect 32510 64542 32562 64594
rect 32622 64542 32674 64594
rect 32958 64542 33010 64594
rect 39230 64542 39282 64594
rect 50318 64542 50370 64594
rect 51662 64542 51714 64594
rect 57374 64542 57426 64594
rect 8990 64430 9042 64482
rect 12798 64430 12850 64482
rect 21422 64430 21474 64482
rect 23214 64430 23266 64482
rect 27246 64430 27298 64482
rect 27358 64430 27410 64482
rect 27470 64430 27522 64482
rect 28702 64430 28754 64482
rect 29598 64430 29650 64482
rect 29710 64430 29762 64482
rect 30830 64430 30882 64482
rect 31054 64430 31106 64482
rect 31502 64430 31554 64482
rect 32286 64430 32338 64482
rect 33070 64430 33122 64482
rect 33294 64430 33346 64482
rect 52782 64430 52834 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 8766 64094 8818 64146
rect 11342 64094 11394 64146
rect 17614 64094 17666 64146
rect 27806 64094 27858 64146
rect 32286 64094 32338 64146
rect 41582 64094 41634 64146
rect 42030 64094 42082 64146
rect 46958 64094 47010 64146
rect 50430 64094 50482 64146
rect 52334 64094 52386 64146
rect 54574 64094 54626 64146
rect 12910 63982 12962 64034
rect 13694 63982 13746 64034
rect 13806 63982 13858 64034
rect 14142 63982 14194 64034
rect 27470 63982 27522 64034
rect 27582 63982 27634 64034
rect 31950 63982 32002 64034
rect 35198 63982 35250 64034
rect 46062 63982 46114 64034
rect 50878 63982 50930 64034
rect 51214 63982 51266 64034
rect 55246 63982 55298 64034
rect 55806 63982 55858 64034
rect 11678 63870 11730 63922
rect 12574 63870 12626 63922
rect 14254 63870 14306 63922
rect 17278 63870 17330 63922
rect 17614 63870 17666 63922
rect 17838 63870 17890 63922
rect 20190 63870 20242 63922
rect 23438 63870 23490 63922
rect 26686 63870 26738 63922
rect 28030 63870 28082 63922
rect 32062 63870 32114 63922
rect 32510 63870 32562 63922
rect 33518 63870 33570 63922
rect 34638 63870 34690 63922
rect 39454 63870 39506 63922
rect 43374 63870 43426 63922
rect 43822 63870 43874 63922
rect 45950 63870 46002 63922
rect 46958 63870 47010 63922
rect 49534 63870 49586 63922
rect 49646 63870 49698 63922
rect 49982 63870 50034 63922
rect 50094 63870 50146 63922
rect 51326 63870 51378 63922
rect 54126 63870 54178 63922
rect 54798 63870 54850 63922
rect 20862 63758 20914 63810
rect 22990 63758 23042 63810
rect 26350 63758 26402 63810
rect 27134 63758 27186 63810
rect 28814 63758 28866 63810
rect 30942 63758 30994 63810
rect 32398 63758 32450 63810
rect 33182 63758 33234 63810
rect 50430 63758 50482 63810
rect 50766 63758 50818 63810
rect 54686 63758 54738 63810
rect 13694 63646 13746 63698
rect 43038 63646 43090 63698
rect 43374 63646 43426 63698
rect 55582 63646 55634 63698
rect 55918 63646 55970 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 19630 63310 19682 63362
rect 22318 63310 22370 63362
rect 53566 63310 53618 63362
rect 54462 63310 54514 63362
rect 6638 63198 6690 63250
rect 12910 63198 12962 63250
rect 17502 63198 17554 63250
rect 26238 63198 26290 63250
rect 32062 63198 32114 63250
rect 45166 63198 45218 63250
rect 47742 63198 47794 63250
rect 51438 63198 51490 63250
rect 51662 63198 51714 63250
rect 53006 63198 53058 63250
rect 53902 63198 53954 63250
rect 54910 63198 54962 63250
rect 55246 63198 55298 63250
rect 57374 63198 57426 63250
rect 6750 63086 6802 63138
rect 7870 63086 7922 63138
rect 8094 63086 8146 63138
rect 15486 63086 15538 63138
rect 16270 63086 16322 63138
rect 18062 63086 18114 63138
rect 19630 63086 19682 63138
rect 21310 63086 21362 63138
rect 26686 63086 26738 63138
rect 27134 63086 27186 63138
rect 27582 63086 27634 63138
rect 27806 63086 27858 63138
rect 28142 63086 28194 63138
rect 30158 63086 30210 63138
rect 30382 63086 30434 63138
rect 32286 63086 32338 63138
rect 32622 63086 32674 63138
rect 41246 63086 41298 63138
rect 43486 63086 43538 63138
rect 44046 63086 44098 63138
rect 44942 63086 44994 63138
rect 46062 63086 46114 63138
rect 46510 63086 46562 63138
rect 50654 63086 50706 63138
rect 50766 63086 50818 63138
rect 51102 63086 51154 63138
rect 51214 63086 51266 63138
rect 51774 63086 51826 63138
rect 53230 63086 53282 63138
rect 54126 63086 54178 63138
rect 58158 63086 58210 63138
rect 6526 62974 6578 63026
rect 7086 62974 7138 63026
rect 7646 62974 7698 63026
rect 12574 62974 12626 63026
rect 12798 62974 12850 63026
rect 14814 62974 14866 63026
rect 16382 62974 16434 63026
rect 17614 62974 17666 63026
rect 19966 62974 20018 63026
rect 26126 62974 26178 63026
rect 26462 62974 26514 63026
rect 28030 62974 28082 63026
rect 29486 62974 29538 63026
rect 31166 62974 31218 63026
rect 31278 62974 31330 63026
rect 41022 62974 41074 63026
rect 42254 62974 42306 63026
rect 44158 62974 44210 63026
rect 45054 62974 45106 63026
rect 45502 62974 45554 63026
rect 45838 62974 45890 63026
rect 17390 62862 17442 62914
rect 18510 62862 18562 62914
rect 27022 62862 27074 62914
rect 27246 62862 27298 62914
rect 28590 62862 28642 62914
rect 31502 62862 31554 62914
rect 32062 62862 32114 62914
rect 32958 62862 33010 62914
rect 42478 62862 42530 62914
rect 42926 62862 42978 62914
rect 44382 62862 44434 62914
rect 45278 62862 45330 62914
rect 47182 62862 47234 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 7198 62526 7250 62578
rect 7310 62526 7362 62578
rect 8542 62526 8594 62578
rect 13134 62526 13186 62578
rect 14926 62526 14978 62578
rect 16494 62526 16546 62578
rect 16718 62526 16770 62578
rect 19406 62526 19458 62578
rect 19966 62526 20018 62578
rect 29038 62526 29090 62578
rect 44046 62526 44098 62578
rect 44718 62526 44770 62578
rect 45502 62526 45554 62578
rect 45614 62526 45666 62578
rect 47182 62526 47234 62578
rect 52110 62526 52162 62578
rect 6862 62414 6914 62466
rect 7870 62414 7922 62466
rect 7982 62414 8034 62466
rect 10894 62414 10946 62466
rect 13582 62414 13634 62466
rect 14814 62414 14866 62466
rect 18958 62414 19010 62466
rect 20862 62414 20914 62466
rect 28926 62414 28978 62466
rect 37886 62414 37938 62466
rect 39454 62414 39506 62466
rect 41918 62414 41970 62466
rect 43262 62414 43314 62466
rect 47294 62414 47346 62466
rect 52446 62414 52498 62466
rect 56590 62414 56642 62466
rect 56702 62414 56754 62466
rect 7086 62302 7138 62354
rect 8206 62302 8258 62354
rect 8430 62302 8482 62354
rect 8766 62302 8818 62354
rect 9438 62302 9490 62354
rect 10222 62302 10274 62354
rect 12910 62302 12962 62354
rect 13694 62302 13746 62354
rect 15150 62302 15202 62354
rect 16382 62302 16434 62354
rect 19182 62302 19234 62354
rect 19518 62302 19570 62354
rect 19854 62302 19906 62354
rect 20078 62302 20130 62354
rect 20414 62302 20466 62354
rect 29150 62302 29202 62354
rect 29374 62302 29426 62354
rect 37214 62302 37266 62354
rect 38782 62302 38834 62354
rect 41246 62302 41298 62354
rect 42814 62302 42866 62354
rect 43486 62302 43538 62354
rect 43934 62302 43986 62354
rect 44158 62302 44210 62354
rect 44606 62302 44658 62354
rect 44942 62302 44994 62354
rect 45054 62302 45106 62354
rect 45726 62302 45778 62354
rect 45950 62302 46002 62354
rect 46286 62302 46338 62354
rect 46510 62302 46562 62354
rect 46958 62302 47010 62354
rect 48862 62302 48914 62354
rect 53454 62302 53506 62354
rect 56926 62302 56978 62354
rect 10558 62190 10610 62242
rect 15598 62190 15650 62242
rect 27694 62190 27746 62242
rect 30830 62190 30882 62242
rect 31278 62190 31330 62242
rect 37438 62190 37490 62242
rect 38558 62190 38610 62242
rect 41022 62190 41074 62242
rect 42478 62190 42530 62242
rect 46174 62190 46226 62242
rect 49534 62190 49586 62242
rect 51662 62190 51714 62242
rect 52894 62190 52946 62242
rect 55358 62190 55410 62242
rect 57262 62190 57314 62242
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 20302 61742 20354 61794
rect 43374 61742 43426 61794
rect 49198 61742 49250 61794
rect 56366 61742 56418 61794
rect 12238 61630 12290 61682
rect 24558 61630 24610 61682
rect 35534 61630 35586 61682
rect 36318 61630 36370 61682
rect 37438 61630 37490 61682
rect 38222 61630 38274 61682
rect 52782 61630 52834 61682
rect 55022 61630 55074 61682
rect 21758 61518 21810 61570
rect 38558 61518 38610 61570
rect 43374 61518 43426 61570
rect 53118 61518 53170 61570
rect 54238 61518 54290 61570
rect 55470 61518 55522 61570
rect 6414 61406 6466 61458
rect 6750 61406 6802 61458
rect 19966 61406 20018 61458
rect 20414 61406 20466 61458
rect 20638 61406 20690 61458
rect 22430 61406 22482 61458
rect 24894 61406 24946 61458
rect 32734 61406 32786 61458
rect 34638 61406 34690 61458
rect 35198 61406 35250 61458
rect 36430 61406 36482 61458
rect 36990 61406 37042 61458
rect 37214 61406 37266 61458
rect 37550 61406 37602 61458
rect 43710 61406 43762 61458
rect 49086 61406 49138 61458
rect 6190 61294 6242 61346
rect 6302 61294 6354 61346
rect 6862 61294 6914 61346
rect 7086 61294 7138 61346
rect 7534 61294 7586 61346
rect 20190 61294 20242 61346
rect 20750 61294 20802 61346
rect 25006 61294 25058 61346
rect 25566 61294 25618 61346
rect 25902 61294 25954 61346
rect 32398 61294 32450 61346
rect 32622 61294 32674 61346
rect 34750 61294 34802 61346
rect 34974 61294 35026 61346
rect 35422 61294 35474 61346
rect 36206 61294 36258 61346
rect 38334 61294 38386 61346
rect 44942 61294 44994 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 7870 60958 7922 61010
rect 25454 60958 25506 61010
rect 26014 60958 26066 61010
rect 32286 60958 32338 61010
rect 40014 60958 40066 61010
rect 42702 60958 42754 61010
rect 49086 60958 49138 61010
rect 49646 60958 49698 61010
rect 50990 60958 51042 61010
rect 57038 60958 57090 61010
rect 57934 60958 57986 61010
rect 6302 60846 6354 60898
rect 11006 60846 11058 60898
rect 11902 60846 11954 60898
rect 13246 60846 13298 60898
rect 17502 60846 17554 60898
rect 17950 60846 18002 60898
rect 18062 60846 18114 60898
rect 20974 60846 21026 60898
rect 27246 60846 27298 60898
rect 27806 60846 27858 60898
rect 29598 60846 29650 60898
rect 35422 60846 35474 60898
rect 36766 60846 36818 60898
rect 39118 60846 39170 60898
rect 54462 60846 54514 60898
rect 55806 60846 55858 60898
rect 56590 60846 56642 60898
rect 2830 60734 2882 60786
rect 6750 60734 6802 60786
rect 7534 60734 7586 60786
rect 10782 60734 10834 60786
rect 11566 60734 11618 60786
rect 11790 60734 11842 60786
rect 12798 60734 12850 60786
rect 13022 60734 13074 60786
rect 13358 60734 13410 60786
rect 17390 60734 17442 60786
rect 17726 60734 17778 60786
rect 21758 60734 21810 60786
rect 22654 60734 22706 60786
rect 25902 60734 25954 60786
rect 26238 60734 26290 60786
rect 27134 60734 27186 60786
rect 27470 60734 27522 60786
rect 27694 60734 27746 60786
rect 27918 60734 27970 60786
rect 28366 60734 28418 60786
rect 28926 60734 28978 60786
rect 31950 60734 32002 60786
rect 33406 60734 33458 60786
rect 34750 60734 34802 60786
rect 35870 60734 35922 60786
rect 36094 60734 36146 60786
rect 37774 60734 37826 60786
rect 39006 60734 39058 60786
rect 39902 60734 39954 60786
rect 41358 60734 41410 60786
rect 42478 60734 42530 60786
rect 48862 60734 48914 60786
rect 49310 60734 49362 60786
rect 49646 60734 49698 60786
rect 50094 60734 50146 60786
rect 51214 60734 51266 60786
rect 53006 60734 53058 60786
rect 54686 60734 54738 60786
rect 56926 60734 56978 60786
rect 57262 60734 57314 60786
rect 3502 60622 3554 60674
rect 5630 60622 5682 60674
rect 11118 60622 11170 60674
rect 13918 60622 13970 60674
rect 14254 60622 14306 60674
rect 18846 60622 18898 60674
rect 23214 60622 23266 60674
rect 28702 60622 28754 60674
rect 30046 60622 30098 60674
rect 30494 60622 30546 60674
rect 31614 60622 31666 60674
rect 33182 60622 33234 60674
rect 34078 60622 34130 60674
rect 34526 60622 34578 60674
rect 37326 60622 37378 60674
rect 37998 60622 38050 60674
rect 38558 60622 38610 60674
rect 41022 60622 41074 60674
rect 49758 60622 49810 60674
rect 53342 60622 53394 60674
rect 56030 60622 56082 60674
rect 57822 60622 57874 60674
rect 18062 60510 18114 60562
rect 25230 60510 25282 60562
rect 25566 60510 25618 60562
rect 29934 60510 29986 60562
rect 41470 60510 41522 60562
rect 42814 60510 42866 60562
rect 57150 60510 57202 60562
rect 57710 60510 57762 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 6974 60174 7026 60226
rect 17614 60174 17666 60226
rect 18958 60174 19010 60226
rect 22654 60174 22706 60226
rect 28366 60174 28418 60226
rect 32510 60174 32562 60226
rect 34414 60174 34466 60226
rect 34750 60174 34802 60226
rect 44270 60174 44322 60226
rect 11230 60062 11282 60114
rect 11790 60062 11842 60114
rect 12798 60062 12850 60114
rect 15710 60062 15762 60114
rect 17054 60062 17106 60114
rect 25454 60062 25506 60114
rect 27806 60062 27858 60114
rect 32062 60062 32114 60114
rect 34190 60062 34242 60114
rect 38670 60062 38722 60114
rect 42478 60062 42530 60114
rect 49870 60062 49922 60114
rect 54910 60062 54962 60114
rect 55246 60062 55298 60114
rect 6526 59950 6578 60002
rect 7086 59950 7138 60002
rect 7422 59950 7474 60002
rect 8430 59950 8482 60002
rect 9102 59950 9154 60002
rect 11678 59950 11730 60002
rect 12462 59950 12514 60002
rect 14142 59950 14194 60002
rect 15262 59950 15314 60002
rect 16494 59950 16546 60002
rect 16942 59950 16994 60002
rect 18846 59950 18898 60002
rect 19854 59950 19906 60002
rect 20190 59950 20242 60002
rect 23998 59950 24050 60002
rect 25902 59950 25954 60002
rect 26462 59950 26514 60002
rect 28030 59950 28082 60002
rect 29038 59950 29090 60002
rect 29374 59950 29426 60002
rect 31166 59950 31218 60002
rect 31614 59950 31666 60002
rect 32398 59950 32450 60002
rect 32846 59950 32898 60002
rect 33182 59950 33234 60002
rect 40238 59950 40290 60002
rect 41246 59950 41298 60002
rect 47070 59950 47122 60002
rect 50990 59950 51042 60002
rect 51214 59950 51266 60002
rect 51662 59950 51714 60002
rect 51886 59950 51938 60002
rect 52110 59950 52162 60002
rect 58046 59950 58098 60002
rect 12014 59838 12066 59890
rect 13806 59838 13858 59890
rect 16158 59838 16210 59890
rect 16270 59838 16322 59890
rect 22990 59838 23042 59890
rect 23326 59838 23378 59890
rect 24894 59838 24946 59890
rect 26574 59838 26626 59890
rect 29262 59838 29314 59890
rect 33070 59838 33122 59890
rect 44158 59838 44210 59890
rect 47742 59838 47794 59890
rect 50206 59838 50258 59890
rect 57374 59838 57426 59890
rect 5854 59726 5906 59778
rect 21982 59726 22034 59778
rect 22766 59726 22818 59778
rect 26014 59726 26066 59778
rect 27470 59726 27522 59778
rect 30382 59726 30434 59778
rect 30718 59726 30770 59778
rect 32510 59726 32562 59778
rect 33630 59726 33682 59778
rect 40014 59726 40066 59778
rect 40686 59726 40738 59778
rect 40798 59726 40850 59778
rect 40910 59726 40962 59778
rect 50542 59726 50594 59778
rect 51102 59726 51154 59778
rect 51998 59726 52050 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 7646 59390 7698 59442
rect 11342 59390 11394 59442
rect 15038 59390 15090 59442
rect 15150 59390 15202 59442
rect 15710 59390 15762 59442
rect 16718 59390 16770 59442
rect 27022 59390 27074 59442
rect 42254 59390 42306 59442
rect 48078 59390 48130 59442
rect 48862 59390 48914 59442
rect 48974 59390 49026 59442
rect 49534 59390 49586 59442
rect 50430 59390 50482 59442
rect 54686 59390 54738 59442
rect 56030 59390 56082 59442
rect 56702 59390 56754 59442
rect 7534 59278 7586 59330
rect 7758 59278 7810 59330
rect 8206 59278 8258 59330
rect 17614 59278 17666 59330
rect 37214 59278 37266 59330
rect 40350 59278 40402 59330
rect 40910 59278 40962 59330
rect 41470 59278 41522 59330
rect 42366 59278 42418 59330
rect 43038 59278 43090 59330
rect 48190 59278 48242 59330
rect 56590 59278 56642 59330
rect 56814 59278 56866 59330
rect 12238 59166 12290 59218
rect 14478 59166 14530 59218
rect 14926 59166 14978 59218
rect 16046 59166 16098 59218
rect 16382 59166 16434 59218
rect 17726 59166 17778 59218
rect 27246 59166 27298 59218
rect 35422 59166 35474 59218
rect 35982 59166 36034 59218
rect 39902 59166 39954 59218
rect 41246 59166 41298 59218
rect 41918 59166 41970 59218
rect 42142 59166 42194 59218
rect 42590 59166 42642 59218
rect 42926 59166 42978 59218
rect 43262 59166 43314 59218
rect 45278 59166 45330 59218
rect 45726 59166 45778 59218
rect 49310 59166 49362 59218
rect 49422 59166 49474 59218
rect 49982 59166 50034 59218
rect 51438 59166 51490 59218
rect 58158 59166 58210 59218
rect 1822 59054 1874 59106
rect 12798 59054 12850 59106
rect 18062 59054 18114 59106
rect 27806 59054 27858 59106
rect 30942 59054 30994 59106
rect 32286 59054 32338 59106
rect 36878 59054 36930 59106
rect 39454 59054 39506 59106
rect 41022 59054 41074 59106
rect 49646 59054 49698 59106
rect 52110 59054 52162 59106
rect 54238 59054 54290 59106
rect 57710 59054 57762 59106
rect 35646 58942 35698 58994
rect 44942 58942 44994 58994
rect 45278 58942 45330 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 16718 58606 16770 58658
rect 43150 58606 43202 58658
rect 52110 58606 52162 58658
rect 10222 58494 10274 58546
rect 27582 58494 27634 58546
rect 36206 58494 36258 58546
rect 39230 58494 39282 58546
rect 41358 58494 41410 58546
rect 41806 58494 41858 58546
rect 44830 58494 44882 58546
rect 46958 58494 47010 58546
rect 48190 58494 48242 58546
rect 51998 58494 52050 58546
rect 54686 58494 54738 58546
rect 58270 58494 58322 58546
rect 2270 58382 2322 58434
rect 4062 58382 4114 58434
rect 4286 58382 4338 58434
rect 11790 58382 11842 58434
rect 13806 58382 13858 58434
rect 16382 58382 16434 58434
rect 26686 58382 26738 58434
rect 27470 58382 27522 58434
rect 38558 58382 38610 58434
rect 43262 58382 43314 58434
rect 47742 58382 47794 58434
rect 53006 58382 53058 58434
rect 1710 58270 1762 58322
rect 3838 58270 3890 58322
rect 5630 58270 5682 58322
rect 10670 58270 10722 58322
rect 13470 58270 13522 58322
rect 16158 58270 16210 58322
rect 28142 58270 28194 58322
rect 29822 58270 29874 58322
rect 30494 58270 30546 58322
rect 35982 58270 36034 58322
rect 43150 58270 43202 58322
rect 3950 58158 4002 58210
rect 4846 58158 4898 58210
rect 5742 58158 5794 58210
rect 5966 58158 6018 58210
rect 12014 58158 12066 58210
rect 14478 58158 14530 58210
rect 15374 58158 15426 58210
rect 15822 58158 15874 58210
rect 26574 58158 26626 58210
rect 29934 58158 29986 58210
rect 30046 58158 30098 58210
rect 30606 58158 30658 58210
rect 30830 58158 30882 58210
rect 36206 58158 36258 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 6862 57822 6914 57874
rect 9886 57822 9938 57874
rect 10558 57822 10610 57874
rect 13806 57822 13858 57874
rect 20526 57822 20578 57874
rect 25230 57822 25282 57874
rect 44942 57822 44994 57874
rect 51662 57822 51714 57874
rect 52558 57822 52610 57874
rect 2494 57710 2546 57762
rect 4958 57710 5010 57762
rect 7982 57710 8034 57762
rect 19630 57710 19682 57762
rect 19742 57710 19794 57762
rect 22878 57710 22930 57762
rect 23998 57710 24050 57762
rect 25454 57710 25506 57762
rect 25566 57710 25618 57762
rect 25902 57710 25954 57762
rect 28254 57710 28306 57762
rect 30046 57710 30098 57762
rect 32286 57710 32338 57762
rect 36430 57710 36482 57762
rect 39006 57710 39058 57762
rect 43262 57710 43314 57762
rect 1822 57598 1874 57650
rect 5630 57598 5682 57650
rect 6302 57598 6354 57650
rect 8318 57598 8370 57650
rect 8542 57598 8594 57650
rect 9438 57598 9490 57650
rect 10110 57598 10162 57650
rect 10334 57598 10386 57650
rect 10670 57598 10722 57650
rect 13918 57598 13970 57650
rect 19406 57598 19458 57650
rect 20078 57598 20130 57650
rect 20302 57598 20354 57650
rect 20750 57598 20802 57650
rect 22766 57598 22818 57650
rect 23662 57598 23714 57650
rect 24670 57598 24722 57650
rect 26238 57598 26290 57650
rect 27022 57598 27074 57650
rect 27582 57598 27634 57650
rect 30270 57598 30322 57650
rect 30942 57598 30994 57650
rect 37662 57598 37714 57650
rect 42142 57598 42194 57650
rect 44494 57598 44546 57650
rect 51438 57598 51490 57650
rect 51998 57598 52050 57650
rect 4622 57486 4674 57538
rect 5854 57486 5906 57538
rect 8094 57486 8146 57538
rect 9998 57486 10050 57538
rect 13358 57486 13410 57538
rect 23774 57486 23826 57538
rect 31614 57486 31666 57538
rect 32062 57486 32114 57538
rect 33182 57486 33234 57538
rect 36206 57486 36258 57538
rect 42590 57486 42642 57538
rect 43150 57486 43202 57538
rect 51102 57486 51154 57538
rect 51550 57486 51602 57538
rect 6526 57374 6578 57426
rect 13806 57374 13858 57426
rect 22654 57374 22706 57426
rect 32398 57374 32450 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 12238 57038 12290 57090
rect 24670 57038 24722 57090
rect 27246 57038 27298 57090
rect 29822 57038 29874 57090
rect 43598 57038 43650 57090
rect 4398 56926 4450 56978
rect 6078 56926 6130 56978
rect 7422 56926 7474 56978
rect 9550 56926 9602 56978
rect 10670 56926 10722 56978
rect 14142 56926 14194 56978
rect 15038 56926 15090 56978
rect 16158 56926 16210 56978
rect 19406 56926 19458 56978
rect 20190 56926 20242 56978
rect 22094 56926 22146 56978
rect 24222 56926 24274 56978
rect 29934 56926 29986 56978
rect 31614 56926 31666 56978
rect 33742 56926 33794 56978
rect 34974 56926 35026 56978
rect 36318 56926 36370 56978
rect 42366 56926 42418 56978
rect 42702 56926 42754 56978
rect 47070 56926 47122 56978
rect 50430 56926 50482 56978
rect 55358 56926 55410 56978
rect 4510 56814 4562 56866
rect 4958 56814 5010 56866
rect 5518 56814 5570 56866
rect 5966 56814 6018 56866
rect 6750 56814 6802 56866
rect 10558 56814 10610 56866
rect 14590 56814 14642 56866
rect 16494 56814 16546 56866
rect 20302 56814 20354 56866
rect 20750 56814 20802 56866
rect 21310 56814 21362 56866
rect 25454 56814 25506 56866
rect 26126 56814 26178 56866
rect 26686 56814 26738 56866
rect 30158 56814 30210 56866
rect 30830 56814 30882 56866
rect 34526 56814 34578 56866
rect 35982 56814 36034 56866
rect 37102 56814 37154 56866
rect 37326 56814 37378 56866
rect 37998 56814 38050 56866
rect 42254 56814 42306 56866
rect 42926 56814 42978 56866
rect 49982 56814 50034 56866
rect 4286 56702 4338 56754
rect 9886 56702 9938 56754
rect 12014 56702 12066 56754
rect 13806 56702 13858 56754
rect 13918 56702 13970 56754
rect 14254 56702 14306 56754
rect 15150 56702 15202 56754
rect 17278 56702 17330 56754
rect 19854 56702 19906 56754
rect 24782 56702 24834 56754
rect 25118 56702 25170 56754
rect 26798 56702 26850 56754
rect 27134 56702 27186 56754
rect 36094 56702 36146 56754
rect 36430 56702 36482 56754
rect 42478 56702 42530 56754
rect 43262 56702 43314 56754
rect 43486 56702 43538 56754
rect 49198 56702 49250 56754
rect 55582 56702 55634 56754
rect 6190 56590 6242 56642
rect 12574 56590 12626 56642
rect 14030 56590 14082 56642
rect 14926 56590 14978 56642
rect 20078 56590 20130 56642
rect 24670 56590 24722 56642
rect 27694 56590 27746 56642
rect 55358 56590 55410 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 8654 56254 8706 56306
rect 8766 56254 8818 56306
rect 9774 56254 9826 56306
rect 10782 56254 10834 56306
rect 11230 56254 11282 56306
rect 12126 56254 12178 56306
rect 13694 56254 13746 56306
rect 14590 56254 14642 56306
rect 22654 56254 22706 56306
rect 28478 56254 28530 56306
rect 46958 56254 47010 56306
rect 48190 56254 48242 56306
rect 48862 56254 48914 56306
rect 49982 56254 50034 56306
rect 54238 56254 54290 56306
rect 8318 56142 8370 56194
rect 12910 56142 12962 56194
rect 13134 56142 13186 56194
rect 13358 56142 13410 56194
rect 13470 56142 13522 56194
rect 13918 56142 13970 56194
rect 14030 56142 14082 56194
rect 17950 56142 18002 56194
rect 19070 56142 19122 56194
rect 20302 56142 20354 56194
rect 23886 56142 23938 56194
rect 31838 56142 31890 56194
rect 32510 56142 32562 56194
rect 35198 56142 35250 56194
rect 35646 56142 35698 56194
rect 37326 56142 37378 56194
rect 48750 56142 48802 56194
rect 51662 56142 51714 56194
rect 8542 56030 8594 56082
rect 10222 56030 10274 56082
rect 10446 56030 10498 56082
rect 11566 56030 11618 56082
rect 12462 56030 12514 56082
rect 12798 56030 12850 56082
rect 14254 56030 14306 56082
rect 15150 56030 15202 56082
rect 22990 56030 23042 56082
rect 32286 56030 32338 56082
rect 33630 56030 33682 56082
rect 34190 56030 34242 56082
rect 35870 56030 35922 56082
rect 37214 56030 37266 56082
rect 38222 56030 38274 56082
rect 39006 56030 39058 56082
rect 47070 56030 47122 56082
rect 47182 56030 47234 56082
rect 47630 56030 47682 56082
rect 48078 56030 48130 56082
rect 50318 56030 50370 56082
rect 50878 56030 50930 56082
rect 54910 56030 54962 56082
rect 4510 55918 4562 55970
rect 5070 55918 5122 55970
rect 15262 55918 15314 55970
rect 17838 55918 17890 55970
rect 18174 55918 18226 55970
rect 18734 55918 18786 55970
rect 20750 55918 20802 55970
rect 24446 55918 24498 55970
rect 25342 55918 25394 55970
rect 31390 55918 31442 55970
rect 45502 55918 45554 55970
rect 47854 55918 47906 55970
rect 53790 55918 53842 55970
rect 55134 55918 55186 55970
rect 15934 55806 15986 55858
rect 45614 55806 45666 55858
rect 55582 55806 55634 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 4734 55470 4786 55522
rect 23550 55470 23602 55522
rect 32286 55470 32338 55522
rect 35198 55470 35250 55522
rect 43150 55470 43202 55522
rect 11790 55358 11842 55410
rect 23774 55358 23826 55410
rect 33182 55358 33234 55410
rect 34862 55358 34914 55410
rect 40462 55358 40514 55410
rect 41582 55358 41634 55410
rect 42142 55358 42194 55410
rect 45614 55358 45666 55410
rect 47742 55358 47794 55410
rect 52782 55358 52834 55410
rect 55582 55358 55634 55410
rect 57710 55358 57762 55410
rect 3390 55246 3442 55298
rect 3838 55246 3890 55298
rect 4398 55246 4450 55298
rect 11006 55246 11058 55298
rect 11342 55246 11394 55298
rect 14478 55246 14530 55298
rect 23886 55246 23938 55298
rect 28366 55246 28418 55298
rect 29262 55246 29314 55298
rect 30158 55246 30210 55298
rect 31726 55246 31778 55298
rect 32958 55246 33010 55298
rect 33854 55246 33906 55298
rect 34750 55246 34802 55298
rect 37662 55246 37714 55298
rect 41470 55246 41522 55298
rect 42366 55246 42418 55298
rect 42814 55246 42866 55298
rect 44942 55246 44994 55298
rect 53342 55246 53394 55298
rect 54910 55246 54962 55298
rect 58158 55246 58210 55298
rect 2830 55134 2882 55186
rect 3166 55134 3218 55186
rect 4846 55134 4898 55186
rect 29374 55134 29426 55186
rect 30718 55134 30770 55186
rect 31390 55134 31442 55186
rect 31502 55134 31554 55186
rect 32286 55134 32338 55186
rect 32398 55134 32450 55186
rect 38334 55134 38386 55186
rect 40798 55134 40850 55186
rect 49982 55134 50034 55186
rect 2942 55022 2994 55074
rect 3726 55022 3778 55074
rect 3950 55022 4002 55074
rect 4734 55022 4786 55074
rect 11118 55022 11170 55074
rect 12686 55022 12738 55074
rect 13582 55022 13634 55074
rect 14590 55022 14642 55074
rect 18398 55022 18450 55074
rect 27694 55022 27746 55074
rect 27806 55022 27858 55074
rect 27918 55022 27970 55074
rect 30158 55022 30210 55074
rect 31054 55022 31106 55074
rect 43038 55022 43090 55074
rect 44270 55022 44322 55074
rect 49198 55022 49250 55074
rect 49534 55022 49586 55074
rect 50318 55022 50370 55074
rect 52782 55022 52834 55074
rect 52894 55022 52946 55074
rect 53118 55022 53170 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 5070 54686 5122 54738
rect 11006 54686 11058 54738
rect 14590 54686 14642 54738
rect 29486 54686 29538 54738
rect 39566 54686 39618 54738
rect 41022 54686 41074 54738
rect 41582 54686 41634 54738
rect 41694 54686 41746 54738
rect 41806 54686 41858 54738
rect 42478 54686 42530 54738
rect 45502 54686 45554 54738
rect 45950 54686 46002 54738
rect 46622 54686 46674 54738
rect 51886 54686 51938 54738
rect 2494 54574 2546 54626
rect 5406 54574 5458 54626
rect 26686 54574 26738 54626
rect 27022 54574 27074 54626
rect 31502 54574 31554 54626
rect 39454 54574 39506 54626
rect 39790 54574 39842 54626
rect 42366 54574 42418 54626
rect 51214 54574 51266 54626
rect 55806 54574 55858 54626
rect 1822 54462 1874 54514
rect 4958 54462 5010 54514
rect 5182 54462 5234 54514
rect 11342 54462 11394 54514
rect 14254 54462 14306 54514
rect 14478 54462 14530 54514
rect 14814 54462 14866 54514
rect 15150 54462 15202 54514
rect 15374 54462 15426 54514
rect 18286 54462 18338 54514
rect 27246 54462 27298 54514
rect 27582 54462 27634 54514
rect 28142 54462 28194 54514
rect 31054 54462 31106 54514
rect 39902 54462 39954 54514
rect 41470 54462 41522 54514
rect 42030 54462 42082 54514
rect 46062 54462 46114 54514
rect 46398 54462 46450 54514
rect 46622 54462 46674 54514
rect 50878 54462 50930 54514
rect 51662 54462 51714 54514
rect 56478 54462 56530 54514
rect 56814 54462 56866 54514
rect 57150 54462 57202 54514
rect 4622 54350 4674 54402
rect 16046 54350 16098 54402
rect 26798 54350 26850 54402
rect 28478 54350 28530 54402
rect 28926 54350 28978 54402
rect 29150 54350 29202 54402
rect 30606 54350 30658 54402
rect 31950 54350 32002 54402
rect 32510 54350 32562 54402
rect 33182 54350 33234 54402
rect 46846 54350 46898 54402
rect 47182 54350 47234 54402
rect 55134 54350 55186 54402
rect 55918 54350 55970 54402
rect 56702 54350 56754 54402
rect 54574 54238 54626 54290
rect 54910 54238 54962 54290
rect 56030 54238 56082 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 8990 53902 9042 53954
rect 23326 53902 23378 53954
rect 29374 53902 29426 53954
rect 29710 53902 29762 53954
rect 36318 53902 36370 53954
rect 52670 53902 52722 53954
rect 2942 53790 2994 53842
rect 5070 53790 5122 53842
rect 18734 53790 18786 53842
rect 22318 53790 22370 53842
rect 24110 53790 24162 53842
rect 26014 53790 26066 53842
rect 28142 53790 28194 53842
rect 29150 53790 29202 53842
rect 36094 53790 36146 53842
rect 37102 53790 37154 53842
rect 39902 53790 39954 53842
rect 53006 53790 53058 53842
rect 53902 53790 53954 53842
rect 56030 53790 56082 53842
rect 58158 53790 58210 53842
rect 3390 53678 3442 53730
rect 3838 53678 3890 53730
rect 4622 53678 4674 53730
rect 8430 53678 8482 53730
rect 8878 53678 8930 53730
rect 17838 53678 17890 53730
rect 18398 53678 18450 53730
rect 19854 53678 19906 53730
rect 19966 53678 20018 53730
rect 23886 53678 23938 53730
rect 24782 53678 24834 53730
rect 25342 53678 25394 53730
rect 34526 53678 34578 53730
rect 35982 53678 36034 53730
rect 37326 53678 37378 53730
rect 37998 53678 38050 53730
rect 39790 53678 39842 53730
rect 40014 53678 40066 53730
rect 51438 53678 51490 53730
rect 54910 53678 54962 53730
rect 55246 53678 55298 53730
rect 4286 53566 4338 53618
rect 4398 53566 4450 53618
rect 7086 53566 7138 53618
rect 7422 53566 7474 53618
rect 7646 53566 7698 53618
rect 10334 53566 10386 53618
rect 17950 53566 18002 53618
rect 19070 53566 19122 53618
rect 20638 53566 20690 53618
rect 22654 53566 22706 53618
rect 23102 53566 23154 53618
rect 24334 53566 24386 53618
rect 30382 53566 30434 53618
rect 40238 53566 40290 53618
rect 40910 53566 40962 53618
rect 41246 53566 41298 53618
rect 41582 53566 41634 53618
rect 41694 53566 41746 53618
rect 54238 53566 54290 53618
rect 54798 53566 54850 53618
rect 7198 53454 7250 53506
rect 8094 53454 8146 53506
rect 8318 53454 8370 53506
rect 8542 53454 8594 53506
rect 8990 53454 9042 53506
rect 10670 53454 10722 53506
rect 18174 53454 18226 53506
rect 18622 53454 18674 53506
rect 18846 53454 18898 53506
rect 19630 53454 19682 53506
rect 20078 53454 20130 53506
rect 20302 53454 20354 53506
rect 20526 53454 20578 53506
rect 22430 53454 22482 53506
rect 23214 53454 23266 53506
rect 30046 53454 30098 53506
rect 33182 53454 33234 53506
rect 39566 53454 39618 53506
rect 41022 53454 41074 53506
rect 41358 53454 41410 53506
rect 51662 53454 51714 53506
rect 52782 53454 52834 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 8542 53118 8594 53170
rect 13134 53118 13186 53170
rect 14590 53118 14642 53170
rect 23998 53118 24050 53170
rect 24670 53118 24722 53170
rect 25342 53118 25394 53170
rect 31278 53118 31330 53170
rect 36430 53118 36482 53170
rect 41022 53118 41074 53170
rect 45838 53118 45890 53170
rect 46622 53118 46674 53170
rect 46846 53118 46898 53170
rect 47518 53118 47570 53170
rect 47966 53118 48018 53170
rect 55022 53118 55074 53170
rect 5966 53006 6018 53058
rect 12014 53006 12066 53058
rect 12574 53006 12626 53058
rect 14814 53006 14866 53058
rect 18174 53006 18226 53058
rect 21422 53006 21474 53058
rect 23886 53006 23938 53058
rect 36206 53006 36258 53058
rect 36654 53006 36706 53058
rect 51550 53006 51602 53058
rect 5294 52894 5346 52946
rect 8430 52894 8482 52946
rect 8654 52894 8706 52946
rect 9102 52894 9154 52946
rect 11566 52894 11618 52946
rect 12350 52894 12402 52946
rect 12686 52894 12738 52946
rect 14926 52894 14978 52946
rect 17502 52894 17554 52946
rect 20638 52894 20690 52946
rect 24222 52894 24274 52946
rect 31502 52894 31554 52946
rect 32174 52894 32226 52946
rect 33742 52894 33794 52946
rect 34414 52894 34466 52946
rect 35646 52894 35698 52946
rect 35982 52894 36034 52946
rect 36766 52894 36818 52946
rect 42478 52894 42530 52946
rect 46398 52894 46450 52946
rect 47070 52894 47122 52946
rect 50766 52894 50818 52946
rect 54126 52894 54178 52946
rect 54462 52894 54514 52946
rect 58158 52894 58210 52946
rect 8094 52782 8146 52834
rect 9774 52782 9826 52834
rect 10110 52782 10162 52834
rect 10670 52782 10722 52834
rect 11118 52782 11170 52834
rect 13694 52782 13746 52834
rect 20302 52782 20354 52834
rect 23550 52782 23602 52834
rect 31950 52782 32002 52834
rect 33518 52782 33570 52834
rect 43262 52782 43314 52834
rect 45390 52782 45442 52834
rect 46510 52782 46562 52834
rect 53678 52782 53730 52834
rect 57374 52782 57426 52834
rect 57598 52782 57650 52834
rect 10334 52670 10386 52722
rect 32510 52670 32562 52722
rect 45614 52670 45666 52722
rect 46174 52670 46226 52722
rect 47294 52670 47346 52722
rect 47630 52670 47682 52722
rect 54014 52670 54066 52722
rect 54350 52670 54402 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 8766 52334 8818 52386
rect 15710 52334 15762 52386
rect 16158 52334 16210 52386
rect 16494 52334 16546 52386
rect 20414 52334 20466 52386
rect 36094 52334 36146 52386
rect 55918 52334 55970 52386
rect 56142 52334 56194 52386
rect 56254 52334 56306 52386
rect 4622 52222 4674 52274
rect 7310 52222 7362 52274
rect 8206 52222 8258 52274
rect 12350 52222 12402 52274
rect 13694 52222 13746 52274
rect 18510 52222 18562 52274
rect 19406 52222 19458 52274
rect 20190 52222 20242 52274
rect 20750 52222 20802 52274
rect 21534 52222 21586 52274
rect 24558 52222 24610 52274
rect 32398 52222 32450 52274
rect 33630 52222 33682 52274
rect 35982 52222 36034 52274
rect 39454 52222 39506 52274
rect 43262 52222 43314 52274
rect 46734 52222 46786 52274
rect 47630 52222 47682 52274
rect 51214 52222 51266 52274
rect 51774 52222 51826 52274
rect 7982 52110 8034 52162
rect 8654 52110 8706 52162
rect 10334 52110 10386 52162
rect 10782 52110 10834 52162
rect 12910 52110 12962 52162
rect 13806 52110 13858 52162
rect 14478 52110 14530 52162
rect 14814 52110 14866 52162
rect 15038 52110 15090 52162
rect 15262 52110 15314 52162
rect 15934 52110 15986 52162
rect 19182 52110 19234 52162
rect 23102 52110 23154 52162
rect 30942 52110 30994 52162
rect 31502 52110 31554 52162
rect 31838 52110 31890 52162
rect 32734 52110 32786 52162
rect 33294 52110 33346 52162
rect 35646 52110 35698 52162
rect 38894 52110 38946 52162
rect 43822 52110 43874 52162
rect 46622 52110 46674 52162
rect 50542 52110 50594 52162
rect 50990 52110 51042 52162
rect 54126 52110 54178 52162
rect 8766 51998 8818 52050
rect 9998 51998 10050 52050
rect 11454 51998 11506 52050
rect 24334 51998 24386 52050
rect 30718 51998 30770 52050
rect 33742 51998 33794 52050
rect 43150 51998 43202 52050
rect 44158 51998 44210 52050
rect 47070 51998 47122 52050
rect 47294 51998 47346 52050
rect 49758 51998 49810 52050
rect 11790 51886 11842 51938
rect 12238 51886 12290 51938
rect 12462 51886 12514 51938
rect 22542 51886 22594 51938
rect 43374 51886 43426 51938
rect 46846 51886 46898 51938
rect 54462 51886 54514 51938
rect 56254 51886 56306 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 3950 51550 4002 51602
rect 12798 51550 12850 51602
rect 13022 51550 13074 51602
rect 13246 51550 13298 51602
rect 15150 51550 15202 51602
rect 32510 51550 32562 51602
rect 36318 51550 36370 51602
rect 43262 51550 43314 51602
rect 47182 51550 47234 51602
rect 48302 51550 48354 51602
rect 48862 51550 48914 51602
rect 51886 51550 51938 51602
rect 52782 51550 52834 51602
rect 55918 51550 55970 51602
rect 56702 51550 56754 51602
rect 3390 51438 3442 51490
rect 5406 51438 5458 51490
rect 37326 51438 37378 51490
rect 38670 51438 38722 51490
rect 41022 51438 41074 51490
rect 41694 51438 41746 51490
rect 48750 51438 48802 51490
rect 53230 51438 53282 51490
rect 55470 51438 55522 51490
rect 3278 51326 3330 51378
rect 3614 51326 3666 51378
rect 4174 51326 4226 51378
rect 4398 51326 4450 51378
rect 5070 51326 5122 51378
rect 5742 51326 5794 51378
rect 13358 51326 13410 51378
rect 14590 51326 14642 51378
rect 15038 51326 15090 51378
rect 15262 51326 15314 51378
rect 28366 51326 28418 51378
rect 28478 51326 28530 51378
rect 29150 51326 29202 51378
rect 30158 51326 30210 51378
rect 36206 51326 36258 51378
rect 36766 51326 36818 51378
rect 37998 51326 38050 51378
rect 41582 51326 41634 51378
rect 43710 51326 43762 51378
rect 46958 51326 47010 51378
rect 47294 51326 47346 51378
rect 47630 51326 47682 51378
rect 52110 51326 52162 51378
rect 52446 51326 52498 51378
rect 55134 51326 55186 51378
rect 55358 51326 55410 51378
rect 56478 51326 56530 51378
rect 56814 51326 56866 51378
rect 57038 51326 57090 51378
rect 4286 51214 4338 51266
rect 5518 51214 5570 51266
rect 29038 51214 29090 51266
rect 29822 51214 29874 51266
rect 37774 51214 37826 51266
rect 42254 51214 42306 51266
rect 44382 51214 44434 51266
rect 46510 51214 46562 51266
rect 47854 51214 47906 51266
rect 48190 51214 48242 51266
rect 40910 51102 40962 51154
rect 41246 51102 41298 51154
rect 41694 51102 41746 51154
rect 51774 51102 51826 51154
rect 53118 51102 53170 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 5070 50766 5122 50818
rect 5742 50766 5794 50818
rect 14366 50766 14418 50818
rect 33406 50766 33458 50818
rect 28366 50710 28418 50762
rect 41806 50766 41858 50818
rect 4622 50654 4674 50706
rect 9326 50654 9378 50706
rect 11678 50654 11730 50706
rect 35198 50654 35250 50706
rect 36318 50654 36370 50706
rect 38558 50654 38610 50706
rect 40686 50654 40738 50706
rect 44942 50654 44994 50706
rect 56030 50654 56082 50706
rect 58158 50654 58210 50706
rect 1822 50542 1874 50594
rect 4958 50542 5010 50594
rect 5630 50542 5682 50594
rect 9102 50542 9154 50594
rect 9774 50542 9826 50594
rect 14030 50542 14082 50594
rect 25454 50542 25506 50594
rect 29262 50542 29314 50594
rect 29486 50542 29538 50594
rect 30158 50542 30210 50594
rect 30382 50542 30434 50594
rect 30942 50542 30994 50594
rect 32286 50542 32338 50594
rect 32510 50542 32562 50594
rect 33294 50542 33346 50594
rect 35086 50542 35138 50594
rect 41470 50542 41522 50594
rect 41918 50542 41970 50594
rect 42142 50542 42194 50594
rect 42254 50542 42306 50594
rect 42814 50542 42866 50594
rect 44830 50542 44882 50594
rect 45502 50542 45554 50594
rect 45838 50542 45890 50594
rect 46734 50542 46786 50594
rect 47182 50542 47234 50594
rect 47406 50542 47458 50594
rect 55246 50542 55298 50594
rect 2494 50430 2546 50482
rect 5742 50430 5794 50482
rect 8766 50430 8818 50482
rect 10782 50430 10834 50482
rect 11118 50430 11170 50482
rect 19630 50430 19682 50482
rect 25118 50430 25170 50482
rect 26238 50430 26290 50482
rect 30606 50430 30658 50482
rect 30830 50430 30882 50482
rect 47854 50430 47906 50482
rect 13694 50318 13746 50370
rect 14254 50318 14306 50370
rect 19742 50318 19794 50370
rect 45054 50318 45106 50370
rect 46958 50318 47010 50370
rect 47070 50318 47122 50370
rect 54910 50318 54962 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4510 49982 4562 50034
rect 9438 49982 9490 50034
rect 12350 49982 12402 50034
rect 28478 49982 28530 50034
rect 28702 49982 28754 50034
rect 29374 49982 29426 50034
rect 29486 49982 29538 50034
rect 30158 49982 30210 50034
rect 35422 49982 35474 50034
rect 41022 49982 41074 50034
rect 41358 49982 41410 50034
rect 51102 49982 51154 50034
rect 4062 49870 4114 49922
rect 9662 49870 9714 49922
rect 10222 49870 10274 49922
rect 19294 49870 19346 49922
rect 20302 49870 20354 49922
rect 21534 49870 21586 49922
rect 28366 49870 28418 49922
rect 29038 49870 29090 49922
rect 29822 49870 29874 49922
rect 29934 49870 29986 49922
rect 34078 49870 34130 49922
rect 37662 49870 37714 49922
rect 39342 49870 39394 49922
rect 41918 49870 41970 49922
rect 47294 49870 47346 49922
rect 50878 49870 50930 49922
rect 51662 49870 51714 49922
rect 51998 49870 52050 49922
rect 52222 49870 52274 49922
rect 3390 49758 3442 49810
rect 3950 49758 4002 49810
rect 4286 49758 4338 49810
rect 4734 49758 4786 49810
rect 4846 49758 4898 49810
rect 8654 49758 8706 49810
rect 8878 49758 8930 49810
rect 9774 49758 9826 49810
rect 9998 49758 10050 49810
rect 10334 49758 10386 49810
rect 12686 49758 12738 49810
rect 13246 49758 13298 49810
rect 14254 49758 14306 49810
rect 19182 49758 19234 49810
rect 19518 49758 19570 49810
rect 20190 49758 20242 49810
rect 21198 49758 21250 49810
rect 21422 49758 21474 49810
rect 23774 49758 23826 49810
rect 29262 49758 29314 49810
rect 31614 49758 31666 49810
rect 32062 49758 32114 49810
rect 33406 49758 33458 49810
rect 35086 49758 35138 49810
rect 38670 49758 38722 49810
rect 41246 49758 41298 49810
rect 41470 49758 41522 49810
rect 50766 49758 50818 49810
rect 52670 49758 52722 49810
rect 5406 49646 5458 49698
rect 7982 49646 8034 49698
rect 14030 49646 14082 49698
rect 20526 49646 20578 49698
rect 23662 49646 23714 49698
rect 30494 49646 30546 49698
rect 31054 49646 31106 49698
rect 32398 49646 32450 49698
rect 33182 49646 33234 49698
rect 34862 49646 34914 49698
rect 37214 49646 37266 49698
rect 41806 49646 41858 49698
rect 42142 49646 42194 49698
rect 49870 49646 49922 49698
rect 50430 49646 50482 49698
rect 52446 49646 52498 49698
rect 14702 49534 14754 49586
rect 21534 49534 21586 49586
rect 23438 49534 23490 49586
rect 47406 49534 47458 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 32958 49198 33010 49250
rect 33294 49198 33346 49250
rect 53006 49198 53058 49250
rect 8878 49086 8930 49138
rect 10222 49086 10274 49138
rect 15822 49086 15874 49138
rect 16270 49086 16322 49138
rect 17390 49086 17442 49138
rect 19518 49086 19570 49138
rect 20078 49086 20130 49138
rect 23662 49086 23714 49138
rect 25790 49086 25842 49138
rect 32734 49086 32786 49138
rect 33742 49086 33794 49138
rect 42142 49086 42194 49138
rect 46734 49086 46786 49138
rect 48862 49086 48914 49138
rect 58158 49086 58210 49138
rect 6078 48974 6130 49026
rect 9102 48974 9154 49026
rect 9662 48974 9714 49026
rect 15598 48974 15650 49026
rect 16718 48974 16770 49026
rect 21982 48974 22034 49026
rect 22542 48974 22594 49026
rect 22990 48974 23042 49026
rect 31726 48974 31778 49026
rect 32174 48974 32226 49026
rect 32398 48974 32450 49026
rect 41918 48974 41970 49026
rect 42030 48974 42082 49026
rect 42254 48974 42306 49026
rect 42814 48974 42866 49026
rect 49646 48974 49698 49026
rect 50878 48974 50930 49026
rect 51102 48974 51154 49026
rect 51550 48974 51602 49026
rect 52782 48974 52834 49026
rect 53230 48974 53282 49026
rect 54126 48974 54178 49026
rect 54462 48974 54514 49026
rect 54910 48974 54962 49026
rect 55246 48974 55298 49026
rect 6750 48862 6802 48914
rect 9326 48862 9378 48914
rect 9550 48862 9602 48914
rect 11118 48862 11170 48914
rect 19966 48862 20018 48914
rect 20302 48862 20354 48914
rect 20526 48862 20578 48914
rect 21422 48862 21474 48914
rect 43150 48862 43202 48914
rect 54686 48862 54738 48914
rect 56030 48862 56082 48914
rect 11230 48750 11282 48802
rect 11342 48750 11394 48802
rect 21310 48750 21362 48802
rect 21534 48750 21586 48802
rect 42366 48750 42418 48802
rect 43038 48750 43090 48802
rect 50990 48750 51042 48802
rect 52110 48750 52162 48802
rect 53118 48750 53170 48802
rect 53902 48750 53954 48802
rect 54798 48750 54850 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 8318 48414 8370 48466
rect 8430 48414 8482 48466
rect 8542 48414 8594 48466
rect 8990 48414 9042 48466
rect 19070 48414 19122 48466
rect 20974 48414 21026 48466
rect 22094 48414 22146 48466
rect 24446 48414 24498 48466
rect 27358 48414 27410 48466
rect 32510 48414 32562 48466
rect 41694 48414 41746 48466
rect 42478 48414 42530 48466
rect 55918 48414 55970 48466
rect 4846 48302 4898 48354
rect 5854 48302 5906 48354
rect 6078 48302 6130 48354
rect 8094 48302 8146 48354
rect 8878 48302 8930 48354
rect 10558 48302 10610 48354
rect 13918 48302 13970 48354
rect 14590 48302 14642 48354
rect 15262 48302 15314 48354
rect 20414 48302 20466 48354
rect 23550 48302 23602 48354
rect 37214 48302 37266 48354
rect 42366 48302 42418 48354
rect 43374 48302 43426 48354
rect 53006 48302 53058 48354
rect 55470 48302 55522 48354
rect 55694 48302 55746 48354
rect 4622 48190 4674 48242
rect 5518 48190 5570 48242
rect 6190 48190 6242 48242
rect 11118 48190 11170 48242
rect 11790 48190 11842 48242
rect 14030 48190 14082 48242
rect 14926 48190 14978 48242
rect 15486 48190 15538 48242
rect 19518 48190 19570 48242
rect 19966 48190 20018 48242
rect 22430 48190 22482 48242
rect 27246 48190 27298 48242
rect 27470 48190 27522 48242
rect 27918 48190 27970 48242
rect 35982 48190 36034 48242
rect 37102 48190 37154 48242
rect 43262 48190 43314 48242
rect 43486 48190 43538 48242
rect 43934 48190 43986 48242
rect 49198 48190 49250 48242
rect 50094 48190 50146 48242
rect 53678 48190 53730 48242
rect 54238 48190 54290 48242
rect 54910 48190 54962 48242
rect 56142 48190 56194 48242
rect 4958 48078 5010 48130
rect 12462 48078 12514 48130
rect 13022 48078 13074 48130
rect 14142 48078 14194 48130
rect 15374 48078 15426 48130
rect 23886 48078 23938 48130
rect 24670 48078 24722 48130
rect 36654 48078 36706 48130
rect 41582 48078 41634 48130
rect 48862 48078 48914 48130
rect 49646 48078 49698 48130
rect 50878 48078 50930 48130
rect 24334 47966 24386 48018
rect 42478 47966 42530 48018
rect 50206 47966 50258 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 5630 47630 5682 47682
rect 11118 47630 11170 47682
rect 12462 47630 12514 47682
rect 22654 47630 22706 47682
rect 28366 47630 28418 47682
rect 35422 47630 35474 47682
rect 4622 47518 4674 47570
rect 5070 47518 5122 47570
rect 11230 47518 11282 47570
rect 15486 47518 15538 47570
rect 17502 47518 17554 47570
rect 23102 47518 23154 47570
rect 25902 47518 25954 47570
rect 29710 47518 29762 47570
rect 34638 47518 34690 47570
rect 37438 47518 37490 47570
rect 37998 47518 38050 47570
rect 44270 47518 44322 47570
rect 47742 47518 47794 47570
rect 56254 47518 56306 47570
rect 1822 47406 1874 47458
rect 11118 47406 11170 47458
rect 12238 47406 12290 47458
rect 12574 47406 12626 47458
rect 15934 47406 15986 47458
rect 17838 47406 17890 47458
rect 22878 47406 22930 47458
rect 23662 47406 23714 47458
rect 24558 47406 24610 47458
rect 24894 47406 24946 47458
rect 27358 47406 27410 47458
rect 27918 47406 27970 47458
rect 34750 47406 34802 47458
rect 37662 47406 37714 47458
rect 38446 47406 38498 47458
rect 39006 47406 39058 47458
rect 41694 47406 41746 47458
rect 42478 47406 42530 47458
rect 44830 47406 44882 47458
rect 52670 47406 52722 47458
rect 2494 47294 2546 47346
rect 5742 47294 5794 47346
rect 5966 47294 6018 47346
rect 13806 47294 13858 47346
rect 15038 47294 15090 47346
rect 15374 47294 15426 47346
rect 15710 47294 15762 47346
rect 18286 47294 18338 47346
rect 23998 47294 24050 47346
rect 24782 47294 24834 47346
rect 26126 47294 26178 47346
rect 28254 47294 28306 47346
rect 29374 47294 29426 47346
rect 39118 47294 39170 47346
rect 42590 47294 42642 47346
rect 45614 47294 45666 47346
rect 53454 47294 53506 47346
rect 12686 47182 12738 47234
rect 14142 47182 14194 47234
rect 14702 47182 14754 47234
rect 24334 47182 24386 47234
rect 25454 47182 25506 47234
rect 28366 47182 28418 47234
rect 29598 47182 29650 47234
rect 38558 47182 38610 47234
rect 41134 47182 41186 47234
rect 48526 47182 48578 47234
rect 49758 47182 49810 47234
rect 55694 47182 55746 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 2606 46846 2658 46898
rect 12574 46846 12626 46898
rect 13358 46846 13410 46898
rect 13694 46846 13746 46898
rect 24558 46846 24610 46898
rect 27246 46846 27298 46898
rect 35310 46846 35362 46898
rect 36094 46846 36146 46898
rect 36430 46846 36482 46898
rect 45950 46846 46002 46898
rect 53566 46846 53618 46898
rect 2494 46734 2546 46786
rect 5294 46734 5346 46786
rect 8878 46734 8930 46786
rect 12798 46734 12850 46786
rect 12910 46734 12962 46786
rect 23662 46734 23714 46786
rect 28590 46734 28642 46786
rect 28702 46734 28754 46786
rect 29822 46734 29874 46786
rect 31054 46734 31106 46786
rect 31950 46734 32002 46786
rect 34750 46734 34802 46786
rect 35870 46734 35922 46786
rect 37438 46734 37490 46786
rect 39902 46734 39954 46786
rect 41022 46734 41074 46786
rect 41246 46734 41298 46786
rect 46174 46734 46226 46786
rect 48750 46734 48802 46786
rect 4062 46622 4114 46674
rect 8766 46622 8818 46674
rect 9102 46622 9154 46674
rect 12350 46622 12402 46674
rect 14030 46622 14082 46674
rect 14702 46622 14754 46674
rect 17838 46622 17890 46674
rect 19406 46622 19458 46674
rect 23550 46622 23602 46674
rect 24446 46622 24498 46674
rect 26014 46622 26066 46674
rect 27470 46622 27522 46674
rect 28926 46622 28978 46674
rect 34974 46622 35026 46674
rect 35758 46622 35810 46674
rect 36654 46622 36706 46674
rect 38894 46622 38946 46674
rect 44494 46622 44546 46674
rect 44830 46622 44882 46674
rect 45390 46622 45442 46674
rect 45726 46622 45778 46674
rect 48078 46622 48130 46674
rect 49310 46622 49362 46674
rect 49758 46622 49810 46674
rect 50542 46622 50594 46674
rect 53342 46622 53394 46674
rect 53678 46622 53730 46674
rect 54126 46622 54178 46674
rect 55022 46622 55074 46674
rect 2718 46510 2770 46562
rect 3390 46510 3442 46562
rect 5406 46510 5458 46562
rect 10110 46510 10162 46562
rect 14926 46510 14978 46562
rect 15374 46510 15426 46562
rect 17726 46510 17778 46562
rect 26238 46510 26290 46562
rect 26798 46510 26850 46562
rect 29374 46510 29426 46562
rect 31390 46510 31442 46562
rect 31726 46510 31778 46562
rect 32510 46510 32562 46562
rect 37102 46510 37154 46562
rect 41694 46510 41746 46562
rect 45838 46510 45890 46562
rect 47630 46510 47682 46562
rect 50206 46510 50258 46562
rect 51102 46510 51154 46562
rect 53006 46510 53058 46562
rect 54798 46510 54850 46562
rect 19742 46398 19794 46450
rect 32062 46398 32114 46450
rect 36318 46398 36370 46450
rect 40910 46398 40962 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 9662 46062 9714 46114
rect 27582 46062 27634 46114
rect 29262 46062 29314 46114
rect 2942 45950 2994 46002
rect 9102 45950 9154 46002
rect 9998 45950 10050 46002
rect 12126 45950 12178 46002
rect 17726 45950 17778 46002
rect 20190 45950 20242 46002
rect 30046 45950 30098 46002
rect 31054 45950 31106 46002
rect 39566 45950 39618 46002
rect 41694 45950 41746 46002
rect 42142 45950 42194 46002
rect 50878 45950 50930 46002
rect 55246 45950 55298 46002
rect 8094 45838 8146 45890
rect 9326 45838 9378 45890
rect 12798 45838 12850 45890
rect 15038 45838 15090 45890
rect 15822 45838 15874 45890
rect 17054 45838 17106 45890
rect 17838 45838 17890 45890
rect 27246 45838 27298 45890
rect 27918 45838 27970 45890
rect 29038 45838 29090 45890
rect 30158 45838 30210 45890
rect 33966 45838 34018 45890
rect 37550 45838 37602 45890
rect 37998 45838 38050 45890
rect 38894 45838 38946 45890
rect 45054 45838 45106 45890
rect 45278 45838 45330 45890
rect 45502 45838 45554 45890
rect 48414 45838 48466 45890
rect 49310 45838 49362 45890
rect 54910 45838 54962 45890
rect 58046 45838 58098 45890
rect 14814 45726 14866 45778
rect 15486 45726 15538 45778
rect 18398 45726 18450 45778
rect 33182 45726 33234 45778
rect 49534 45726 49586 45778
rect 49982 45726 50034 45778
rect 51214 45726 51266 45778
rect 57374 45726 57426 45778
rect 7982 45614 8034 45666
rect 8206 45614 8258 45666
rect 8430 45614 8482 45666
rect 13582 45614 13634 45666
rect 15598 45614 15650 45666
rect 20750 45614 20802 45666
rect 21422 45614 21474 45666
rect 23102 45614 23154 45666
rect 28590 45614 28642 45666
rect 34414 45614 34466 45666
rect 45390 45614 45442 45666
rect 45950 45614 46002 45666
rect 48078 45614 48130 45666
rect 50654 45614 50706 45666
rect 50990 45614 51042 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 3054 45278 3106 45330
rect 9662 45278 9714 45330
rect 9774 45278 9826 45330
rect 22318 45278 22370 45330
rect 23662 45278 23714 45330
rect 24110 45278 24162 45330
rect 28702 45278 28754 45330
rect 36654 45278 36706 45330
rect 38446 45278 38498 45330
rect 48302 45278 48354 45330
rect 48750 45278 48802 45330
rect 53342 45278 53394 45330
rect 55918 45278 55970 45330
rect 58158 45278 58210 45330
rect 4958 45166 5010 45218
rect 14590 45166 14642 45218
rect 15598 45166 15650 45218
rect 21758 45166 21810 45218
rect 22206 45166 22258 45218
rect 25230 45166 25282 45218
rect 31502 45166 31554 45218
rect 49086 45166 49138 45218
rect 50766 45166 50818 45218
rect 55134 45166 55186 45218
rect 57150 45166 57202 45218
rect 5070 45054 5122 45106
rect 6078 45054 6130 45106
rect 9550 45054 9602 45106
rect 10110 45054 10162 45106
rect 14926 45054 14978 45106
rect 15822 45054 15874 45106
rect 21646 45054 21698 45106
rect 21982 45054 22034 45106
rect 22430 45054 22482 45106
rect 22878 45054 22930 45106
rect 23326 45054 23378 45106
rect 25342 45054 25394 45106
rect 25790 45054 25842 45106
rect 28478 45054 28530 45106
rect 31726 45054 31778 45106
rect 32510 45054 32562 45106
rect 36206 45054 36258 45106
rect 43822 45054 43874 45106
rect 49982 45054 50034 45106
rect 55470 45054 55522 45106
rect 55694 45054 55746 45106
rect 56030 45054 56082 45106
rect 56590 45054 56642 45106
rect 56814 45054 56866 45106
rect 57038 45054 57090 45106
rect 6750 44942 6802 44994
rect 8878 44942 8930 44994
rect 15710 44942 15762 44994
rect 20974 44942 21026 44994
rect 23102 44942 23154 44994
rect 24670 44942 24722 44994
rect 29150 44942 29202 44994
rect 31950 44942 32002 44994
rect 33294 44942 33346 44994
rect 35422 44942 35474 44994
rect 52894 44942 52946 44994
rect 57710 44942 57762 44994
rect 4958 44830 5010 44882
rect 24446 44830 24498 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 3502 44494 3554 44546
rect 9326 44494 9378 44546
rect 9662 44494 9714 44546
rect 16270 44494 16322 44546
rect 31726 44494 31778 44546
rect 45390 44494 45442 44546
rect 51214 44494 51266 44546
rect 54574 44494 54626 44546
rect 55246 44494 55298 44546
rect 56142 44494 56194 44546
rect 4062 44382 4114 44434
rect 5630 44382 5682 44434
rect 5966 44382 6018 44434
rect 7310 44382 7362 44434
rect 8094 44382 8146 44434
rect 8990 44382 9042 44434
rect 9550 44382 9602 44434
rect 16830 44382 16882 44434
rect 19630 44382 19682 44434
rect 24110 44382 24162 44434
rect 31390 44382 31442 44434
rect 32286 44382 32338 44434
rect 43598 44382 43650 44434
rect 45502 44382 45554 44434
rect 51774 44382 51826 44434
rect 54238 44382 54290 44434
rect 57598 44382 57650 44434
rect 58270 44382 58322 44434
rect 2494 44270 2546 44322
rect 4510 44270 4562 44322
rect 4958 44270 5010 44322
rect 6190 44270 6242 44322
rect 7534 44270 7586 44322
rect 7758 44270 7810 44322
rect 8766 44270 8818 44322
rect 15486 44270 15538 44322
rect 16158 44270 16210 44322
rect 17278 44270 17330 44322
rect 17838 44270 17890 44322
rect 18510 44270 18562 44322
rect 21758 44270 21810 44322
rect 22094 44270 22146 44322
rect 23326 44270 23378 44322
rect 24782 44270 24834 44322
rect 25790 44270 25842 44322
rect 31166 44270 31218 44322
rect 32398 44270 32450 44322
rect 33070 44270 33122 44322
rect 33742 44270 33794 44322
rect 34302 44270 34354 44322
rect 34750 44270 34802 44322
rect 35310 44270 35362 44322
rect 40798 44270 40850 44322
rect 44270 44270 44322 44322
rect 44718 44270 44770 44322
rect 45614 44270 45666 44322
rect 46510 44270 46562 44322
rect 46958 44270 47010 44322
rect 51886 44270 51938 44322
rect 55470 44270 55522 44322
rect 56590 44270 56642 44322
rect 2830 44158 2882 44210
rect 3502 44158 3554 44210
rect 3614 44158 3666 44210
rect 3950 44158 4002 44210
rect 7198 44158 7250 44210
rect 13470 44158 13522 44210
rect 16942 44158 16994 44210
rect 22318 44158 22370 44210
rect 22654 44158 22706 44210
rect 24446 44158 24498 44210
rect 25566 44158 25618 44210
rect 34078 44158 34130 44210
rect 41470 44158 41522 44210
rect 43934 44158 43986 44210
rect 44046 44158 44098 44210
rect 46846 44158 46898 44210
rect 56702 44158 56754 44210
rect 56814 44158 56866 44210
rect 2718 44046 2770 44098
rect 13806 44046 13858 44098
rect 22766 44046 22818 44098
rect 22878 44046 22930 44098
rect 23662 44046 23714 44098
rect 33966 44046 34018 44098
rect 34638 44046 34690 44098
rect 34862 44046 34914 44098
rect 35646 44046 35698 44098
rect 37886 44046 37938 44098
rect 46622 44046 46674 44098
rect 54350 44046 54402 44098
rect 54910 44046 54962 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4958 43710 5010 43762
rect 23214 43710 23266 43762
rect 32398 43710 32450 43762
rect 37662 43710 37714 43762
rect 2494 43598 2546 43650
rect 5070 43598 5122 43650
rect 5518 43598 5570 43650
rect 15374 43598 15426 43650
rect 15598 43598 15650 43650
rect 16382 43598 16434 43650
rect 17726 43598 17778 43650
rect 18286 43598 18338 43650
rect 22206 43598 22258 43650
rect 22542 43598 22594 43650
rect 22766 43598 22818 43650
rect 29822 43598 29874 43650
rect 36654 43598 36706 43650
rect 38558 43598 38610 43650
rect 46062 43598 46114 43650
rect 57374 43598 57426 43650
rect 57822 43598 57874 43650
rect 1822 43486 1874 43538
rect 15710 43486 15762 43538
rect 17614 43486 17666 43538
rect 19070 43486 19122 43538
rect 29710 43486 29762 43538
rect 29934 43486 29986 43538
rect 30270 43486 30322 43538
rect 31838 43486 31890 43538
rect 32062 43486 32114 43538
rect 37102 43486 37154 43538
rect 37774 43486 37826 43538
rect 39678 43486 39730 43538
rect 41022 43486 41074 43538
rect 41470 43486 41522 43538
rect 45390 43486 45442 43538
rect 52782 43486 52834 43538
rect 53230 43486 53282 43538
rect 4622 43374 4674 43426
rect 16494 43374 16546 43426
rect 17390 43374 17442 43426
rect 19742 43374 19794 43426
rect 21870 43374 21922 43426
rect 22318 43374 22370 43426
rect 38222 43374 38274 43426
rect 40350 43374 40402 43426
rect 42478 43374 42530 43426
rect 44942 43374 44994 43426
rect 48190 43374 48242 43426
rect 54798 43374 54850 43426
rect 57150 43374 57202 43426
rect 16158 43262 16210 43314
rect 57598 43262 57650 43314
rect 57822 43262 57874 43314
rect 58158 43262 58210 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 10110 42926 10162 42978
rect 20190 42926 20242 42978
rect 33182 42926 33234 42978
rect 34078 42926 34130 42978
rect 37102 42926 37154 42978
rect 45614 42926 45666 42978
rect 50094 42926 50146 42978
rect 53566 42926 53618 42978
rect 53678 42926 53730 42978
rect 53902 42926 53954 42978
rect 2942 42814 2994 42866
rect 3726 42814 3778 42866
rect 13022 42814 13074 42866
rect 16830 42814 16882 42866
rect 22094 42814 22146 42866
rect 25342 42814 25394 42866
rect 31054 42814 31106 42866
rect 33182 42814 33234 42866
rect 34078 42814 34130 42866
rect 40126 42814 40178 42866
rect 41582 42814 41634 42866
rect 44158 42814 44210 42866
rect 46734 42814 46786 42866
rect 51662 42814 51714 42866
rect 53118 42814 53170 42866
rect 57038 42814 57090 42866
rect 3614 42702 3666 42754
rect 8430 42702 8482 42754
rect 8766 42702 8818 42754
rect 9662 42702 9714 42754
rect 10110 42702 10162 42754
rect 10558 42702 10610 42754
rect 14030 42702 14082 42754
rect 14478 42702 14530 42754
rect 15374 42702 15426 42754
rect 15710 42702 15762 42754
rect 15934 42702 15986 42754
rect 16494 42702 16546 42754
rect 18174 42702 18226 42754
rect 19406 42702 19458 42754
rect 25230 42702 25282 42754
rect 26014 42702 26066 42754
rect 26238 42702 26290 42754
rect 27134 42702 27186 42754
rect 27470 42702 27522 42754
rect 27694 42702 27746 42754
rect 28366 42702 28418 42754
rect 29150 42702 29202 42754
rect 30046 42702 30098 42754
rect 30942 42702 30994 42754
rect 37550 42702 37602 42754
rect 38110 42702 38162 42754
rect 39230 42702 39282 42754
rect 39454 42702 39506 42754
rect 46622 42702 46674 42754
rect 51550 42702 51602 42754
rect 51774 42702 51826 42754
rect 55918 42702 55970 42754
rect 56478 42702 56530 42754
rect 9102 42590 9154 42642
rect 13918 42590 13970 42642
rect 16830 42590 16882 42642
rect 20302 42590 20354 42642
rect 20750 42590 20802 42642
rect 25118 42590 25170 42642
rect 30494 42590 30546 42642
rect 31278 42590 31330 42642
rect 37214 42590 37266 42642
rect 38558 42590 38610 42642
rect 41694 42590 41746 42642
rect 42030 42590 42082 42642
rect 42254 42590 42306 42642
rect 43934 42590 43986 42642
rect 45614 42590 45666 42642
rect 45726 42590 45778 42642
rect 50206 42590 50258 42642
rect 54014 42590 54066 42642
rect 55470 42590 55522 42642
rect 56926 42590 56978 42642
rect 8990 42478 9042 42530
rect 14366 42478 14418 42530
rect 20526 42478 20578 42530
rect 21422 42478 21474 42530
rect 28478 42478 28530 42530
rect 28702 42478 28754 42530
rect 29262 42478 29314 42530
rect 29486 42478 29538 42530
rect 33630 42478 33682 42530
rect 36430 42478 36482 42530
rect 37102 42478 37154 42530
rect 37662 42478 37714 42530
rect 41022 42478 41074 42530
rect 41470 42478 41522 42530
rect 45166 42478 45218 42530
rect 46398 42478 46450 42530
rect 46846 42478 46898 42530
rect 49646 42478 49698 42530
rect 50094 42478 50146 42530
rect 51998 42478 52050 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 14478 42142 14530 42194
rect 20974 42142 21026 42194
rect 28030 42142 28082 42194
rect 28478 42142 28530 42194
rect 58158 42142 58210 42194
rect 8766 42030 8818 42082
rect 9662 42030 9714 42082
rect 11566 42030 11618 42082
rect 15598 42030 15650 42082
rect 18398 42030 18450 42082
rect 20526 42030 20578 42082
rect 23886 42030 23938 42082
rect 24110 42030 24162 42082
rect 24446 42030 24498 42082
rect 24558 42030 24610 42082
rect 27246 42030 27298 42082
rect 34078 42030 34130 42082
rect 35534 42030 35586 42082
rect 43486 42030 43538 42082
rect 53790 42030 53842 42082
rect 57038 42030 57090 42082
rect 57598 42030 57650 42082
rect 5406 41918 5458 41970
rect 6078 41918 6130 41970
rect 8878 41918 8930 41970
rect 9550 41918 9602 41970
rect 9886 41918 9938 41970
rect 10222 41918 10274 41970
rect 12798 41918 12850 41970
rect 14142 41918 14194 41970
rect 14478 41918 14530 41970
rect 14814 41918 14866 41970
rect 15262 41918 15314 41970
rect 15486 41918 15538 41970
rect 15934 41918 15986 41970
rect 16718 41918 16770 41970
rect 18286 41918 18338 41970
rect 19854 41918 19906 41970
rect 20638 41918 20690 41970
rect 21422 41918 21474 41970
rect 23550 41918 23602 41970
rect 24782 41918 24834 41970
rect 25118 41918 25170 41970
rect 25902 41918 25954 41970
rect 26910 41918 26962 41970
rect 27918 41918 27970 41970
rect 28142 41918 28194 41970
rect 28590 41918 28642 41970
rect 28702 41918 28754 41970
rect 29038 41918 29090 41970
rect 29486 41918 29538 41970
rect 29710 41918 29762 41970
rect 30382 41918 30434 41970
rect 33742 41918 33794 41970
rect 35870 41918 35922 41970
rect 36878 41918 36930 41970
rect 38782 41918 38834 41970
rect 40350 41918 40402 41970
rect 41134 41918 41186 41970
rect 41358 41918 41410 41970
rect 41806 41918 41858 41970
rect 43822 41918 43874 41970
rect 49198 41918 49250 41970
rect 52446 41918 52498 41970
rect 53118 41918 53170 41970
rect 56702 41918 56754 41970
rect 57374 41918 57426 41970
rect 3278 41806 3330 41858
rect 8206 41806 8258 41858
rect 11006 41806 11058 41858
rect 21198 41806 21250 41858
rect 25790 41806 25842 41858
rect 32510 41806 32562 41858
rect 34414 41806 34466 41858
rect 37214 41806 37266 41858
rect 38110 41806 38162 41858
rect 38894 41806 38946 41858
rect 39454 41806 39506 41858
rect 41246 41806 41298 41858
rect 44494 41806 44546 41858
rect 49870 41806 49922 41858
rect 51998 41806 52050 41858
rect 55918 41806 55970 41858
rect 57486 41806 57538 41858
rect 8990 41694 9042 41746
rect 13806 41694 13858 41746
rect 19966 41694 20018 41746
rect 24222 41694 24274 41746
rect 25678 41694 25730 41746
rect 27694 41694 27746 41746
rect 33406 41694 33458 41746
rect 33742 41694 33794 41746
rect 34638 41694 34690 41746
rect 43822 41694 43874 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14030 41358 14082 41410
rect 27134 41358 27186 41410
rect 27358 41358 27410 41410
rect 32174 41358 32226 41410
rect 33518 41358 33570 41410
rect 44158 41358 44210 41410
rect 50318 41358 50370 41410
rect 52894 41358 52946 41410
rect 2718 41246 2770 41298
rect 4510 41246 4562 41298
rect 9998 41246 10050 41298
rect 14702 41246 14754 41298
rect 20078 41246 20130 41298
rect 21310 41246 21362 41298
rect 23214 41246 23266 41298
rect 23774 41246 23826 41298
rect 25566 41246 25618 41298
rect 32510 41246 32562 41298
rect 34862 41246 34914 41298
rect 36990 41246 37042 41298
rect 38558 41246 38610 41298
rect 40126 41246 40178 41298
rect 43486 41246 43538 41298
rect 45166 41246 45218 41298
rect 45502 41246 45554 41298
rect 48638 41246 48690 41298
rect 50542 41246 50594 41298
rect 52670 41246 52722 41298
rect 4062 41134 4114 41186
rect 5182 41134 5234 41186
rect 5518 41134 5570 41186
rect 8654 41134 8706 41186
rect 12126 41134 12178 41186
rect 15822 41134 15874 41186
rect 17390 41134 17442 41186
rect 19070 41134 19122 41186
rect 19854 41134 19906 41186
rect 23326 41134 23378 41186
rect 25230 41134 25282 41186
rect 25454 41134 25506 41186
rect 25902 41134 25954 41186
rect 26574 41134 26626 41186
rect 29038 41134 29090 41186
rect 32062 41134 32114 41186
rect 33182 41134 33234 41186
rect 33518 41134 33570 41186
rect 33966 41134 34018 41186
rect 34638 41134 34690 41186
rect 35534 41134 35586 41186
rect 35758 41134 35810 41186
rect 36094 41134 36146 41186
rect 37102 41134 37154 41186
rect 37662 41134 37714 41186
rect 43038 41134 43090 41186
rect 50654 41134 50706 41186
rect 51662 41134 51714 41186
rect 51886 41134 51938 41186
rect 51998 41134 52050 41186
rect 53118 41134 53170 41186
rect 55694 41134 55746 41186
rect 57598 41134 57650 41186
rect 2830 41022 2882 41074
rect 3054 41022 3106 41074
rect 3726 41022 3778 41074
rect 5854 41022 5906 41074
rect 9662 41022 9714 41074
rect 12350 41022 12402 41074
rect 12462 41022 12514 41074
rect 13470 41022 13522 41074
rect 13918 41022 13970 41074
rect 16382 41022 16434 41074
rect 17502 41022 17554 41074
rect 18846 41022 18898 41074
rect 20302 41022 20354 41074
rect 20526 41022 20578 41074
rect 26462 41022 26514 41074
rect 26686 41022 26738 41074
rect 27918 41022 27970 41074
rect 29374 41022 29426 41074
rect 34750 41022 34802 41074
rect 42254 41022 42306 41074
rect 44270 41022 44322 41074
rect 51550 41022 51602 41074
rect 55358 41022 55410 41074
rect 57262 41022 57314 41074
rect 5742 40910 5794 40962
rect 8318 40910 8370 40962
rect 13694 40910 13746 40962
rect 15150 40910 15202 40962
rect 21870 40910 21922 40962
rect 22318 40910 22370 40962
rect 27470 40910 27522 40962
rect 27694 40910 27746 40962
rect 29262 40910 29314 40962
rect 34974 40910 35026 40962
rect 35086 40910 35138 40962
rect 44158 40910 44210 40962
rect 45390 40910 45442 40962
rect 49086 40910 49138 40962
rect 53566 40910 53618 40962
rect 56030 40910 56082 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 2718 40574 2770 40626
rect 5070 40574 5122 40626
rect 8094 40574 8146 40626
rect 14030 40574 14082 40626
rect 19406 40574 19458 40626
rect 20414 40574 20466 40626
rect 20974 40574 21026 40626
rect 21422 40574 21474 40626
rect 41134 40574 41186 40626
rect 55694 40574 55746 40626
rect 55918 40574 55970 40626
rect 58158 40574 58210 40626
rect 4286 40462 4338 40514
rect 5294 40462 5346 40514
rect 16718 40462 16770 40514
rect 17950 40462 18002 40514
rect 22878 40462 22930 40514
rect 34862 40462 34914 40514
rect 35646 40462 35698 40514
rect 38782 40462 38834 40514
rect 40238 40462 40290 40514
rect 40350 40462 40402 40514
rect 44046 40462 44098 40514
rect 45838 40462 45890 40514
rect 56926 40462 56978 40514
rect 3054 40350 3106 40402
rect 3950 40350 4002 40402
rect 7758 40350 7810 40402
rect 15038 40350 15090 40402
rect 15822 40350 15874 40402
rect 17502 40350 17554 40402
rect 20302 40350 20354 40402
rect 23438 40350 23490 40402
rect 23886 40350 23938 40402
rect 27134 40350 27186 40402
rect 27806 40350 27858 40402
rect 28926 40350 28978 40402
rect 29262 40350 29314 40402
rect 31390 40350 31442 40402
rect 34190 40350 34242 40402
rect 35758 40350 35810 40402
rect 37886 40350 37938 40402
rect 40798 40350 40850 40402
rect 41246 40350 41298 40402
rect 41358 40350 41410 40402
rect 43822 40350 43874 40402
rect 44606 40350 44658 40402
rect 45054 40350 45106 40402
rect 51662 40350 51714 40402
rect 56030 40350 56082 40402
rect 57038 40350 57090 40402
rect 57486 40350 57538 40402
rect 4958 40238 5010 40290
rect 19182 40238 19234 40290
rect 22990 40238 23042 40290
rect 27582 40238 27634 40290
rect 28030 40238 28082 40290
rect 29486 40238 29538 40290
rect 31166 40238 31218 40290
rect 35870 40238 35922 40290
rect 38110 40238 38162 40290
rect 43598 40238 43650 40290
rect 47966 40238 48018 40290
rect 50990 40238 51042 40290
rect 51774 40238 51826 40290
rect 57262 40238 57314 40290
rect 15150 40126 15202 40178
rect 16494 40126 16546 40178
rect 20414 40126 20466 40178
rect 22654 40126 22706 40178
rect 40238 40126 40290 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 14926 39790 14978 39842
rect 26014 39790 26066 39842
rect 45838 39790 45890 39842
rect 51326 39790 51378 39842
rect 57486 39790 57538 39842
rect 57822 39790 57874 39842
rect 2494 39678 2546 39730
rect 4622 39678 4674 39730
rect 5070 39678 5122 39730
rect 6862 39678 6914 39730
rect 17726 39678 17778 39730
rect 18846 39678 18898 39730
rect 20750 39678 20802 39730
rect 22206 39678 22258 39730
rect 26126 39678 26178 39730
rect 27918 39678 27970 39730
rect 32174 39678 32226 39730
rect 32510 39678 32562 39730
rect 34638 39678 34690 39730
rect 35198 39678 35250 39730
rect 43374 39678 43426 39730
rect 45278 39678 45330 39730
rect 47518 39678 47570 39730
rect 50990 39678 51042 39730
rect 56478 39678 56530 39730
rect 1822 39566 1874 39618
rect 11454 39566 11506 39618
rect 12350 39566 12402 39618
rect 14142 39566 14194 39618
rect 14926 39566 14978 39618
rect 15486 39566 15538 39618
rect 17502 39566 17554 39618
rect 18958 39566 19010 39618
rect 19294 39566 19346 39618
rect 22654 39566 22706 39618
rect 23774 39566 23826 39618
rect 25566 39566 25618 39618
rect 26238 39566 26290 39618
rect 26574 39566 26626 39618
rect 31278 39566 31330 39618
rect 31502 39566 31554 39618
rect 34862 39566 34914 39618
rect 41694 39566 41746 39618
rect 43822 39566 43874 39618
rect 45390 39566 45442 39618
rect 47406 39566 47458 39618
rect 53678 39566 53730 39618
rect 57038 39566 57090 39618
rect 12910 39454 12962 39506
rect 16494 39454 16546 39506
rect 25006 39454 25058 39506
rect 37550 39454 37602 39506
rect 44270 39454 44322 39506
rect 45054 39454 45106 39506
rect 45726 39454 45778 39506
rect 49310 39454 49362 39506
rect 54350 39454 54402 39506
rect 57598 39454 57650 39506
rect 11678 39342 11730 39394
rect 12574 39342 12626 39394
rect 17390 39342 17442 39394
rect 20190 39342 20242 39394
rect 24110 39342 24162 39394
rect 27470 39342 27522 39394
rect 33070 39342 33122 39394
rect 37886 39342 37938 39394
rect 42254 39342 42306 39394
rect 45838 39342 45890 39394
rect 48974 39342 49026 39394
rect 49758 39342 49810 39394
rect 50654 39342 50706 39394
rect 51102 39342 51154 39394
rect 56814 39342 56866 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 6190 39006 6242 39058
rect 8206 39006 8258 39058
rect 13022 39006 13074 39058
rect 27694 39006 27746 39058
rect 27918 39006 27970 39058
rect 44718 39006 44770 39058
rect 53566 39006 53618 39058
rect 54126 39006 54178 39058
rect 7870 38894 7922 38946
rect 7982 38894 8034 38946
rect 12014 38894 12066 38946
rect 12238 38894 12290 38946
rect 19854 38894 19906 38946
rect 20414 38894 20466 38946
rect 20974 38894 21026 38946
rect 30382 38894 30434 38946
rect 36542 38894 36594 38946
rect 38110 38894 38162 38946
rect 39006 38894 39058 38946
rect 50990 38894 51042 38946
rect 57822 38894 57874 38946
rect 6414 38782 6466 38834
rect 6638 38782 6690 38834
rect 7086 38782 7138 38834
rect 11454 38782 11506 38834
rect 12462 38782 12514 38834
rect 12574 38782 12626 38834
rect 15598 38782 15650 38834
rect 16382 38782 16434 38834
rect 18062 38782 18114 38834
rect 18510 38782 18562 38834
rect 18846 38782 18898 38834
rect 20750 38782 20802 38834
rect 23438 38782 23490 38834
rect 23662 38782 23714 38834
rect 23886 38782 23938 38834
rect 24110 38782 24162 38834
rect 25678 38782 25730 38834
rect 26350 38782 26402 38834
rect 27022 38782 27074 38834
rect 27246 38782 27298 38834
rect 28030 38782 28082 38834
rect 30046 38782 30098 38834
rect 30606 38782 30658 38834
rect 32510 38782 32562 38834
rect 34078 38782 34130 38834
rect 34750 38782 34802 38834
rect 36878 38782 36930 38834
rect 37438 38782 37490 38834
rect 39678 38782 39730 38834
rect 40014 38782 40066 38834
rect 48862 38782 48914 38834
rect 50206 38782 50258 38834
rect 57598 38782 57650 38834
rect 58046 38782 58098 38834
rect 6526 38670 6578 38722
rect 7534 38670 7586 38722
rect 11678 38670 11730 38722
rect 15822 38670 15874 38722
rect 18622 38670 18674 38722
rect 25566 38670 25618 38722
rect 29934 38670 29986 38722
rect 32174 38670 32226 38722
rect 34302 38670 34354 38722
rect 34862 38670 34914 38722
rect 39230 38670 39282 38722
rect 45950 38670 46002 38722
rect 46174 38670 46226 38722
rect 49422 38670 49474 38722
rect 53118 38670 53170 38722
rect 53902 38670 53954 38722
rect 54238 38670 54290 38722
rect 56702 38670 56754 38722
rect 11118 38558 11170 38610
rect 15374 38558 15426 38610
rect 24222 38558 24274 38610
rect 26798 38558 26850 38610
rect 30270 38558 30322 38610
rect 30830 38558 30882 38610
rect 31950 38558 32002 38610
rect 46510 38558 46562 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 3950 38222 4002 38274
rect 9886 38222 9938 38274
rect 11790 38222 11842 38274
rect 12238 38222 12290 38274
rect 12574 38222 12626 38274
rect 13694 38222 13746 38274
rect 15374 38222 15426 38274
rect 16718 38222 16770 38274
rect 19070 38222 19122 38274
rect 24558 38222 24610 38274
rect 26014 38222 26066 38274
rect 27358 38222 27410 38274
rect 29262 38222 29314 38274
rect 30494 38222 30546 38274
rect 35534 38222 35586 38274
rect 4510 38110 4562 38162
rect 6750 38110 6802 38162
rect 12798 38110 12850 38162
rect 16606 38110 16658 38162
rect 18622 38110 18674 38162
rect 27022 38110 27074 38162
rect 28142 38110 28194 38162
rect 38782 38110 38834 38162
rect 46398 38110 46450 38162
rect 58158 38110 58210 38162
rect 4062 37998 4114 38050
rect 5854 37998 5906 38050
rect 6190 37998 6242 38050
rect 6414 37998 6466 38050
rect 7198 37998 7250 38050
rect 8878 37998 8930 38050
rect 9550 37998 9602 38050
rect 11454 37998 11506 38050
rect 14030 37998 14082 38050
rect 14814 37998 14866 38050
rect 15374 37998 15426 38050
rect 18510 37998 18562 38050
rect 20750 37998 20802 38050
rect 24222 37998 24274 38050
rect 26126 37998 26178 38050
rect 27134 37998 27186 38050
rect 27470 37998 27522 38050
rect 28590 37998 28642 38050
rect 31278 37998 31330 38050
rect 32958 37998 33010 38050
rect 34414 37998 34466 38050
rect 38110 37998 38162 38050
rect 40238 37998 40290 38050
rect 41582 37998 41634 38050
rect 42142 37998 42194 38050
rect 45390 37998 45442 38050
rect 45838 37998 45890 38050
rect 49310 37998 49362 38050
rect 54910 37998 54962 38050
rect 55358 37998 55410 38050
rect 8766 37886 8818 37938
rect 10670 37886 10722 37938
rect 11230 37886 11282 37938
rect 14702 37886 14754 37938
rect 17054 37886 17106 37938
rect 21310 37886 21362 37938
rect 23998 37886 24050 37938
rect 28142 37886 28194 37938
rect 29262 37886 29314 37938
rect 29374 37886 29426 37938
rect 30606 37886 30658 37938
rect 31838 37886 31890 37938
rect 35086 37886 35138 37938
rect 35646 37886 35698 37938
rect 37214 37886 37266 37938
rect 37998 37886 38050 37938
rect 39006 37886 39058 37938
rect 46062 37886 46114 37938
rect 48526 37886 48578 37938
rect 56030 37886 56082 37938
rect 3950 37774 4002 37826
rect 5966 37774 6018 37826
rect 21646 37774 21698 37826
rect 22206 37774 22258 37826
rect 26014 37774 26066 37826
rect 28366 37774 28418 37826
rect 30158 37774 30210 37826
rect 30494 37774 30546 37826
rect 30830 37774 30882 37826
rect 35534 37774 35586 37826
rect 37438 37774 37490 37826
rect 40798 37774 40850 37826
rect 45278 37774 45330 37826
rect 45950 37774 46002 37826
rect 49758 37774 49810 37826
rect 53566 37774 53618 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 3614 37438 3666 37490
rect 12686 37438 12738 37490
rect 15150 37438 15202 37490
rect 15486 37438 15538 37490
rect 24558 37438 24610 37490
rect 25342 37438 25394 37490
rect 30718 37438 30770 37490
rect 37102 37438 37154 37490
rect 39006 37438 39058 37490
rect 39902 37438 39954 37490
rect 44270 37438 44322 37490
rect 46622 37438 46674 37490
rect 46734 37438 46786 37490
rect 56702 37438 56754 37490
rect 2718 37326 2770 37378
rect 3054 37326 3106 37378
rect 5294 37326 5346 37378
rect 8542 37326 8594 37378
rect 8654 37326 8706 37378
rect 8766 37326 8818 37378
rect 9886 37326 9938 37378
rect 11342 37326 11394 37378
rect 12014 37326 12066 37378
rect 12462 37326 12514 37378
rect 14814 37326 14866 37378
rect 14926 37326 14978 37378
rect 18286 37326 18338 37378
rect 18958 37326 19010 37378
rect 23662 37326 23714 37378
rect 26014 37326 26066 37378
rect 26126 37326 26178 37378
rect 26798 37326 26850 37378
rect 35758 37326 35810 37378
rect 37214 37326 37266 37378
rect 37774 37326 37826 37378
rect 39566 37326 39618 37378
rect 39678 37326 39730 37378
rect 46510 37326 46562 37378
rect 3166 37214 3218 37266
rect 3726 37214 3778 37266
rect 3838 37214 3890 37266
rect 4286 37214 4338 37266
rect 4622 37214 4674 37266
rect 7870 37214 7922 37266
rect 8990 37214 9042 37266
rect 9438 37214 9490 37266
rect 10222 37214 10274 37266
rect 11902 37214 11954 37266
rect 15486 37214 15538 37266
rect 15598 37214 15650 37266
rect 16382 37214 16434 37266
rect 17390 37214 17442 37266
rect 17950 37214 18002 37266
rect 19630 37214 19682 37266
rect 20414 37214 20466 37266
rect 20862 37214 20914 37266
rect 24670 37214 24722 37266
rect 26574 37214 26626 37266
rect 27134 37214 27186 37266
rect 27582 37214 27634 37266
rect 29150 37214 29202 37266
rect 31278 37214 31330 37266
rect 33518 37214 33570 37266
rect 33854 37214 33906 37266
rect 35982 37214 36034 37266
rect 37998 37214 38050 37266
rect 39230 37214 39282 37266
rect 43822 37214 43874 37266
rect 2830 37102 2882 37154
rect 7422 37102 7474 37154
rect 8766 37102 8818 37154
rect 15822 37102 15874 37154
rect 16718 37102 16770 37154
rect 18398 37102 18450 37154
rect 19742 37102 19794 37154
rect 20750 37102 20802 37154
rect 22878 37102 22930 37154
rect 25230 37102 25282 37154
rect 34078 37102 34130 37154
rect 40910 37102 40962 37154
rect 43038 37102 43090 37154
rect 11118 36990 11170 37042
rect 27246 36990 27298 37042
rect 31054 36990 31106 37042
rect 38894 36990 38946 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 8878 36654 8930 36706
rect 16158 36654 16210 36706
rect 16942 36654 16994 36706
rect 23102 36654 23154 36706
rect 24558 36654 24610 36706
rect 27358 36654 27410 36706
rect 35646 36654 35698 36706
rect 36878 36654 36930 36706
rect 40910 36654 40962 36706
rect 41246 36654 41298 36706
rect 2494 36542 2546 36594
rect 4622 36542 4674 36594
rect 5182 36542 5234 36594
rect 9326 36542 9378 36594
rect 12014 36542 12066 36594
rect 15934 36542 15986 36594
rect 16830 36542 16882 36594
rect 18510 36542 18562 36594
rect 22542 36542 22594 36594
rect 24110 36542 24162 36594
rect 28254 36542 28306 36594
rect 30718 36542 30770 36594
rect 35534 36542 35586 36594
rect 37886 36542 37938 36594
rect 52110 36542 52162 36594
rect 52894 36542 52946 36594
rect 56142 36542 56194 36594
rect 1822 36430 1874 36482
rect 11118 36430 11170 36482
rect 11454 36430 11506 36482
rect 12350 36430 12402 36482
rect 15710 36430 15762 36482
rect 17166 36430 17218 36482
rect 17502 36430 17554 36482
rect 18846 36430 18898 36482
rect 20190 36430 20242 36482
rect 22766 36430 22818 36482
rect 23998 36430 24050 36482
rect 24334 36430 24386 36482
rect 24670 36430 24722 36482
rect 26910 36430 26962 36482
rect 27246 36430 27298 36482
rect 31502 36430 31554 36482
rect 33294 36430 33346 36482
rect 35422 36430 35474 36482
rect 36094 36430 36146 36482
rect 37102 36430 37154 36482
rect 37550 36430 37602 36482
rect 37662 36430 37714 36482
rect 38558 36430 38610 36482
rect 49310 36430 49362 36482
rect 53342 36430 53394 36482
rect 57038 36430 57090 36482
rect 57374 36430 57426 36482
rect 8766 36318 8818 36370
rect 11566 36318 11618 36370
rect 19070 36318 19122 36370
rect 23662 36318 23714 36370
rect 32062 36318 32114 36370
rect 38222 36318 38274 36370
rect 44046 36318 44098 36370
rect 49982 36318 50034 36370
rect 54014 36318 54066 36370
rect 56702 36318 56754 36370
rect 8878 36206 8930 36258
rect 9886 36206 9938 36258
rect 10782 36206 10834 36258
rect 11006 36206 11058 36258
rect 12686 36206 12738 36258
rect 21310 36206 21362 36258
rect 21646 36206 21698 36258
rect 27806 36206 27858 36258
rect 31166 36206 31218 36258
rect 32958 36206 33010 36258
rect 41134 36206 41186 36258
rect 41694 36206 41746 36258
rect 43822 36206 43874 36258
rect 43934 36206 43986 36258
rect 57150 36206 57202 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 11678 35870 11730 35922
rect 15598 35870 15650 35922
rect 18958 35870 19010 35922
rect 23326 35870 23378 35922
rect 24222 35870 24274 35922
rect 25230 35870 25282 35922
rect 27246 35870 27298 35922
rect 28366 35870 28418 35922
rect 31502 35870 31554 35922
rect 37662 35870 37714 35922
rect 38222 35870 38274 35922
rect 39006 35870 39058 35922
rect 39230 35870 39282 35922
rect 50430 35870 50482 35922
rect 51214 35870 51266 35922
rect 55134 35870 55186 35922
rect 56702 35870 56754 35922
rect 57262 35870 57314 35922
rect 57486 35870 57538 35922
rect 57822 35870 57874 35922
rect 58046 35870 58098 35922
rect 17950 35758 18002 35810
rect 27358 35758 27410 35810
rect 30942 35758 30994 35810
rect 32398 35758 32450 35810
rect 34974 35758 35026 35810
rect 37214 35758 37266 35810
rect 37438 35758 37490 35810
rect 38334 35758 38386 35810
rect 44830 35758 44882 35810
rect 51998 35758 52050 35810
rect 1822 35646 1874 35698
rect 11342 35646 11394 35698
rect 11678 35646 11730 35698
rect 12014 35646 12066 35698
rect 16158 35646 16210 35698
rect 18846 35646 18898 35698
rect 20302 35646 20354 35698
rect 22766 35646 22818 35698
rect 23998 35646 24050 35698
rect 30494 35646 30546 35698
rect 31390 35646 31442 35698
rect 32510 35646 32562 35698
rect 35870 35646 35922 35698
rect 37886 35646 37938 35698
rect 38558 35646 38610 35698
rect 38894 35646 38946 35698
rect 39342 35646 39394 35698
rect 42478 35646 42530 35698
rect 45502 35646 45554 35698
rect 50654 35646 50706 35698
rect 52894 35646 52946 35698
rect 54910 35646 54962 35698
rect 55358 35646 55410 35698
rect 55582 35646 55634 35698
rect 56478 35646 56530 35698
rect 56814 35646 56866 35698
rect 57150 35646 57202 35698
rect 57710 35646 57762 35698
rect 2270 35534 2322 35586
rect 19182 35534 19234 35586
rect 20750 35534 20802 35586
rect 21310 35534 21362 35586
rect 25678 35534 25730 35586
rect 33630 35534 33682 35586
rect 34190 35534 34242 35586
rect 42702 35534 42754 35586
rect 51998 35534 52050 35586
rect 15934 35422 15986 35474
rect 32398 35422 32450 35474
rect 50318 35422 50370 35474
rect 50878 35422 50930 35474
rect 51214 35422 51266 35474
rect 51774 35422 51826 35474
rect 53118 35422 53170 35474
rect 53454 35422 53506 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 10446 35086 10498 35138
rect 12126 35086 12178 35138
rect 14254 35086 14306 35138
rect 17278 35086 17330 35138
rect 44942 35086 44994 35138
rect 1822 34974 1874 35026
rect 8654 34974 8706 35026
rect 15822 34974 15874 35026
rect 19070 34974 19122 35026
rect 19518 34974 19570 35026
rect 20862 34974 20914 35026
rect 24222 34974 24274 35026
rect 27918 34974 27970 35026
rect 29710 34974 29762 35026
rect 33742 34974 33794 35026
rect 35758 34974 35810 35026
rect 37662 34974 37714 35026
rect 38222 34974 38274 35026
rect 44046 34974 44098 35026
rect 45502 34974 45554 35026
rect 46062 34974 46114 35026
rect 49982 34974 50034 35026
rect 7870 34862 7922 34914
rect 8206 34862 8258 34914
rect 8430 34862 8482 34914
rect 9550 34862 9602 34914
rect 9998 34862 10050 34914
rect 10558 34862 10610 34914
rect 10894 34862 10946 34914
rect 11454 34862 11506 34914
rect 12574 34862 12626 34914
rect 13470 34862 13522 34914
rect 16270 34862 16322 34914
rect 16606 34862 16658 34914
rect 16830 34862 16882 34914
rect 17838 34862 17890 34914
rect 19966 34862 20018 34914
rect 21310 34862 21362 34914
rect 29822 34862 29874 34914
rect 30158 34862 30210 34914
rect 36206 34862 36258 34914
rect 37214 34862 37266 34914
rect 38334 34862 38386 34914
rect 48862 34862 48914 34914
rect 53230 34862 53282 34914
rect 8766 34750 8818 34802
rect 12910 34750 12962 34802
rect 13694 34750 13746 34802
rect 13806 34750 13858 34802
rect 17950 34750 18002 34802
rect 18510 34750 18562 34802
rect 22094 34750 22146 34802
rect 37998 34750 38050 34802
rect 43598 34750 43650 34802
rect 43822 34750 43874 34802
rect 44158 34750 44210 34802
rect 44942 34750 44994 34802
rect 48190 34750 48242 34802
rect 49422 34750 49474 34802
rect 7982 34638 8034 34690
rect 11790 34638 11842 34690
rect 12014 34638 12066 34690
rect 12686 34638 12738 34690
rect 28366 34638 28418 34690
rect 29374 34638 29426 34690
rect 29598 34638 29650 34690
rect 38782 34638 38834 34690
rect 45054 34694 45106 34746
rect 49534 34750 49586 34802
rect 56926 34750 56978 34802
rect 57038 34750 57090 34802
rect 53454 34638 53506 34690
rect 56702 34638 56754 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 9662 34302 9714 34354
rect 11118 34302 11170 34354
rect 18622 34302 18674 34354
rect 29150 34302 29202 34354
rect 29822 34302 29874 34354
rect 30046 34302 30098 34354
rect 34078 34302 34130 34354
rect 41470 34302 41522 34354
rect 42366 34302 42418 34354
rect 44270 34302 44322 34354
rect 44494 34302 44546 34354
rect 54686 34302 54738 34354
rect 10558 34190 10610 34242
rect 10782 34190 10834 34242
rect 14814 34190 14866 34242
rect 30270 34190 30322 34242
rect 30942 34190 30994 34242
rect 31390 34190 31442 34242
rect 34638 34190 34690 34242
rect 35982 34190 36034 34242
rect 37102 34190 37154 34242
rect 47182 34190 47234 34242
rect 54910 34190 54962 34242
rect 56702 34190 56754 34242
rect 8542 34078 8594 34130
rect 9886 34078 9938 34130
rect 11342 34078 11394 34130
rect 11790 34078 11842 34130
rect 12238 34078 12290 34130
rect 13918 34078 13970 34130
rect 17838 34078 17890 34130
rect 18286 34078 18338 34130
rect 19182 34078 19234 34130
rect 23886 34078 23938 34130
rect 28366 34078 28418 34130
rect 28702 34078 28754 34130
rect 28926 34078 28978 34130
rect 30382 34078 30434 34130
rect 30718 34078 30770 34130
rect 31838 34078 31890 34130
rect 34190 34078 34242 34130
rect 36542 34078 36594 34130
rect 36766 34078 36818 34130
rect 37438 34078 37490 34130
rect 38782 34078 38834 34130
rect 39230 34078 39282 34130
rect 40350 34078 40402 34130
rect 41022 34078 41074 34130
rect 41694 34078 41746 34130
rect 42030 34078 42082 34130
rect 43934 34078 43986 34130
rect 44606 34078 44658 34130
rect 45726 34078 45778 34130
rect 45950 34078 46002 34130
rect 55022 34078 55074 34130
rect 57038 34078 57090 34130
rect 57262 34078 57314 34130
rect 8878 33966 8930 34018
rect 14478 33966 14530 34018
rect 23550 33966 23602 34018
rect 25454 33966 25506 34018
rect 27582 33966 27634 34018
rect 28814 33966 28866 34018
rect 31614 33966 31666 34018
rect 33854 33966 33906 34018
rect 37326 33966 37378 34018
rect 38334 33966 38386 34018
rect 39678 33966 39730 34018
rect 41582 33966 41634 34018
rect 46622 33966 46674 34018
rect 46958 33966 47010 34018
rect 47294 33966 47346 34018
rect 47742 33966 47794 34018
rect 56814 33966 56866 34018
rect 9550 33854 9602 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 12798 33518 12850 33570
rect 57038 33518 57090 33570
rect 57598 33518 57650 33570
rect 13918 33406 13970 33458
rect 18062 33406 18114 33458
rect 24222 33406 24274 33458
rect 27918 33406 27970 33458
rect 51214 33406 51266 33458
rect 55582 33406 55634 33458
rect 11678 33294 11730 33346
rect 12238 33294 12290 33346
rect 12798 33294 12850 33346
rect 15150 33294 15202 33346
rect 18846 33294 18898 33346
rect 19630 33294 19682 33346
rect 20078 33294 20130 33346
rect 21422 33294 21474 33346
rect 22094 33294 22146 33346
rect 28142 33294 28194 33346
rect 28366 33294 28418 33346
rect 31278 33294 31330 33346
rect 31838 33294 31890 33346
rect 33630 33294 33682 33346
rect 34302 33294 34354 33346
rect 35086 33294 35138 33346
rect 36990 33294 37042 33346
rect 38446 33294 38498 33346
rect 38894 33294 38946 33346
rect 39790 33294 39842 33346
rect 40238 33294 40290 33346
rect 41246 33294 41298 33346
rect 41694 33294 41746 33346
rect 42030 33294 42082 33346
rect 42366 33294 42418 33346
rect 43934 33294 43986 33346
rect 48302 33294 48354 33346
rect 51886 33294 51938 33346
rect 52782 33294 52834 33346
rect 57486 33294 57538 33346
rect 15934 33182 15986 33234
rect 18510 33182 18562 33234
rect 18622 33182 18674 33234
rect 19070 33182 19122 33234
rect 25790 33182 25842 33234
rect 27806 33182 27858 33234
rect 32398 33182 32450 33234
rect 38110 33182 38162 33234
rect 39118 33182 39170 33234
rect 43710 33182 43762 33234
rect 49086 33182 49138 33234
rect 51550 33182 51602 33234
rect 51998 33182 52050 33234
rect 52110 33182 52162 33234
rect 53454 33182 53506 33234
rect 57150 33182 57202 33234
rect 13470 33070 13522 33122
rect 14814 33070 14866 33122
rect 19406 33070 19458 33122
rect 19518 33070 19570 33122
rect 20526 33070 20578 33122
rect 24670 33070 24722 33122
rect 25118 33070 25170 33122
rect 25454 33070 25506 33122
rect 27582 33070 27634 33122
rect 29486 33070 29538 33122
rect 30942 33070 30994 33122
rect 31502 33070 31554 33122
rect 36206 33070 36258 33122
rect 37102 33070 37154 33122
rect 42030 33070 42082 33122
rect 56030 33070 56082 33122
rect 57038 33070 57090 33122
rect 57598 33070 57650 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 8990 32734 9042 32786
rect 13134 32734 13186 32786
rect 18734 32734 18786 32786
rect 24110 32734 24162 32786
rect 24446 32734 24498 32786
rect 32062 32734 32114 32786
rect 34078 32734 34130 32786
rect 38110 32734 38162 32786
rect 39342 32734 39394 32786
rect 43374 32734 43426 32786
rect 49086 32734 49138 32786
rect 51774 32734 51826 32786
rect 53902 32734 53954 32786
rect 55134 32734 55186 32786
rect 11006 32622 11058 32674
rect 13022 32622 13074 32674
rect 50654 32622 50706 32674
rect 51998 32622 52050 32674
rect 52110 32622 52162 32674
rect 52894 32622 52946 32674
rect 53230 32622 53282 32674
rect 54014 32622 54066 32674
rect 54798 32622 54850 32674
rect 8766 32510 8818 32562
rect 9550 32510 9602 32562
rect 10894 32510 10946 32562
rect 11454 32510 11506 32562
rect 12462 32510 12514 32562
rect 12798 32510 12850 32562
rect 31726 32510 31778 32562
rect 31838 32510 31890 32562
rect 33966 32510 34018 32562
rect 34190 32510 34242 32562
rect 34974 32510 35026 32562
rect 37214 32510 37266 32562
rect 38446 32510 38498 32562
rect 39902 32510 39954 32562
rect 43934 32510 43986 32562
rect 44158 32510 44210 32562
rect 44494 32510 44546 32562
rect 44942 32510 44994 32562
rect 46734 32510 46786 32562
rect 47406 32510 47458 32562
rect 48974 32510 49026 32562
rect 49198 32510 49250 32562
rect 49646 32510 49698 32562
rect 50318 32510 50370 32562
rect 50430 32510 50482 32562
rect 50878 32510 50930 32562
rect 9886 32398 9938 32450
rect 18622 32398 18674 32450
rect 19406 32398 19458 32450
rect 20190 32398 20242 32450
rect 28590 32398 28642 32450
rect 31054 32398 31106 32450
rect 31502 32398 31554 32450
rect 34526 32398 34578 32450
rect 36878 32398 36930 32450
rect 37662 32398 37714 32450
rect 38894 32398 38946 32450
rect 43598 32398 43650 32450
rect 44046 32398 44098 32450
rect 46510 32398 46562 32450
rect 51438 32398 51490 32450
rect 58158 32398 58210 32450
rect 43262 32286 43314 32338
rect 53902 32286 53954 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 9326 31950 9378 32002
rect 10782 31950 10834 32002
rect 12238 31950 12290 32002
rect 35758 31950 35810 32002
rect 43710 31950 43762 32002
rect 44046 31950 44098 32002
rect 49870 31950 49922 32002
rect 8542 31838 8594 31890
rect 10334 31838 10386 31890
rect 14254 31838 14306 31890
rect 15038 31838 15090 31890
rect 18286 31838 18338 31890
rect 19070 31838 19122 31890
rect 26798 31838 26850 31890
rect 31838 31838 31890 31890
rect 34750 31838 34802 31890
rect 37102 31838 37154 31890
rect 37886 31838 37938 31890
rect 39566 31838 39618 31890
rect 41694 31838 41746 31890
rect 42142 31838 42194 31890
rect 45390 31838 45442 31890
rect 48750 31838 48802 31890
rect 56030 31838 56082 31890
rect 58158 31838 58210 31890
rect 8430 31726 8482 31778
rect 10446 31726 10498 31778
rect 11342 31726 11394 31778
rect 13470 31726 13522 31778
rect 14030 31726 14082 31778
rect 15374 31726 15426 31778
rect 18622 31726 18674 31778
rect 23886 31726 23938 31778
rect 32062 31726 32114 31778
rect 34190 31726 34242 31778
rect 34302 31726 34354 31778
rect 35422 31726 35474 31778
rect 37550 31726 37602 31778
rect 37998 31726 38050 31778
rect 38894 31726 38946 31778
rect 44270 31726 44322 31778
rect 48302 31726 48354 31778
rect 49310 31726 49362 31778
rect 49534 31726 49586 31778
rect 50094 31726 50146 31778
rect 55246 31726 55298 31778
rect 8094 31614 8146 31666
rect 8654 31614 8706 31666
rect 8990 31614 9042 31666
rect 12574 31614 12626 31666
rect 14142 31614 14194 31666
rect 16158 31614 16210 31666
rect 24670 31614 24722 31666
rect 33070 31614 33122 31666
rect 35198 31614 35250 31666
rect 47518 31614 47570 31666
rect 49422 31614 49474 31666
rect 9214 31502 9266 31554
rect 12350 31502 12402 31554
rect 27246 31502 27298 31554
rect 32062 31502 32114 31554
rect 50430 31502 50482 31554
rect 50766 31502 50818 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 9886 31166 9938 31218
rect 12462 31166 12514 31218
rect 22766 31166 22818 31218
rect 23326 31166 23378 31218
rect 24110 31166 24162 31218
rect 31054 31166 31106 31218
rect 32062 31166 32114 31218
rect 34862 31166 34914 31218
rect 35870 31166 35922 31218
rect 49086 31166 49138 31218
rect 56926 31166 56978 31218
rect 13470 31054 13522 31106
rect 21982 31054 22034 31106
rect 22094 31054 22146 31106
rect 22206 31054 22258 31106
rect 35310 31054 35362 31106
rect 43038 31054 43090 31106
rect 49982 31054 50034 31106
rect 55358 31054 55410 31106
rect 57822 31054 57874 31106
rect 58158 31054 58210 31106
rect 7646 30942 7698 30994
rect 8542 30942 8594 30994
rect 8878 30942 8930 30994
rect 9886 30942 9938 30994
rect 10222 30942 10274 30994
rect 11454 30942 11506 30994
rect 12910 30942 12962 30994
rect 21534 30942 21586 30994
rect 22318 30942 22370 30994
rect 22542 30942 22594 30994
rect 22878 30942 22930 30994
rect 23102 30942 23154 30994
rect 23438 30942 23490 30994
rect 23998 30942 24050 30994
rect 24334 30942 24386 30994
rect 28142 30942 28194 30994
rect 42366 30942 42418 30994
rect 55134 30942 55186 30994
rect 56590 30942 56642 30994
rect 56814 30942 56866 30994
rect 57262 30942 57314 30994
rect 8206 30830 8258 30882
rect 9774 30830 9826 30882
rect 11118 30830 11170 30882
rect 12686 30830 12738 30882
rect 21198 30830 21250 30882
rect 25454 30830 25506 30882
rect 27694 30830 27746 30882
rect 28814 30830 28866 30882
rect 31614 30830 31666 30882
rect 45166 30830 45218 30882
rect 45614 30830 45666 30882
rect 49870 30830 49922 30882
rect 50206 30830 50258 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 46510 30382 46562 30434
rect 9214 30270 9266 30322
rect 11118 30270 11170 30322
rect 19182 30270 19234 30322
rect 21534 30270 21586 30322
rect 25006 30270 25058 30322
rect 28590 30270 28642 30322
rect 29150 30270 29202 30322
rect 39902 30270 39954 30322
rect 46958 30270 47010 30322
rect 56030 30270 56082 30322
rect 58158 30270 58210 30322
rect 8990 30158 9042 30210
rect 12910 30158 12962 30210
rect 13582 30158 13634 30210
rect 13806 30158 13858 30210
rect 14142 30158 14194 30210
rect 14814 30158 14866 30210
rect 19630 30158 19682 30210
rect 22318 30158 22370 30210
rect 25790 30158 25842 30210
rect 30158 30158 30210 30210
rect 34078 30158 34130 30210
rect 34638 30158 34690 30210
rect 37102 30158 37154 30210
rect 46622 30158 46674 30210
rect 49870 30158 49922 30210
rect 50206 30158 50258 30210
rect 50878 30158 50930 30210
rect 51550 30158 51602 30210
rect 52670 30158 52722 30210
rect 55358 30158 55410 30210
rect 7982 30046 8034 30098
rect 9774 30046 9826 30098
rect 11902 30046 11954 30098
rect 21758 30046 21810 30098
rect 21982 30046 22034 30098
rect 22094 30046 22146 30098
rect 24222 30046 24274 30098
rect 24558 30046 24610 30098
rect 24782 30046 24834 30098
rect 26462 30046 26514 30098
rect 29486 30046 29538 30098
rect 29598 30046 29650 30098
rect 30382 30046 30434 30098
rect 30494 30046 30546 30098
rect 31278 30046 31330 30098
rect 35422 30046 35474 30098
rect 37774 30046 37826 30098
rect 49086 30046 49138 30098
rect 50318 30046 50370 30098
rect 51774 30046 51826 30098
rect 12798 29934 12850 29986
rect 15598 29934 15650 29986
rect 22878 29934 22930 29986
rect 24446 29934 24498 29986
rect 29710 29934 29762 29986
rect 29934 29934 29986 29986
rect 31390 29934 31442 29986
rect 31614 29934 31666 29986
rect 35086 29934 35138 29986
rect 35758 29934 35810 29986
rect 40350 29934 40402 29986
rect 46510 29934 46562 29986
rect 50542 29934 50594 29986
rect 53006 29934 53058 29986
rect 54574 29934 54626 29986
rect 54910 29934 54962 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 16606 29598 16658 29650
rect 17502 29598 17554 29650
rect 18062 29598 18114 29650
rect 21870 29598 21922 29650
rect 22318 29598 22370 29650
rect 22878 29598 22930 29650
rect 23214 29598 23266 29650
rect 24334 29598 24386 29650
rect 25566 29598 25618 29650
rect 26910 29598 26962 29650
rect 27806 29598 27858 29650
rect 28702 29598 28754 29650
rect 30830 29598 30882 29650
rect 31838 29598 31890 29650
rect 37214 29598 37266 29650
rect 42926 29598 42978 29650
rect 43486 29598 43538 29650
rect 51102 29598 51154 29650
rect 53118 29598 53170 29650
rect 56702 29598 56754 29650
rect 56926 29598 56978 29650
rect 57822 29598 57874 29650
rect 8990 29486 9042 29538
rect 14814 29486 14866 29538
rect 16494 29486 16546 29538
rect 17278 29486 17330 29538
rect 21534 29486 21586 29538
rect 21646 29486 21698 29538
rect 22094 29486 22146 29538
rect 22430 29486 22482 29538
rect 23662 29486 23714 29538
rect 25230 29486 25282 29538
rect 27582 29486 27634 29538
rect 27694 29486 27746 29538
rect 28478 29486 28530 29538
rect 31166 29486 31218 29538
rect 36990 29486 37042 29538
rect 51550 29486 51602 29538
rect 53454 29486 53506 29538
rect 57038 29486 57090 29538
rect 4398 29374 4450 29426
rect 8318 29374 8370 29426
rect 8766 29374 8818 29426
rect 11230 29374 11282 29426
rect 12014 29374 12066 29426
rect 13022 29374 13074 29426
rect 14254 29374 14306 29426
rect 14590 29374 14642 29426
rect 15038 29374 15090 29426
rect 15374 29374 15426 29426
rect 16046 29374 16098 29426
rect 16830 29374 16882 29426
rect 17614 29374 17666 29426
rect 21086 29374 21138 29426
rect 23998 29374 24050 29426
rect 24558 29374 24610 29426
rect 28030 29374 28082 29426
rect 28814 29374 28866 29426
rect 30606 29374 30658 29426
rect 31054 29374 31106 29426
rect 35646 29374 35698 29426
rect 36878 29374 36930 29426
rect 37438 29374 37490 29426
rect 50990 29374 51042 29426
rect 51214 29374 51266 29426
rect 5070 29262 5122 29314
rect 7198 29262 7250 29314
rect 7870 29262 7922 29314
rect 10446 29262 10498 29314
rect 13918 29262 13970 29314
rect 14702 29262 14754 29314
rect 16494 29262 16546 29314
rect 20750 29262 20802 29314
rect 21534 29262 21586 29314
rect 27694 29262 27746 29314
rect 29262 29262 29314 29314
rect 29710 29262 29762 29314
rect 31390 29262 31442 29314
rect 35982 29262 36034 29314
rect 40238 29262 40290 29314
rect 44046 29262 44098 29314
rect 53902 29262 53954 29314
rect 58158 29262 58210 29314
rect 40126 29150 40178 29202
rect 42814 29150 42866 29202
rect 43150 29150 43202 29202
rect 43822 29150 43874 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 12014 28814 12066 28866
rect 29038 28814 29090 28866
rect 29374 28814 29426 28866
rect 8094 28702 8146 28754
rect 9998 28702 10050 28754
rect 15934 28702 15986 28754
rect 19630 28702 19682 28754
rect 29374 28702 29426 28754
rect 31950 28702 32002 28754
rect 34078 28702 34130 28754
rect 34862 28702 34914 28754
rect 36430 28702 36482 28754
rect 37886 28702 37938 28754
rect 41470 28702 41522 28754
rect 41918 28702 41970 28754
rect 43486 28702 43538 28754
rect 45278 28702 45330 28754
rect 48526 28702 48578 28754
rect 49534 28702 49586 28754
rect 49758 28702 49810 28754
rect 50654 28702 50706 28754
rect 56590 28702 56642 28754
rect 7646 28590 7698 28642
rect 9326 28590 9378 28642
rect 11006 28590 11058 28642
rect 12350 28590 12402 28642
rect 13918 28590 13970 28642
rect 14702 28590 14754 28642
rect 15150 28590 15202 28642
rect 16830 28590 16882 28642
rect 28142 28590 28194 28642
rect 30270 28590 30322 28642
rect 30606 28590 30658 28642
rect 30942 28590 30994 28642
rect 31166 28590 31218 28642
rect 35310 28590 35362 28642
rect 35870 28590 35922 28642
rect 37326 28590 37378 28642
rect 38670 28590 38722 28642
rect 42702 28590 42754 28642
rect 42926 28590 42978 28642
rect 45614 28590 45666 28642
rect 52670 28590 52722 28642
rect 53230 28590 53282 28642
rect 54462 28590 54514 28642
rect 10446 28478 10498 28530
rect 12574 28478 12626 28530
rect 14142 28478 14194 28530
rect 14254 28478 14306 28530
rect 16158 28478 16210 28530
rect 16270 28478 16322 28530
rect 17502 28478 17554 28530
rect 28366 28478 28418 28530
rect 30718 28478 30770 28530
rect 37774 28478 37826 28530
rect 39342 28478 39394 28530
rect 46398 28478 46450 28530
rect 53006 28478 53058 28530
rect 53566 28478 53618 28530
rect 7198 28366 7250 28418
rect 14030 28366 14082 28418
rect 16494 28366 16546 28418
rect 34414 28366 34466 28418
rect 37102 28366 37154 28418
rect 37998 28366 38050 28418
rect 43374 28366 43426 28418
rect 43598 28366 43650 28418
rect 50094 28366 50146 28418
rect 53454 28366 53506 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 11454 28030 11506 28082
rect 11790 28030 11842 28082
rect 12798 28030 12850 28082
rect 14142 28030 14194 28082
rect 14926 28030 14978 28082
rect 16382 28030 16434 28082
rect 17390 28030 17442 28082
rect 17502 28030 17554 28082
rect 18846 28030 18898 28082
rect 19182 28030 19234 28082
rect 28478 28030 28530 28082
rect 28926 28030 28978 28082
rect 30830 28030 30882 28082
rect 34526 28030 34578 28082
rect 36094 28030 36146 28082
rect 38894 28030 38946 28082
rect 44382 28030 44434 28082
rect 54686 28030 54738 28082
rect 56590 28030 56642 28082
rect 57374 28030 57426 28082
rect 5518 27918 5570 27970
rect 10446 27918 10498 27970
rect 14366 27918 14418 27970
rect 17614 27918 17666 27970
rect 17726 27918 17778 27970
rect 20302 27918 20354 27970
rect 31054 27918 31106 27970
rect 32062 27918 32114 27970
rect 38110 27918 38162 27970
rect 38222 27918 38274 27970
rect 38446 27918 38498 27970
rect 39006 27918 39058 27970
rect 39118 27918 39170 27970
rect 41806 27918 41858 27970
rect 55470 27918 55522 27970
rect 56926 27918 56978 27970
rect 57262 27918 57314 27970
rect 57934 27918 57986 27970
rect 4846 27806 4898 27858
rect 8094 27806 8146 27858
rect 9550 27806 9602 27858
rect 10894 27806 10946 27858
rect 11342 27806 11394 27858
rect 12686 27806 12738 27858
rect 12910 27806 12962 27858
rect 14478 27806 14530 27858
rect 14814 27806 14866 27858
rect 18174 27806 18226 27858
rect 19630 27806 19682 27858
rect 22878 27806 22930 27858
rect 25790 27806 25842 27858
rect 28142 27806 28194 27858
rect 31278 27806 31330 27858
rect 31502 27806 31554 27858
rect 32510 27806 32562 27858
rect 35758 27806 35810 27858
rect 38670 27806 38722 27858
rect 41134 27806 41186 27858
rect 51438 27806 51490 27858
rect 55134 27806 55186 27858
rect 57822 27806 57874 27858
rect 7646 27694 7698 27746
rect 9998 27694 10050 27746
rect 12350 27694 12402 27746
rect 22430 27694 22482 27746
rect 26350 27694 26402 27746
rect 31614 27694 31666 27746
rect 34974 27694 35026 27746
rect 37774 27694 37826 27746
rect 39454 27694 39506 27746
rect 43934 27694 43986 27746
rect 52110 27694 52162 27746
rect 54238 27694 54290 27746
rect 14926 27582 14978 27634
rect 57374 27582 57426 27634
rect 57934 27582 57986 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 24558 27246 24610 27298
rect 26686 27246 26738 27298
rect 9662 27134 9714 27186
rect 12462 27134 12514 27186
rect 18174 27134 18226 27186
rect 18622 27134 18674 27186
rect 19518 27134 19570 27186
rect 31726 27134 31778 27186
rect 33854 27134 33906 27186
rect 41918 27134 41970 27186
rect 52782 27134 52834 27186
rect 58158 27134 58210 27186
rect 12910 27022 12962 27074
rect 14142 27022 14194 27074
rect 14926 27022 14978 27074
rect 26014 27022 26066 27074
rect 26238 27022 26290 27074
rect 30606 27022 30658 27074
rect 30942 27022 30994 27074
rect 37998 27022 38050 27074
rect 40014 27022 40066 27074
rect 40910 27022 40962 27074
rect 52558 27022 52610 27074
rect 53230 27022 53282 27074
rect 53790 27022 53842 27074
rect 55358 27022 55410 27074
rect 9214 26910 9266 26962
rect 13470 26910 13522 26962
rect 13806 26910 13858 26962
rect 14254 26910 14306 26962
rect 24670 26910 24722 26962
rect 25790 26910 25842 26962
rect 26574 26910 26626 26962
rect 29374 26910 29426 26962
rect 38222 26910 38274 26962
rect 38670 26910 38722 26962
rect 44270 26910 44322 26962
rect 44830 26910 44882 26962
rect 45166 26910 45218 26962
rect 45390 26910 45442 26962
rect 53006 26910 53058 26962
rect 53454 26910 53506 26962
rect 56030 26910 56082 26962
rect 8878 26798 8930 26850
rect 14478 26798 14530 26850
rect 14590 26798 14642 26850
rect 14814 26798 14866 26850
rect 24558 26798 24610 26850
rect 25566 26798 25618 26850
rect 25678 26798 25730 26850
rect 26686 26798 26738 26850
rect 28590 26798 28642 26850
rect 29822 26798 29874 26850
rect 43934 26798 43986 26850
rect 44158 26798 44210 26850
rect 44942 26798 44994 26850
rect 53678 26798 53730 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 9774 26462 9826 26514
rect 10670 26462 10722 26514
rect 16494 26462 16546 26514
rect 22318 26462 22370 26514
rect 22654 26462 22706 26514
rect 25342 26462 25394 26514
rect 26462 26462 26514 26514
rect 27358 26462 27410 26514
rect 28478 26462 28530 26514
rect 29038 26462 29090 26514
rect 30270 26462 30322 26514
rect 30830 26462 30882 26514
rect 34414 26462 34466 26514
rect 39230 26462 39282 26514
rect 52334 26462 52386 26514
rect 57038 26462 57090 26514
rect 15598 26350 15650 26402
rect 15934 26350 15986 26402
rect 17390 26350 17442 26402
rect 18174 26350 18226 26402
rect 18622 26350 18674 26402
rect 25118 26350 25170 26402
rect 25454 26350 25506 26402
rect 28814 26350 28866 26402
rect 29598 26350 29650 26402
rect 33966 26350 34018 26402
rect 39790 26350 39842 26402
rect 41470 26350 41522 26402
rect 52558 26350 52610 26402
rect 52670 26350 52722 26402
rect 6078 26238 6130 26290
rect 9550 26238 9602 26290
rect 10222 26238 10274 26290
rect 11790 26238 11842 26290
rect 13246 26238 13298 26290
rect 16830 26238 16882 26290
rect 17726 26238 17778 26290
rect 18062 26238 18114 26290
rect 19182 26238 19234 26290
rect 23774 26238 23826 26290
rect 24222 26238 24274 26290
rect 26350 26238 26402 26290
rect 26574 26238 26626 26290
rect 27134 26238 27186 26290
rect 27470 26238 27522 26290
rect 28254 26238 28306 26290
rect 28590 26238 28642 26290
rect 29150 26238 29202 26290
rect 30158 26238 30210 26290
rect 39454 26238 39506 26290
rect 40126 26238 40178 26290
rect 41134 26238 41186 26290
rect 42590 26238 42642 26290
rect 47630 26238 47682 26290
rect 48190 26238 48242 26290
rect 56590 26238 56642 26290
rect 56926 26238 56978 26290
rect 57262 26238 57314 26290
rect 6750 26126 6802 26178
rect 8878 26126 8930 26178
rect 9662 26126 9714 26178
rect 11006 26126 11058 26178
rect 12238 26126 12290 26178
rect 13918 26126 13970 26178
rect 23214 26126 23266 26178
rect 24334 26126 24386 26178
rect 26126 26126 26178 26178
rect 27246 26126 27298 26178
rect 36766 26126 36818 26178
rect 37662 26126 37714 26178
rect 41918 26126 41970 26178
rect 43262 26126 43314 26178
rect 45390 26126 45442 26178
rect 58158 26126 58210 26178
rect 18174 26014 18226 26066
rect 25902 26014 25954 26066
rect 27806 26014 27858 26066
rect 29486 26014 29538 26066
rect 30270 26014 30322 26066
rect 33854 26014 33906 26066
rect 39118 26014 39170 26066
rect 41022 26014 41074 26066
rect 41358 26014 41410 26066
rect 47294 26014 47346 26066
rect 47630 26014 47682 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 24670 25678 24722 25730
rect 27694 25678 27746 25730
rect 39790 25678 39842 25730
rect 39902 25678 39954 25730
rect 40686 25678 40738 25730
rect 43598 25678 43650 25730
rect 43934 25678 43986 25730
rect 44046 25678 44098 25730
rect 8318 25566 8370 25618
rect 9438 25566 9490 25618
rect 15486 25566 15538 25618
rect 15934 25566 15986 25618
rect 19742 25566 19794 25618
rect 23326 25566 23378 25618
rect 26126 25566 26178 25618
rect 27806 25566 27858 25618
rect 28590 25566 28642 25618
rect 33854 25566 33906 25618
rect 34190 25566 34242 25618
rect 36206 25566 36258 25618
rect 38334 25566 38386 25618
rect 39006 25566 39058 25618
rect 39342 25566 39394 25618
rect 45054 25566 45106 25618
rect 46622 25566 46674 25618
rect 46958 25566 47010 25618
rect 49086 25566 49138 25618
rect 50318 25566 50370 25618
rect 8542 25454 8594 25506
rect 8766 25454 8818 25506
rect 12238 25454 12290 25506
rect 12798 25454 12850 25506
rect 16270 25454 16322 25506
rect 16830 25454 16882 25506
rect 21422 25454 21474 25506
rect 23886 25454 23938 25506
rect 24222 25454 24274 25506
rect 25566 25454 25618 25506
rect 25902 25454 25954 25506
rect 26014 25454 26066 25506
rect 26910 25454 26962 25506
rect 29150 25454 29202 25506
rect 32398 25454 32450 25506
rect 32734 25454 32786 25506
rect 33294 25454 33346 25506
rect 34974 25454 35026 25506
rect 36990 25454 37042 25506
rect 37214 25454 37266 25506
rect 37550 25454 37602 25506
rect 38446 25454 38498 25506
rect 40126 25454 40178 25506
rect 41918 25454 41970 25506
rect 43710 25454 43762 25506
rect 45726 25454 45778 25506
rect 45950 25454 46002 25506
rect 49870 25454 49922 25506
rect 52558 25454 52610 25506
rect 53006 25454 53058 25506
rect 53118 25454 53170 25506
rect 53454 25454 53506 25506
rect 53790 25454 53842 25506
rect 8206 25342 8258 25394
rect 11566 25342 11618 25394
rect 14030 25342 14082 25394
rect 14254 25342 14306 25394
rect 14478 25342 14530 25394
rect 17614 25342 17666 25394
rect 21758 25342 21810 25394
rect 21982 25342 22034 25394
rect 24110 25342 24162 25394
rect 24558 25342 24610 25394
rect 26686 25342 26738 25394
rect 27358 25342 27410 25394
rect 29486 25342 29538 25394
rect 30942 25342 30994 25394
rect 32622 25342 32674 25394
rect 32958 25342 33010 25394
rect 34638 25342 34690 25394
rect 35422 25342 35474 25394
rect 39230 25342 39282 25394
rect 40238 25342 40290 25394
rect 40574 25342 40626 25394
rect 40686 25342 40738 25394
rect 41470 25342 41522 25394
rect 44830 25342 44882 25394
rect 45054 25342 45106 25394
rect 45278 25342 45330 25394
rect 56590 25342 56642 25394
rect 56702 25342 56754 25394
rect 58158 25342 58210 25394
rect 13918 25230 13970 25282
rect 14142 25230 14194 25282
rect 16382 25230 16434 25282
rect 16606 25230 16658 25282
rect 21534 25230 21586 25282
rect 22542 25230 22594 25282
rect 26238 25230 26290 25282
rect 29710 25230 29762 25282
rect 31278 25230 31330 25282
rect 33182 25230 33234 25282
rect 34078 25230 34130 25282
rect 35758 25230 35810 25282
rect 37102 25230 37154 25282
rect 37998 25230 38050 25282
rect 38222 25230 38274 25282
rect 41694 25230 41746 25282
rect 42478 25230 42530 25282
rect 42926 25230 42978 25282
rect 52782 25230 52834 25282
rect 53678 25230 53730 25282
rect 56366 25230 56418 25282
rect 57598 25230 57650 25282
rect 57822 25230 57874 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 8990 24894 9042 24946
rect 13358 24894 13410 24946
rect 13918 24894 13970 24946
rect 15150 24894 15202 24946
rect 16046 24894 16098 24946
rect 17390 24894 17442 24946
rect 17502 24894 17554 24946
rect 19070 24894 19122 24946
rect 25566 24894 25618 24946
rect 28142 24894 28194 24946
rect 29934 24894 29986 24946
rect 31390 24894 31442 24946
rect 39230 24894 39282 24946
rect 44382 24894 44434 24946
rect 45838 24894 45890 24946
rect 52558 24894 52610 24946
rect 14142 24782 14194 24834
rect 14478 24782 14530 24834
rect 16270 24782 16322 24834
rect 17614 24782 17666 24834
rect 18622 24782 18674 24834
rect 20526 24782 20578 24834
rect 25342 24782 25394 24834
rect 27694 24782 27746 24834
rect 28926 24782 28978 24834
rect 36094 24782 36146 24834
rect 40910 24782 40962 24834
rect 41134 24782 41186 24834
rect 42142 24782 42194 24834
rect 50206 24782 50258 24834
rect 52782 24782 52834 24834
rect 52894 24782 52946 24834
rect 53342 24838 53394 24890
rect 56814 24894 56866 24946
rect 53454 24782 53506 24834
rect 57822 24782 57874 24834
rect 10110 24670 10162 24722
rect 14366 24670 14418 24722
rect 16494 24670 16546 24722
rect 16718 24670 16770 24722
rect 17838 24670 17890 24722
rect 18062 24670 18114 24722
rect 19742 24670 19794 24722
rect 23438 24670 23490 24722
rect 25230 24670 25282 24722
rect 27470 24670 27522 24722
rect 28702 24670 28754 24722
rect 29150 24670 29202 24722
rect 29486 24670 29538 24722
rect 32958 24670 33010 24722
rect 33294 24670 33346 24722
rect 33630 24670 33682 24722
rect 34190 24670 34242 24722
rect 35422 24670 35474 24722
rect 42702 24670 42754 24722
rect 43038 24670 43090 24722
rect 49534 24670 49586 24722
rect 56478 24670 56530 24722
rect 56926 24670 56978 24722
rect 57150 24670 57202 24722
rect 10782 24558 10834 24610
rect 12910 24558 12962 24610
rect 14030 24558 14082 24610
rect 15598 24558 15650 24610
rect 16158 24558 16210 24610
rect 22654 24558 22706 24610
rect 22990 24558 23042 24610
rect 23998 24558 24050 24610
rect 29038 24558 29090 24610
rect 31838 24558 31890 24610
rect 38222 24558 38274 24610
rect 38670 24558 38722 24610
rect 41022 24558 41074 24610
rect 41806 24558 41858 24610
rect 43486 24558 43538 24610
rect 44830 24558 44882 24610
rect 45278 24558 45330 24610
rect 52334 24558 52386 24610
rect 53902 24558 53954 24610
rect 57486 24558 57538 24610
rect 27134 24446 27186 24498
rect 53342 24446 53394 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 31502 24110 31554 24162
rect 17838 23998 17890 24050
rect 19406 23998 19458 24050
rect 22318 23998 22370 24050
rect 27694 23998 27746 24050
rect 29150 23998 29202 24050
rect 38446 23998 38498 24050
rect 45166 23998 45218 24050
rect 55134 23998 55186 24050
rect 57262 23998 57314 24050
rect 18958 23886 19010 23938
rect 19854 23886 19906 23938
rect 20302 23886 20354 23938
rect 22206 23886 22258 23938
rect 24894 23886 24946 23938
rect 26910 23886 26962 23938
rect 27918 23886 27970 23938
rect 33742 23886 33794 23938
rect 35758 23886 35810 23938
rect 45502 23886 45554 23938
rect 46062 23886 46114 23938
rect 52782 23886 52834 23938
rect 53006 23886 53058 23938
rect 53342 23886 53394 23938
rect 53790 23886 53842 23938
rect 58046 23886 58098 23938
rect 17278 23774 17330 23826
rect 24334 23774 24386 23826
rect 26350 23774 26402 23826
rect 28254 23774 28306 23826
rect 31614 23774 31666 23826
rect 32062 23774 32114 23826
rect 35982 23774 36034 23826
rect 20750 23662 20802 23714
rect 21982 23662 22034 23714
rect 22430 23662 22482 23714
rect 22654 23662 22706 23714
rect 26798 23662 26850 23714
rect 29262 23662 29314 23714
rect 33406 23662 33458 23714
rect 45838 23662 45890 23714
rect 46510 23662 46562 23714
rect 46622 23662 46674 23714
rect 46734 23662 46786 23714
rect 53006 23662 53058 23714
rect 53454 23662 53506 23714
rect 53678 23662 53730 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 23438 23326 23490 23378
rect 25342 23326 25394 23378
rect 25566 23326 25618 23378
rect 25790 23326 25842 23378
rect 27582 23326 27634 23378
rect 33630 23326 33682 23378
rect 34078 23326 34130 23378
rect 41022 23326 41074 23378
rect 41806 23326 41858 23378
rect 42030 23326 42082 23378
rect 42478 23326 42530 23378
rect 43374 23326 43426 23378
rect 44158 23326 44210 23378
rect 44606 23326 44658 23378
rect 56702 23326 56754 23378
rect 56926 23326 56978 23378
rect 16046 23214 16098 23266
rect 22766 23214 22818 23266
rect 24334 23214 24386 23266
rect 25230 23214 25282 23266
rect 30046 23214 30098 23266
rect 39230 23214 39282 23266
rect 44942 23214 44994 23266
rect 51438 23214 51490 23266
rect 54126 23214 54178 23266
rect 54350 23214 54402 23266
rect 56590 23214 56642 23266
rect 16830 23102 16882 23154
rect 17502 23102 17554 23154
rect 22318 23102 22370 23154
rect 22990 23102 23042 23154
rect 23662 23102 23714 23154
rect 24110 23102 24162 23154
rect 24222 23102 24274 23154
rect 25902 23102 25954 23154
rect 30718 23102 30770 23154
rect 38110 23102 38162 23154
rect 38446 23102 38498 23154
rect 38782 23102 38834 23154
rect 42254 23102 42306 23154
rect 45278 23102 45330 23154
rect 50766 23102 50818 23154
rect 54014 23102 54066 23154
rect 13918 22990 13970 23042
rect 19742 22990 19794 23042
rect 22542 22990 22594 23042
rect 27918 22990 27970 23042
rect 33070 22990 33122 23042
rect 38334 22990 38386 23042
rect 42142 22990 42194 23042
rect 43710 22990 43762 23042
rect 46062 22990 46114 23042
rect 48190 22990 48242 23042
rect 53566 22990 53618 23042
rect 54686 22990 54738 23042
rect 58158 22990 58210 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 33182 22430 33234 22482
rect 36430 22430 36482 22482
rect 40686 22430 40738 22482
rect 44158 22430 44210 22482
rect 45054 22430 45106 22482
rect 45502 22430 45554 22482
rect 45838 22430 45890 22482
rect 47518 22430 47570 22482
rect 50766 22430 50818 22482
rect 51214 22430 51266 22482
rect 24446 22318 24498 22370
rect 26462 22318 26514 22370
rect 26910 22318 26962 22370
rect 33518 22318 33570 22370
rect 37886 22318 37938 22370
rect 38558 22318 38610 22370
rect 41246 22318 41298 22370
rect 45614 22318 45666 22370
rect 45950 22318 46002 22370
rect 46286 22318 46338 22370
rect 46734 22318 46786 22370
rect 47966 22318 48018 22370
rect 54910 22318 54962 22370
rect 56814 22318 56866 22370
rect 57374 22318 57426 22370
rect 57934 22318 57986 22370
rect 23886 22206 23938 22258
rect 25342 22206 25394 22258
rect 27918 22206 27970 22258
rect 34302 22206 34354 22258
rect 37214 22206 37266 22258
rect 37326 22206 37378 22258
rect 37438 22206 37490 22258
rect 42030 22206 42082 22258
rect 47070 22206 47122 22258
rect 47182 22206 47234 22258
rect 48638 22206 48690 22258
rect 54574 22206 54626 22258
rect 55134 22206 55186 22258
rect 56702 22206 56754 22258
rect 57038 22206 57090 22258
rect 28478 22094 28530 22146
rect 46958 22094 47010 22146
rect 54686 22094 54738 22146
rect 56478 22094 56530 22146
rect 57262 22094 57314 22146
rect 57598 22094 57650 22146
rect 57822 22094 57874 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 18622 21758 18674 21810
rect 19294 21758 19346 21810
rect 19966 21758 20018 21810
rect 25342 21758 25394 21810
rect 33630 21758 33682 21810
rect 34414 21758 34466 21810
rect 35534 21758 35586 21810
rect 36766 21758 36818 21810
rect 40350 21758 40402 21810
rect 41470 21758 41522 21810
rect 46398 21758 46450 21810
rect 47070 21758 47122 21810
rect 47294 21758 47346 21810
rect 49646 21758 49698 21810
rect 18286 21646 18338 21698
rect 18958 21646 19010 21698
rect 19630 21646 19682 21698
rect 22430 21646 22482 21698
rect 26350 21646 26402 21698
rect 27806 21646 27858 21698
rect 33966 21646 34018 21698
rect 36094 21646 36146 21698
rect 37102 21646 37154 21698
rect 38110 21646 38162 21698
rect 41806 21646 41858 21698
rect 49758 21646 49810 21698
rect 54350 21646 54402 21698
rect 56926 21646 56978 21698
rect 57150 21646 57202 21698
rect 21758 21534 21810 21586
rect 26798 21534 26850 21586
rect 27246 21534 27298 21586
rect 34190 21534 34242 21586
rect 34526 21534 34578 21586
rect 34862 21534 34914 21586
rect 35086 21534 35138 21586
rect 35646 21534 35698 21586
rect 35758 21534 35810 21586
rect 36318 21534 36370 21586
rect 38334 21534 38386 21586
rect 39006 21534 39058 21586
rect 41134 21534 41186 21586
rect 41470 21534 41522 21586
rect 47406 21534 47458 21586
rect 55134 21534 55186 21586
rect 55582 21534 55634 21586
rect 56478 21534 56530 21586
rect 24558 21422 24610 21474
rect 37774 21422 37826 21474
rect 45390 21422 45442 21474
rect 47854 21422 47906 21474
rect 52222 21422 52274 21474
rect 56702 21422 56754 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 14702 20862 14754 20914
rect 17950 20862 18002 20914
rect 19294 20862 19346 20914
rect 24894 20862 24946 20914
rect 30158 20862 30210 20914
rect 33518 20862 33570 20914
rect 56030 20862 56082 20914
rect 58158 20862 58210 20914
rect 15038 20750 15090 20802
rect 18286 20750 18338 20802
rect 18622 20750 18674 20802
rect 18734 20750 18786 20802
rect 20078 20750 20130 20802
rect 20526 20750 20578 20802
rect 22542 20750 22594 20802
rect 22878 20750 22930 20802
rect 28030 20750 28082 20802
rect 29038 20750 29090 20802
rect 29374 20750 29426 20802
rect 30718 20750 30770 20802
rect 33966 20750 34018 20802
rect 55246 20750 55298 20802
rect 15822 20638 15874 20690
rect 18398 20638 18450 20690
rect 20750 20638 20802 20690
rect 21982 20638 22034 20690
rect 29710 20638 29762 20690
rect 31390 20638 31442 20690
rect 20302 20526 20354 20578
rect 21870 20526 21922 20578
rect 22094 20526 22146 20578
rect 28254 20526 28306 20578
rect 29262 20526 29314 20578
rect 41582 20526 41634 20578
rect 47294 20526 47346 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 18510 20190 18562 20242
rect 31278 20190 31330 20242
rect 58158 20190 58210 20242
rect 18062 20078 18114 20130
rect 18398 20078 18450 20130
rect 20190 20078 20242 20130
rect 26798 20078 26850 20130
rect 27470 20078 27522 20130
rect 31614 20078 31666 20130
rect 32062 20078 32114 20130
rect 32398 20078 32450 20130
rect 40350 20078 40402 20130
rect 41246 20078 41298 20130
rect 46622 20078 46674 20130
rect 47966 20078 48018 20130
rect 18622 19966 18674 20018
rect 18958 19966 19010 20018
rect 19406 19966 19458 20018
rect 26574 19966 26626 20018
rect 27246 19966 27298 20018
rect 27918 19966 27970 20018
rect 28590 19966 28642 20018
rect 31054 19966 31106 20018
rect 31390 19966 31442 20018
rect 31950 19966 32002 20018
rect 32174 19966 32226 20018
rect 40910 19966 40962 20018
rect 41470 19966 41522 20018
rect 41806 19966 41858 20018
rect 46846 19966 46898 20018
rect 47070 19966 47122 20018
rect 47518 19966 47570 20018
rect 47742 19966 47794 20018
rect 22318 19854 22370 19906
rect 30718 19854 30770 19906
rect 37774 19854 37826 19906
rect 41022 19854 41074 19906
rect 42590 19854 42642 19906
rect 44718 19854 44770 19906
rect 46286 19854 46338 19906
rect 46734 19854 46786 19906
rect 47630 19854 47682 19906
rect 50318 19854 50370 19906
rect 51214 19854 51266 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 17278 19294 17330 19346
rect 17838 19294 17890 19346
rect 26238 19294 26290 19346
rect 30046 19294 30098 19346
rect 39790 19294 39842 19346
rect 42142 19294 42194 19346
rect 47854 19294 47906 19346
rect 49982 19294 50034 19346
rect 14478 19182 14530 19234
rect 18286 19182 18338 19234
rect 18958 19182 19010 19234
rect 23662 19182 23714 19234
rect 24334 19182 24386 19234
rect 26574 19182 26626 19234
rect 26798 19182 26850 19234
rect 33742 19182 33794 19234
rect 34302 19182 34354 19234
rect 36990 19182 37042 19234
rect 37214 19182 37266 19234
rect 37550 19182 37602 19234
rect 37998 19182 38050 19234
rect 38782 19182 38834 19234
rect 39118 19182 39170 19234
rect 42254 19182 42306 19234
rect 45614 19182 45666 19234
rect 46174 19182 46226 19234
rect 47182 19182 47234 19234
rect 50766 19182 50818 19234
rect 50990 19182 51042 19234
rect 15150 19070 15202 19122
rect 27134 19070 27186 19122
rect 35422 19070 35474 19122
rect 39342 19070 39394 19122
rect 45950 19070 46002 19122
rect 50542 19070 50594 19122
rect 51886 19070 51938 19122
rect 18398 18958 18450 19010
rect 18510 18958 18562 19010
rect 23998 18958 24050 19010
rect 26686 18958 26738 19010
rect 29934 18958 29986 19010
rect 30158 18958 30210 19010
rect 30382 18958 30434 19010
rect 30942 18958 30994 19010
rect 34638 18958 34690 19010
rect 34974 18958 35026 19010
rect 35982 18958 36034 19010
rect 37102 18958 37154 19010
rect 37886 18958 37938 19010
rect 38110 18958 38162 19010
rect 38334 18958 38386 19010
rect 38894 18958 38946 19010
rect 41806 18958 41858 19010
rect 42030 18958 42082 19010
rect 45278 18958 45330 19010
rect 45838 18958 45890 19010
rect 50766 18958 50818 19010
rect 51438 18958 51490 19010
rect 51550 18958 51602 19010
rect 51662 18958 51714 19010
rect 52782 18958 52834 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 21758 18622 21810 18674
rect 28478 18622 28530 18674
rect 33854 18622 33906 18674
rect 39566 18622 39618 18674
rect 39678 18622 39730 18674
rect 41246 18622 41298 18674
rect 51326 18622 51378 18674
rect 18510 18510 18562 18562
rect 24446 18510 24498 18562
rect 26014 18510 26066 18562
rect 28702 18510 28754 18562
rect 39790 18510 39842 18562
rect 45838 18510 45890 18562
rect 50878 18510 50930 18562
rect 52670 18510 52722 18562
rect 17950 18398 18002 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 19070 18398 19122 18450
rect 21982 18398 22034 18450
rect 22318 18398 22370 18450
rect 22990 18398 23042 18450
rect 23214 18398 23266 18450
rect 24222 18398 24274 18450
rect 25342 18398 25394 18450
rect 28590 18398 28642 18450
rect 29038 18398 29090 18450
rect 33630 18398 33682 18450
rect 34190 18398 34242 18450
rect 34750 18398 34802 18450
rect 35310 18398 35362 18450
rect 35982 18398 36034 18450
rect 40238 18398 40290 18450
rect 41358 18398 41410 18450
rect 41470 18398 41522 18450
rect 41806 18398 41858 18450
rect 42030 18398 42082 18450
rect 42366 18398 42418 18450
rect 42590 18398 42642 18450
rect 43150 18398 43202 18450
rect 43934 18398 43986 18450
rect 44494 18398 44546 18450
rect 45054 18398 45106 18450
rect 50430 18398 50482 18450
rect 51326 18398 51378 18450
rect 52222 18398 52274 18450
rect 52894 18398 52946 18450
rect 53118 18398 53170 18450
rect 53790 18398 53842 18450
rect 21870 18286 21922 18338
rect 22318 18286 22370 18338
rect 22766 18286 22818 18338
rect 23774 18286 23826 18338
rect 28142 18286 28194 18338
rect 31390 18286 31442 18338
rect 38110 18286 38162 18338
rect 38558 18286 38610 18338
rect 42254 18286 42306 18338
rect 43598 18286 43650 18338
rect 47966 18286 48018 18338
rect 53230 18286 53282 18338
rect 53566 18286 53618 18338
rect 54462 18286 54514 18338
rect 55134 18286 55186 18338
rect 52334 18174 52386 18226
rect 54126 18174 54178 18226
rect 54574 18174 54626 18226
rect 55246 18174 55298 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 51550 17838 51602 17890
rect 51886 17838 51938 17890
rect 52782 17838 52834 17890
rect 22318 17726 22370 17778
rect 40686 17726 40738 17778
rect 42142 17726 42194 17778
rect 44270 17726 44322 17778
rect 47070 17726 47122 17778
rect 54350 17726 54402 17778
rect 56478 17726 56530 17778
rect 17390 17614 17442 17666
rect 17950 17614 18002 17666
rect 18398 17614 18450 17666
rect 18958 17614 19010 17666
rect 19182 17614 19234 17666
rect 19854 17614 19906 17666
rect 21198 17614 21250 17666
rect 21646 17614 21698 17666
rect 21870 17614 21922 17666
rect 23102 17614 23154 17666
rect 30494 17614 30546 17666
rect 30942 17614 30994 17666
rect 31166 17614 31218 17666
rect 31502 17614 31554 17666
rect 31614 17614 31666 17666
rect 32174 17614 32226 17666
rect 35086 17614 35138 17666
rect 35534 17614 35586 17666
rect 37774 17614 37826 17666
rect 38558 17614 38610 17666
rect 41470 17614 41522 17666
rect 44942 17614 44994 17666
rect 46958 17614 47010 17666
rect 47182 17614 47234 17666
rect 50318 17614 50370 17666
rect 50654 17614 50706 17666
rect 50990 17614 51042 17666
rect 52670 17614 52722 17666
rect 57150 17614 57202 17666
rect 51326 17558 51378 17610
rect 53342 17558 53394 17610
rect 17726 17502 17778 17554
rect 22766 17502 22818 17554
rect 53566 17502 53618 17554
rect 57822 17502 57874 17554
rect 58158 17502 58210 17554
rect 17502 17390 17554 17442
rect 18286 17390 18338 17442
rect 18510 17390 18562 17442
rect 19294 17390 19346 17442
rect 19406 17390 19458 17442
rect 21422 17390 21474 17442
rect 28366 17390 28418 17442
rect 30718 17390 30770 17442
rect 31726 17390 31778 17442
rect 35982 17390 36034 17442
rect 46622 17390 46674 17442
rect 47406 17390 47458 17442
rect 50654 17390 50706 17442
rect 53118 17390 53170 17442
rect 53454 17390 53506 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 18286 17054 18338 17106
rect 27582 17054 27634 17106
rect 28030 17054 28082 17106
rect 33182 17054 33234 17106
rect 51214 17054 51266 17106
rect 51662 17054 51714 17106
rect 51886 17054 51938 17106
rect 52110 17054 52162 17106
rect 57486 17054 57538 17106
rect 58270 17054 58322 17106
rect 14702 16942 14754 16994
rect 18622 16942 18674 16994
rect 18846 16942 18898 16994
rect 19070 16942 19122 16994
rect 20638 16942 20690 16994
rect 28142 16942 28194 16994
rect 28702 16942 28754 16994
rect 30382 16942 30434 16994
rect 48974 16942 49026 16994
rect 14030 16830 14082 16882
rect 17614 16830 17666 16882
rect 18398 16830 18450 16882
rect 19630 16830 19682 16882
rect 19854 16830 19906 16882
rect 27694 16830 27746 16882
rect 28254 16830 28306 16882
rect 28926 16830 28978 16882
rect 29374 16830 29426 16882
rect 29710 16830 29762 16882
rect 49310 16830 49362 16882
rect 52670 16830 52722 16882
rect 52894 16830 52946 16882
rect 53566 16830 53618 16882
rect 16830 16718 16882 16770
rect 22766 16718 22818 16770
rect 28814 16718 28866 16770
rect 32510 16718 32562 16770
rect 33630 16718 33682 16770
rect 41022 16718 41074 16770
rect 41470 16718 41522 16770
rect 51998 16718 52050 16770
rect 53342 16718 53394 16770
rect 53790 16718 53842 16770
rect 54014 16718 54066 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 36094 16270 36146 16322
rect 36430 16270 36482 16322
rect 37774 16270 37826 16322
rect 38334 16270 38386 16322
rect 16606 16158 16658 16210
rect 18734 16158 18786 16210
rect 19742 16158 19794 16210
rect 22430 16158 22482 16210
rect 32174 16158 32226 16210
rect 35646 16158 35698 16210
rect 36094 16158 36146 16210
rect 38334 16158 38386 16210
rect 41470 16158 41522 16210
rect 49310 16158 49362 16210
rect 54910 16158 54962 16210
rect 55246 16158 55298 16210
rect 57374 16158 57426 16210
rect 15822 16046 15874 16098
rect 22766 16046 22818 16098
rect 22990 16046 23042 16098
rect 27694 16046 27746 16098
rect 29262 16046 29314 16098
rect 32510 16046 32562 16098
rect 32734 16046 32786 16098
rect 33630 16046 33682 16098
rect 33966 16046 34018 16098
rect 49534 16046 49586 16098
rect 51662 16046 51714 16098
rect 58046 16046 58098 16098
rect 19294 15934 19346 15986
rect 23326 15934 23378 15986
rect 24446 15934 24498 15986
rect 27470 15934 27522 15986
rect 28142 15934 28194 15986
rect 28366 15934 28418 15986
rect 29374 15934 29426 15986
rect 29710 15934 29762 15986
rect 34302 15934 34354 15986
rect 35310 15934 35362 15986
rect 35534 15934 35586 15986
rect 47854 15934 47906 15986
rect 50542 15934 50594 15986
rect 22990 15822 23042 15874
rect 24558 15822 24610 15874
rect 24670 15822 24722 15874
rect 25230 15822 25282 15874
rect 27918 15822 27970 15874
rect 29486 15822 29538 15874
rect 33182 15822 33234 15874
rect 33966 15822 34018 15874
rect 37998 15822 38050 15874
rect 45390 15822 45442 15874
rect 45726 15822 45778 15874
rect 52110 15822 52162 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 21870 15486 21922 15538
rect 38222 15486 38274 15538
rect 47742 15486 47794 15538
rect 52110 15486 52162 15538
rect 52334 15486 52386 15538
rect 24222 15374 24274 15426
rect 27358 15374 27410 15426
rect 34638 15374 34690 15426
rect 35758 15374 35810 15426
rect 39230 15374 39282 15426
rect 45054 15374 45106 15426
rect 49086 15374 49138 15426
rect 49422 15374 49474 15426
rect 23774 15262 23826 15314
rect 26686 15262 26738 15314
rect 31502 15262 31554 15314
rect 34078 15262 34130 15314
rect 35086 15262 35138 15314
rect 38558 15262 38610 15314
rect 39678 15262 39730 15314
rect 40238 15262 40290 15314
rect 40910 15262 40962 15314
rect 41134 15262 41186 15314
rect 41918 15262 41970 15314
rect 45278 15262 45330 15314
rect 45614 15262 45666 15314
rect 46846 15262 46898 15314
rect 47294 15262 47346 15314
rect 48974 15262 49026 15314
rect 49982 15262 50034 15314
rect 50318 15262 50370 15314
rect 50654 15262 50706 15314
rect 51662 15262 51714 15314
rect 52558 15262 52610 15314
rect 22430 15150 22482 15202
rect 23662 15150 23714 15202
rect 29486 15150 29538 15202
rect 29934 15150 29986 15202
rect 31726 15150 31778 15202
rect 33966 15150 34018 15202
rect 37886 15150 37938 15202
rect 38782 15150 38834 15202
rect 39790 15150 39842 15202
rect 42590 15150 42642 15202
rect 44718 15150 44770 15202
rect 45166 15150 45218 15202
rect 46622 15150 46674 15202
rect 47070 15150 47122 15202
rect 49310 15150 49362 15202
rect 50206 15150 50258 15202
rect 51438 15150 51490 15202
rect 52446 15150 52498 15202
rect 54126 15150 54178 15202
rect 22206 15038 22258 15090
rect 32062 15038 32114 15090
rect 41470 15038 41522 15090
rect 51102 15038 51154 15090
rect 54238 15038 54290 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 50542 14702 50594 14754
rect 52670 14702 52722 14754
rect 18286 14590 18338 14642
rect 22654 14590 22706 14642
rect 24334 14590 24386 14642
rect 26462 14590 26514 14642
rect 27582 14590 27634 14642
rect 38334 14590 38386 14642
rect 41470 14590 41522 14642
rect 43710 14590 43762 14642
rect 47854 14590 47906 14642
rect 50766 14590 50818 14642
rect 52782 14590 52834 14642
rect 53678 14590 53730 14642
rect 54350 14590 54402 14642
rect 56478 14590 56530 14642
rect 57710 14590 57762 14642
rect 18510 14478 18562 14530
rect 23550 14478 23602 14530
rect 26798 14478 26850 14530
rect 37550 14478 37602 14530
rect 39790 14478 39842 14530
rect 41694 14478 41746 14530
rect 41918 14478 41970 14530
rect 42590 14478 42642 14530
rect 42814 14478 42866 14530
rect 45054 14478 45106 14530
rect 46734 14478 46786 14530
rect 46846 14478 46898 14530
rect 48078 14478 48130 14530
rect 50206 14478 50258 14530
rect 51102 14478 51154 14530
rect 51214 14478 51266 14530
rect 52110 14478 52162 14530
rect 53566 14478 53618 14530
rect 57262 14478 57314 14530
rect 39118 14366 39170 14418
rect 39566 14366 39618 14418
rect 40910 14366 40962 14418
rect 43038 14366 43090 14418
rect 44718 14366 44770 14418
rect 47182 14366 47234 14418
rect 51774 14366 51826 14418
rect 53342 14366 53394 14418
rect 18846 14254 18898 14306
rect 22094 14254 22146 14306
rect 23214 14254 23266 14306
rect 27134 14254 27186 14306
rect 33742 14254 33794 14306
rect 37214 14254 37266 14306
rect 37886 14254 37938 14306
rect 39006 14254 39058 14306
rect 42702 14254 42754 14306
rect 44942 14254 44994 14306
rect 47070 14254 47122 14306
rect 47518 14254 47570 14306
rect 51550 14254 51602 14306
rect 51886 14254 51938 14306
rect 53118 14254 53170 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 20750 13918 20802 13970
rect 23886 13918 23938 13970
rect 24334 13918 24386 13970
rect 34190 13918 34242 13970
rect 40014 13918 40066 13970
rect 42478 13918 42530 13970
rect 43262 13918 43314 13970
rect 44158 13918 44210 13970
rect 47630 13918 47682 13970
rect 47854 13918 47906 13970
rect 50654 13918 50706 13970
rect 50766 13918 50818 13970
rect 56702 13918 56754 13970
rect 14702 13806 14754 13858
rect 18734 13806 18786 13858
rect 22654 13806 22706 13858
rect 27918 13806 27970 13858
rect 34302 13806 34354 13858
rect 35310 13806 35362 13858
rect 35758 13806 35810 13858
rect 37550 13806 37602 13858
rect 38446 13806 38498 13858
rect 41470 13806 41522 13858
rect 42814 13806 42866 13858
rect 44046 13806 44098 13858
rect 44942 13806 44994 13858
rect 45166 13806 45218 13858
rect 47406 13806 47458 13858
rect 14030 13694 14082 13746
rect 18286 13694 18338 13746
rect 18846 13694 18898 13746
rect 18958 13694 19010 13746
rect 19854 13694 19906 13746
rect 20190 13694 20242 13746
rect 20862 13694 20914 13746
rect 21086 13694 21138 13746
rect 21310 13694 21362 13746
rect 21422 13694 21474 13746
rect 21758 13694 21810 13746
rect 22430 13694 22482 13746
rect 22766 13694 22818 13746
rect 22990 13694 23042 13746
rect 23326 13694 23378 13746
rect 23662 13694 23714 13746
rect 27134 13694 27186 13746
rect 33070 13694 33122 13746
rect 33854 13694 33906 13746
rect 34526 13694 34578 13746
rect 34750 13694 34802 13746
rect 35086 13694 35138 13746
rect 39342 13694 39394 13746
rect 39566 13694 39618 13746
rect 41694 13694 41746 13746
rect 41918 13694 41970 13746
rect 42366 13694 42418 13746
rect 42702 13694 42754 13746
rect 44382 13694 44434 13746
rect 50206 13694 50258 13746
rect 50878 13694 50930 13746
rect 52670 13694 52722 13746
rect 56030 13694 56082 13746
rect 16830 13582 16882 13634
rect 17502 13582 17554 13634
rect 19406 13582 19458 13634
rect 22206 13582 22258 13634
rect 23774 13582 23826 13634
rect 30046 13582 30098 13634
rect 30494 13582 30546 13634
rect 32062 13582 32114 13634
rect 32398 13582 32450 13634
rect 38110 13582 38162 13634
rect 42142 13582 42194 13634
rect 43710 13582 43762 13634
rect 44942 13582 44994 13634
rect 47742 13582 47794 13634
rect 52782 13582 52834 13634
rect 53118 13582 53170 13634
rect 55246 13582 55298 13634
rect 20414 13470 20466 13522
rect 21982 13470 22034 13522
rect 22206 13470 22258 13522
rect 32510 13470 32562 13522
rect 33070 13470 33122 13522
rect 33406 13470 33458 13522
rect 34974 13470 35026 13522
rect 37662 13470 37714 13522
rect 38110 13470 38162 13522
rect 39006 13470 39058 13522
rect 39118 13470 39170 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17838 13134 17890 13186
rect 19966 13134 20018 13186
rect 20526 13134 20578 13186
rect 21310 13134 21362 13186
rect 23550 13134 23602 13186
rect 23774 13134 23826 13186
rect 34638 13134 34690 13186
rect 34750 13134 34802 13186
rect 44830 13134 44882 13186
rect 44942 13134 44994 13186
rect 48190 13134 48242 13186
rect 19518 13022 19570 13074
rect 20414 13022 20466 13074
rect 21422 13022 21474 13074
rect 32398 13022 32450 13074
rect 33630 13022 33682 13074
rect 34974 13022 35026 13074
rect 36430 13022 36482 13074
rect 37102 13022 37154 13074
rect 41022 13022 41074 13074
rect 42814 13022 42866 13074
rect 43374 13022 43426 13074
rect 48078 13022 48130 13074
rect 18398 12910 18450 12962
rect 18622 12910 18674 12962
rect 19854 12910 19906 12962
rect 21646 12910 21698 12962
rect 22542 12910 22594 12962
rect 23326 12910 23378 12962
rect 24222 12910 24274 12962
rect 24446 12910 24498 12962
rect 24782 12910 24834 12962
rect 25230 12910 25282 12962
rect 29486 12910 29538 12962
rect 33294 12910 33346 12962
rect 33518 12910 33570 12962
rect 35646 12910 35698 12962
rect 38782 12910 38834 12962
rect 39678 12910 39730 12962
rect 42366 12910 42418 12962
rect 43710 12910 43762 12962
rect 45838 12910 45890 12962
rect 47182 12910 47234 12962
rect 52894 12910 52946 12962
rect 17950 12798 18002 12850
rect 18734 12798 18786 12850
rect 18846 12798 18898 12850
rect 19182 12798 19234 12850
rect 22094 12798 22146 12850
rect 22430 12798 22482 12850
rect 22766 12798 22818 12850
rect 22990 12798 23042 12850
rect 30270 12798 30322 12850
rect 35422 12798 35474 12850
rect 35982 12798 36034 12850
rect 42030 12798 42082 12850
rect 44046 12798 44098 12850
rect 45278 12798 45330 12850
rect 45502 12798 45554 12850
rect 47518 12798 47570 12850
rect 47854 12798 47906 12850
rect 17838 12686 17890 12738
rect 19406 12686 19458 12738
rect 19966 12686 20018 12738
rect 23438 12686 23490 12738
rect 24334 12686 24386 12738
rect 27470 12686 27522 12738
rect 33966 12686 34018 12738
rect 34638 12686 34690 12738
rect 35646 12686 35698 12738
rect 45614 12686 45666 12738
rect 47406 12686 47458 12738
rect 51102 12686 51154 12738
rect 51438 12686 51490 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 20862 12350 20914 12402
rect 23326 12350 23378 12402
rect 24222 12350 24274 12402
rect 27022 12350 27074 12402
rect 33070 12350 33122 12402
rect 33518 12350 33570 12402
rect 34526 12350 34578 12402
rect 39006 12350 39058 12402
rect 39902 12350 39954 12402
rect 41134 12350 41186 12402
rect 42590 12350 42642 12402
rect 49758 12350 49810 12402
rect 50654 12350 50706 12402
rect 51662 12350 51714 12402
rect 52110 12350 52162 12402
rect 24558 12238 24610 12290
rect 26686 12238 26738 12290
rect 27694 12238 27746 12290
rect 35982 12238 36034 12290
rect 40910 12238 40962 12290
rect 44718 12238 44770 12290
rect 47742 12238 47794 12290
rect 50990 12238 51042 12290
rect 52222 12238 52274 12290
rect 52670 12238 52722 12290
rect 18286 12126 18338 12178
rect 27022 12126 27074 12178
rect 27246 12126 27298 12178
rect 27470 12126 27522 12178
rect 27806 12126 27858 12178
rect 30158 12126 30210 12178
rect 33294 12126 33346 12178
rect 34302 12126 34354 12178
rect 34638 12126 34690 12178
rect 34750 12126 34802 12178
rect 35310 12126 35362 12178
rect 38782 12126 38834 12178
rect 39118 12126 39170 12178
rect 39230 12126 39282 12178
rect 39566 12126 39618 12178
rect 39902 12126 39954 12178
rect 40238 12126 40290 12178
rect 50318 12126 50370 12178
rect 51326 12126 51378 12178
rect 51886 12126 51938 12178
rect 53230 12126 53282 12178
rect 18846 12014 18898 12066
rect 21198 12014 21250 12066
rect 28254 12014 28306 12066
rect 30942 12014 30994 12066
rect 33182 12014 33234 12066
rect 38110 12014 38162 12066
rect 41246 12014 41298 12066
rect 41694 12014 41746 12066
rect 42142 12014 42194 12066
rect 55358 12014 55410 12066
rect 44606 11902 44658 11954
rect 47854 11902 47906 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19518 11566 19570 11618
rect 19630 11566 19682 11618
rect 32734 11566 32786 11618
rect 33182 11566 33234 11618
rect 57262 11566 57314 11618
rect 17278 11454 17330 11506
rect 24670 11454 24722 11506
rect 26798 11454 26850 11506
rect 29262 11454 29314 11506
rect 29710 11454 29762 11506
rect 31838 11454 31890 11506
rect 33070 11454 33122 11506
rect 33518 11454 33570 11506
rect 35086 11454 35138 11506
rect 37886 11454 37938 11506
rect 38334 11454 38386 11506
rect 40238 11454 40290 11506
rect 42366 11454 42418 11506
rect 43038 11454 43090 11506
rect 46734 11454 46786 11506
rect 48862 11454 48914 11506
rect 50094 11454 50146 11506
rect 50654 11454 50706 11506
rect 52670 11454 52722 11506
rect 56030 11454 56082 11506
rect 14366 11342 14418 11394
rect 21534 11342 21586 11394
rect 24334 11342 24386 11394
rect 27470 11342 27522 11394
rect 28254 11342 28306 11394
rect 31614 11342 31666 11394
rect 32062 11342 32114 11394
rect 32286 11342 32338 11394
rect 32622 11342 32674 11394
rect 38670 11342 38722 11394
rect 39454 11342 39506 11394
rect 49646 11342 49698 11394
rect 50990 11342 51042 11394
rect 51886 11342 51938 11394
rect 52110 11342 52162 11394
rect 55582 11342 55634 11394
rect 15150 11230 15202 11282
rect 18734 11230 18786 11282
rect 18958 11230 19010 11282
rect 21310 11230 21362 11282
rect 33966 11230 34018 11282
rect 51326 11230 51378 11282
rect 51550 11230 51602 11282
rect 54798 11230 54850 11282
rect 57374 11230 57426 11282
rect 57822 11230 57874 11282
rect 58158 11230 58210 11282
rect 17726 11118 17778 11170
rect 18846 11118 18898 11170
rect 19182 11118 19234 11170
rect 20190 11118 20242 11170
rect 23998 11118 24050 11170
rect 27918 11118 27970 11170
rect 30606 11118 30658 11170
rect 31502 11118 31554 11170
rect 39006 11118 39058 11170
rect 51102 11118 51154 11170
rect 51774 11118 51826 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 15822 10782 15874 10834
rect 18174 10782 18226 10834
rect 26686 10782 26738 10834
rect 27246 10782 27298 10834
rect 31166 10782 31218 10834
rect 31726 10782 31778 10834
rect 41694 10782 41746 10834
rect 42814 10782 42866 10834
rect 47182 10782 47234 10834
rect 51998 10782 52050 10834
rect 15934 10670 15986 10722
rect 18062 10670 18114 10722
rect 18398 10670 18450 10722
rect 18734 10670 18786 10722
rect 23774 10670 23826 10722
rect 27022 10670 27074 10722
rect 43934 10670 43986 10722
rect 50206 10670 50258 10722
rect 51326 10670 51378 10722
rect 51438 10670 51490 10722
rect 17838 10558 17890 10610
rect 24558 10558 24610 10610
rect 25342 10558 25394 10610
rect 26910 10558 26962 10610
rect 30270 10558 30322 10610
rect 30942 10558 30994 10610
rect 31278 10558 31330 10610
rect 42254 10558 42306 10610
rect 43150 10558 43202 10610
rect 46846 10558 46898 10610
rect 49870 10558 49922 10610
rect 51662 10558 51714 10610
rect 58158 10558 58210 10610
rect 21646 10446 21698 10498
rect 27470 10446 27522 10498
rect 29598 10446 29650 10498
rect 46062 10446 46114 10498
rect 49534 10446 49586 10498
rect 50654 10446 50706 10498
rect 18958 10334 19010 10386
rect 19182 10334 19234 10386
rect 19406 10334 19458 10386
rect 19854 10334 19906 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 17950 9998 18002 10050
rect 15934 9886 15986 9938
rect 17614 9886 17666 9938
rect 18622 9886 18674 9938
rect 19966 9886 20018 9938
rect 22206 9886 22258 9938
rect 26686 9886 26738 9938
rect 30494 9886 30546 9938
rect 32286 9886 32338 9938
rect 35422 9886 35474 9938
rect 42590 9886 42642 9938
rect 43486 9886 43538 9938
rect 52110 9886 52162 9938
rect 18174 9774 18226 9826
rect 18846 9774 18898 9826
rect 19406 9774 19458 9826
rect 19518 9774 19570 9826
rect 21758 9774 21810 9826
rect 24894 9774 24946 9826
rect 25342 9774 25394 9826
rect 27582 9774 27634 9826
rect 28030 9774 28082 9826
rect 31166 9774 31218 9826
rect 31838 9774 31890 9826
rect 32958 9774 33010 9826
rect 33294 9774 33346 9826
rect 33518 9774 33570 9826
rect 33854 9774 33906 9826
rect 35646 9774 35698 9826
rect 35870 9774 35922 9826
rect 36094 9774 36146 9826
rect 37662 9774 37714 9826
rect 41470 9774 41522 9826
rect 42926 9774 42978 9826
rect 43822 9774 43874 9826
rect 50766 9774 50818 9826
rect 52558 9774 52610 9826
rect 52894 9774 52946 9826
rect 53230 9774 53282 9826
rect 18622 9662 18674 9714
rect 23438 9662 23490 9714
rect 26462 9662 26514 9714
rect 28590 9662 28642 9714
rect 29934 9662 29986 9714
rect 30718 9662 30770 9714
rect 31502 9662 31554 9714
rect 32846 9662 32898 9714
rect 34190 9662 34242 9714
rect 34526 9662 34578 9714
rect 36542 9662 36594 9714
rect 37774 9662 37826 9714
rect 39566 9662 39618 9714
rect 40350 9662 40402 9714
rect 50878 9662 50930 9714
rect 51102 9662 51154 9714
rect 51438 9662 51490 9714
rect 15822 9550 15874 9602
rect 19070 9550 19122 9602
rect 21422 9550 21474 9602
rect 27582 9550 27634 9602
rect 30046 9550 30098 9602
rect 30382 9550 30434 9602
rect 30606 9550 30658 9602
rect 32622 9550 32674 9602
rect 33518 9550 33570 9602
rect 44158 9550 44210 9602
rect 50430 9550 50482 9602
rect 52894 9550 52946 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 17502 9214 17554 9266
rect 18734 9214 18786 9266
rect 18846 9214 18898 9266
rect 22094 9214 22146 9266
rect 31390 9214 31442 9266
rect 33294 9214 33346 9266
rect 33854 9214 33906 9266
rect 39230 9214 39282 9266
rect 40238 9214 40290 9266
rect 41918 9214 41970 9266
rect 42478 9214 42530 9266
rect 42814 9214 42866 9266
rect 43486 9214 43538 9266
rect 44382 9214 44434 9266
rect 50206 9214 50258 9266
rect 55694 9214 55746 9266
rect 14702 9102 14754 9154
rect 18958 9102 19010 9154
rect 31054 9102 31106 9154
rect 33518 9102 33570 9154
rect 33630 9102 33682 9154
rect 35534 9102 35586 9154
rect 37102 9102 37154 9154
rect 37326 9102 37378 9154
rect 37662 9102 37714 9154
rect 39566 9102 39618 9154
rect 39902 9102 39954 9154
rect 42142 9102 42194 9154
rect 43150 9102 43202 9154
rect 43822 9102 43874 9154
rect 54462 9102 54514 9154
rect 14030 8990 14082 9042
rect 19294 8990 19346 9042
rect 22430 8990 22482 9042
rect 35086 8990 35138 9042
rect 35310 8990 35362 9042
rect 44718 8990 44770 9042
rect 49758 8990 49810 9042
rect 50430 8990 50482 9042
rect 55246 8990 55298 9042
rect 16830 8878 16882 8930
rect 35422 8878 35474 8930
rect 37550 8878 37602 8930
rect 45502 8878 45554 8930
rect 47630 8878 47682 8930
rect 50318 8878 50370 8930
rect 52334 8878 52386 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 35310 8430 35362 8482
rect 33630 8318 33682 8370
rect 47518 8318 47570 8370
rect 50206 8318 50258 8370
rect 51102 8318 51154 8370
rect 26910 8206 26962 8258
rect 27358 8206 27410 8258
rect 30942 8206 30994 8258
rect 31502 8206 31554 8258
rect 32174 8206 32226 8258
rect 33966 8206 34018 8258
rect 35534 8206 35586 8258
rect 35870 8206 35922 8258
rect 44942 8206 44994 8258
rect 45166 8206 45218 8258
rect 45614 8206 45666 8258
rect 45838 8206 45890 8258
rect 46286 8206 46338 8258
rect 46398 8206 46450 8258
rect 47294 8206 47346 8258
rect 47630 8206 47682 8258
rect 48526 8206 48578 8258
rect 48750 8206 48802 8258
rect 48974 8206 49026 8258
rect 49646 8206 49698 8258
rect 50766 8206 50818 8258
rect 51326 8206 51378 8258
rect 30606 8094 30658 8146
rect 31166 8094 31218 8146
rect 36318 8094 36370 8146
rect 39006 8094 39058 8146
rect 39678 8094 39730 8146
rect 47966 8094 48018 8146
rect 48302 8094 48354 8146
rect 49982 8094 50034 8146
rect 26686 7982 26738 8034
rect 26798 7982 26850 8034
rect 30718 7982 30770 8034
rect 31614 7982 31666 8034
rect 31726 7982 31778 8034
rect 32510 7982 32562 8034
rect 33742 7982 33794 8034
rect 34974 7982 35026 8034
rect 35982 7982 36034 8034
rect 36094 7982 36146 8034
rect 39342 7982 39394 8034
rect 45502 7982 45554 8034
rect 46174 7982 46226 8034
rect 46622 7982 46674 8034
rect 49422 7982 49474 8034
rect 51662 7982 51714 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 19070 7646 19122 7698
rect 24782 7646 24834 7698
rect 31502 7646 31554 7698
rect 38446 7646 38498 7698
rect 38894 7646 38946 7698
rect 40014 7646 40066 7698
rect 41246 7646 41298 7698
rect 41470 7646 41522 7698
rect 43598 7646 43650 7698
rect 45838 7646 45890 7698
rect 50094 7646 50146 7698
rect 18734 7534 18786 7586
rect 19294 7534 19346 7586
rect 26798 7534 26850 7586
rect 29822 7534 29874 7586
rect 33966 7534 34018 7586
rect 35646 7534 35698 7586
rect 36430 7534 36482 7586
rect 39790 7534 39842 7586
rect 40126 7534 40178 7586
rect 43262 7534 43314 7586
rect 50878 7534 50930 7586
rect 51214 7534 51266 7586
rect 18958 7422 19010 7474
rect 19630 7422 19682 7474
rect 23326 7422 23378 7474
rect 24334 7422 24386 7474
rect 26350 7422 26402 7474
rect 26574 7422 26626 7474
rect 27022 7422 27074 7474
rect 27246 7422 27298 7474
rect 30494 7422 30546 7474
rect 33630 7422 33682 7474
rect 33742 7422 33794 7474
rect 34302 7422 34354 7474
rect 34414 7422 34466 7474
rect 34638 7422 34690 7474
rect 35086 7422 35138 7474
rect 35310 7422 35362 7474
rect 35422 7422 35474 7474
rect 36094 7422 36146 7474
rect 36766 7422 36818 7474
rect 37886 7422 37938 7474
rect 38110 7422 38162 7474
rect 38670 7422 38722 7474
rect 40350 7422 40402 7474
rect 40798 7422 40850 7474
rect 42926 7422 42978 7474
rect 43822 7422 43874 7474
rect 44158 7422 44210 7474
rect 49646 7422 49698 7474
rect 49870 7422 49922 7474
rect 50542 7422 50594 7474
rect 50654 7422 50706 7474
rect 51438 7422 51490 7474
rect 20190 7310 20242 7362
rect 21086 7310 21138 7362
rect 21310 7310 21362 7362
rect 23662 7310 23714 7362
rect 25790 7310 25842 7362
rect 27694 7310 27746 7362
rect 31838 7310 31890 7362
rect 38558 7310 38610 7362
rect 41358 7310 41410 7362
rect 42590 7310 42642 7362
rect 43710 7310 43762 7362
rect 44158 7310 44210 7362
rect 19966 7198 20018 7250
rect 20750 7198 20802 7250
rect 22766 7198 22818 7250
rect 23102 7198 23154 7250
rect 23886 7198 23938 7250
rect 24110 7198 24162 7250
rect 26126 7198 26178 7250
rect 35982 7198 36034 7250
rect 37550 7198 37602 7250
rect 44606 7310 44658 7362
rect 49758 7310 49810 7362
rect 51550 7310 51602 7362
rect 52446 7310 52498 7362
rect 44606 7198 44658 7250
rect 52558 7198 52610 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19518 6862 19570 6914
rect 21422 6862 21474 6914
rect 23550 6862 23602 6914
rect 26798 6862 26850 6914
rect 26910 6862 26962 6914
rect 32286 6862 32338 6914
rect 38782 6862 38834 6914
rect 38894 6862 38946 6914
rect 40798 6862 40850 6914
rect 40910 6862 40962 6914
rect 41582 6862 41634 6914
rect 50318 6862 50370 6914
rect 18286 6750 18338 6802
rect 18622 6750 18674 6802
rect 22206 6750 22258 6802
rect 24334 6750 24386 6802
rect 31950 6750 32002 6802
rect 32286 6750 32338 6802
rect 36206 6750 36258 6802
rect 46398 6750 46450 6802
rect 48750 6750 48802 6802
rect 49758 6750 49810 6802
rect 50430 6750 50482 6802
rect 52670 6750 52722 6802
rect 15486 6638 15538 6690
rect 18734 6638 18786 6690
rect 19630 6638 19682 6690
rect 20526 6638 20578 6690
rect 20638 6638 20690 6690
rect 21310 6638 21362 6690
rect 22318 6638 22370 6690
rect 23438 6638 23490 6690
rect 24446 6638 24498 6690
rect 25454 6638 25506 6690
rect 25902 6638 25954 6690
rect 27582 6638 27634 6690
rect 28030 6638 28082 6690
rect 30942 6638 30994 6690
rect 31278 6638 31330 6690
rect 31950 6638 32002 6690
rect 37886 6638 37938 6690
rect 38222 6638 38274 6690
rect 41246 6638 41298 6690
rect 41806 6638 41858 6690
rect 43486 6638 43538 6690
rect 43934 6638 43986 6690
rect 46846 6638 46898 6690
rect 48414 6638 48466 6690
rect 49982 6638 50034 6690
rect 50990 6638 51042 6690
rect 54798 6638 54850 6690
rect 55470 6638 55522 6690
rect 56030 6638 56082 6690
rect 16158 6526 16210 6578
rect 18958 6526 19010 6578
rect 19294 6526 19346 6578
rect 21982 6526 22034 6578
rect 24110 6526 24162 6578
rect 24782 6526 24834 6578
rect 25006 6526 25058 6578
rect 26238 6526 26290 6578
rect 27246 6526 27298 6578
rect 31502 6526 31554 6578
rect 38558 6526 38610 6578
rect 40014 6526 40066 6578
rect 40238 6526 40290 6578
rect 40462 6526 40514 6578
rect 42926 6526 42978 6578
rect 43262 6526 43314 6578
rect 48526 6526 48578 6578
rect 48862 6526 48914 6578
rect 49422 6526 49474 6578
rect 50766 6526 50818 6578
rect 51214 6526 51266 6578
rect 20302 6414 20354 6466
rect 20750 6414 20802 6466
rect 21758 6414 21810 6466
rect 23886 6414 23938 6466
rect 25118 6414 25170 6466
rect 26126 6414 26178 6466
rect 26462 6414 26514 6466
rect 30158 6414 30210 6466
rect 30494 6414 30546 6466
rect 30718 6414 30770 6466
rect 30830 6414 30882 6466
rect 31390 6414 31442 6466
rect 38110 6414 38162 6466
rect 40126 6414 40178 6466
rect 43150 6414 43202 6466
rect 51102 6414 51154 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 17390 6078 17442 6130
rect 18510 6078 18562 6130
rect 18846 6078 18898 6130
rect 21646 6078 21698 6130
rect 23662 6078 23714 6130
rect 23774 6078 23826 6130
rect 23998 6078 24050 6130
rect 17502 5966 17554 6018
rect 19070 5966 19122 6018
rect 21534 5966 21586 6018
rect 22094 5966 22146 6018
rect 19406 5854 19458 5906
rect 21758 5854 21810 5906
rect 23550 5854 23602 5906
rect 30382 5854 30434 5906
rect 30830 6078 30882 6130
rect 31278 6078 31330 6130
rect 32174 6078 32226 6130
rect 32510 6078 32562 6130
rect 46286 6078 46338 6130
rect 31614 5966 31666 6018
rect 33854 5966 33906 6018
rect 35422 5966 35474 6018
rect 43710 5966 43762 6018
rect 46174 5966 46226 6018
rect 46510 5966 46562 6018
rect 46958 5966 47010 6018
rect 47070 5966 47122 6018
rect 47182 5966 47234 6018
rect 30942 5854 30994 5906
rect 31390 5854 31442 5906
rect 44382 5854 44434 5906
rect 45054 5854 45106 5906
rect 45278 5854 45330 5906
rect 45614 5854 45666 5906
rect 46734 5854 46786 5906
rect 18958 5742 19010 5794
rect 27582 5742 27634 5794
rect 29710 5742 29762 5794
rect 30718 5742 30770 5794
rect 41246 5742 41298 5794
rect 41582 5742 41634 5794
rect 45166 5742 45218 5794
rect 47518 5742 47570 5794
rect 33742 5630 33794 5682
rect 35534 5630 35586 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 20190 5182 20242 5234
rect 21422 5182 21474 5234
rect 23214 5182 23266 5234
rect 26126 5182 26178 5234
rect 31054 5182 31106 5234
rect 31614 5182 31666 5234
rect 32062 5182 32114 5234
rect 33518 5182 33570 5234
rect 35646 5182 35698 5234
rect 36990 5182 37042 5234
rect 40350 5182 40402 5234
rect 40686 5182 40738 5234
rect 44046 5182 44098 5234
rect 44942 5182 44994 5234
rect 47742 5182 47794 5234
rect 49870 5182 49922 5234
rect 51214 5182 51266 5234
rect 30718 5070 30770 5122
rect 30942 5070 30994 5122
rect 31166 5070 31218 5122
rect 32734 5070 32786 5122
rect 39118 5070 39170 5122
rect 39790 5070 39842 5122
rect 45502 5070 45554 5122
rect 45838 5070 45890 5122
rect 46398 5070 46450 5122
rect 47070 5070 47122 5122
rect 50318 5070 50370 5122
rect 20078 4846 20130 4898
rect 23102 4846 23154 4898
rect 26014 4846 26066 4898
rect 40798 4846 40850 4898
rect 45950 4846 46002 4898
rect 46062 4846 46114 4898
rect 51326 4846 51378 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 28590 4510 28642 4562
rect 33182 4510 33234 4562
rect 37662 4510 37714 4562
rect 38222 4510 38274 4562
rect 48750 4510 48802 4562
rect 53902 4510 53954 4562
rect 19182 4398 19234 4450
rect 22430 4398 22482 4450
rect 26014 4398 26066 4450
rect 31502 4398 31554 4450
rect 36430 4398 36482 4450
rect 38110 4398 38162 4450
rect 41694 4398 41746 4450
rect 44942 4398 44994 4450
rect 48862 4398 48914 4450
rect 52670 4398 52722 4450
rect 18510 4286 18562 4338
rect 21646 4286 21698 4338
rect 25342 4286 25394 4338
rect 32286 4286 32338 4338
rect 37214 4286 37266 4338
rect 40910 4286 40962 4338
rect 44158 4286 44210 4338
rect 53342 4286 53394 4338
rect 57598 4286 57650 4338
rect 58158 4286 58210 4338
rect 21310 4174 21362 4226
rect 24558 4174 24610 4226
rect 28142 4174 28194 4226
rect 29374 4174 29426 4226
rect 34302 4174 34354 4226
rect 43822 4174 43874 4226
rect 47070 4174 47122 4226
rect 50542 4174 50594 4226
rect 57374 4174 57426 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 21646 3614 21698 3666
rect 43934 3614 43986 3666
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2688 69200 2800 70000
rect 4704 69200 4816 70000
rect 6720 69200 6832 70000
rect 8736 69200 8848 70000
rect 10752 69200 10864 70000
rect 12768 69200 12880 70000
rect 14784 69200 14896 70000
rect 16800 69200 16912 70000
rect 18816 69200 18928 70000
rect 20832 69200 20944 70000
rect 22848 69200 22960 70000
rect 24864 69200 24976 70000
rect 26880 69200 26992 70000
rect 28896 69200 29008 70000
rect 30912 69200 31024 70000
rect 32928 69200 33040 70000
rect 34944 69200 35056 70000
rect 36960 69200 37072 70000
rect 38976 69200 39088 70000
rect 40992 69200 41104 70000
rect 43008 69200 43120 70000
rect 45024 69200 45136 70000
rect 47040 69200 47152 70000
rect 49056 69200 49168 70000
rect 51072 69200 51184 70000
rect 53088 69200 53200 70000
rect 55104 69200 55216 70000
rect 57120 69200 57232 70000
rect 2716 67228 2772 69200
rect 2716 67172 2996 67228
rect 2940 66162 2996 67172
rect 4732 66836 4788 69200
rect 6748 67228 6804 69200
rect 6748 67172 7028 67228
rect 4732 66770 4788 66780
rect 5516 66836 5572 66846
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 2940 66110 2942 66162
rect 2994 66110 2996 66162
rect 2940 66098 2996 66110
rect 5516 66162 5572 66780
rect 5516 66110 5518 66162
rect 5570 66110 5572 66162
rect 5516 66098 5572 66110
rect 6972 66162 7028 67172
rect 8764 66834 8820 69200
rect 10780 67228 10836 69200
rect 12796 67228 12852 69200
rect 14812 67228 14868 69200
rect 16828 67228 16884 69200
rect 10780 67172 11060 67228
rect 12796 67172 13188 67228
rect 14812 67172 15092 67228
rect 16828 67172 17108 67228
rect 8764 66782 8766 66834
rect 8818 66782 8820 66834
rect 8764 66770 8820 66782
rect 9324 66834 9380 66846
rect 9324 66782 9326 66834
rect 9378 66782 9380 66834
rect 6972 66110 6974 66162
rect 7026 66110 7028 66162
rect 6972 66098 7028 66110
rect 9324 66162 9380 66782
rect 9324 66110 9326 66162
rect 9378 66110 9380 66162
rect 9324 66098 9380 66110
rect 11004 66162 11060 67172
rect 11004 66110 11006 66162
rect 11058 66110 11060 66162
rect 11004 66098 11060 66110
rect 13132 66162 13188 67172
rect 13132 66110 13134 66162
rect 13186 66110 13188 66162
rect 13132 66098 13188 66110
rect 15036 66162 15092 67172
rect 15036 66110 15038 66162
rect 15090 66110 15092 66162
rect 15036 66098 15092 66110
rect 17052 66162 17108 67172
rect 18844 66386 18900 69200
rect 20860 67228 20916 69200
rect 20860 67172 21140 67228
rect 18844 66334 18846 66386
rect 18898 66334 18900 66386
rect 18844 66322 18900 66334
rect 17612 66276 17668 66286
rect 17052 66110 17054 66162
rect 17106 66110 17108 66162
rect 17052 66098 17108 66110
rect 17388 66274 17668 66276
rect 17388 66222 17614 66274
rect 17666 66222 17668 66274
rect 17388 66220 17668 66222
rect 12572 65380 12628 65390
rect 12572 65378 12740 65380
rect 12572 65326 12574 65378
rect 12626 65326 12740 65378
rect 12572 65324 12740 65326
rect 12572 65314 12628 65324
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 8540 64876 8932 64932
rect 8540 64818 8596 64876
rect 8540 64766 8542 64818
rect 8594 64766 8596 64818
rect 8540 64754 8596 64766
rect 5740 64706 5796 64718
rect 5740 64654 5742 64706
rect 5794 64654 5796 64706
rect 5740 63924 5796 64654
rect 8764 64708 8820 64718
rect 6412 64596 6468 64606
rect 6412 64594 6692 64596
rect 6412 64542 6414 64594
rect 6466 64542 6692 64594
rect 6412 64540 6692 64542
rect 6412 64530 6468 64540
rect 5740 63858 5796 63868
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 6636 63250 6692 64540
rect 8764 64146 8820 64652
rect 8876 64706 8932 64876
rect 10108 64820 10164 64830
rect 10108 64726 10164 64764
rect 12236 64818 12292 64830
rect 12236 64766 12238 64818
rect 12290 64766 12292 64818
rect 8876 64654 8878 64706
rect 8930 64654 8932 64706
rect 8876 64642 8932 64654
rect 9436 64708 9492 64718
rect 9436 64614 9492 64652
rect 11340 64596 11396 64606
rect 8764 64094 8766 64146
rect 8818 64094 8820 64146
rect 8764 63924 8820 64094
rect 6636 63198 6638 63250
rect 6690 63198 6692 63250
rect 6636 63186 6692 63198
rect 8652 63868 8764 63924
rect 6748 63138 6804 63150
rect 6748 63086 6750 63138
rect 6802 63086 6804 63138
rect 6524 63028 6580 63038
rect 6524 62934 6580 62972
rect 6748 62356 6804 63086
rect 7868 63138 7924 63150
rect 8092 63140 8148 63150
rect 7868 63086 7870 63138
rect 7922 63086 7924 63138
rect 7084 63028 7140 63038
rect 7308 63028 7364 63038
rect 7084 63026 7252 63028
rect 7084 62974 7086 63026
rect 7138 62974 7252 63026
rect 7084 62972 7252 62974
rect 7084 62962 7140 62972
rect 7196 62578 7252 62972
rect 7196 62526 7198 62578
rect 7250 62526 7252 62578
rect 7196 62514 7252 62526
rect 7308 62578 7364 62972
rect 7644 63028 7700 63038
rect 7644 62934 7700 62972
rect 7308 62526 7310 62578
rect 7362 62526 7364 62578
rect 7308 62514 7364 62526
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 6748 61684 6804 62300
rect 6860 62466 6916 62478
rect 6860 62414 6862 62466
rect 6914 62414 6916 62466
rect 6860 62188 6916 62414
rect 7868 62468 7924 63086
rect 7868 62374 7924 62412
rect 7980 63138 8148 63140
rect 7980 63086 8094 63138
rect 8146 63086 8148 63138
rect 7980 63084 8148 63086
rect 7980 62466 8036 63084
rect 8092 63074 8148 63084
rect 8540 62580 8596 62590
rect 8540 62486 8596 62524
rect 7980 62414 7982 62466
rect 8034 62414 8036 62466
rect 7084 62356 7140 62366
rect 7084 62262 7140 62300
rect 7980 62356 8036 62414
rect 7980 62290 8036 62300
rect 8204 62356 8260 62366
rect 8428 62356 8484 62366
rect 8204 62354 8484 62356
rect 8204 62302 8206 62354
rect 8258 62302 8430 62354
rect 8482 62302 8484 62354
rect 8204 62300 8484 62302
rect 8204 62290 8260 62300
rect 8428 62290 8484 62300
rect 6860 62132 7588 62188
rect 6748 61628 7028 61684
rect 6412 61460 6468 61470
rect 6748 61460 6804 61470
rect 6412 61458 6804 61460
rect 6412 61406 6414 61458
rect 6466 61406 6750 61458
rect 6802 61406 6804 61458
rect 6412 61404 6804 61406
rect 6412 61394 6468 61404
rect 6188 61348 6244 61358
rect 6188 60900 6244 61292
rect 6300 61346 6356 61358
rect 6300 61294 6302 61346
rect 6354 61294 6356 61346
rect 6300 61124 6356 61294
rect 6300 61068 6580 61124
rect 6300 60900 6356 60910
rect 6188 60898 6356 60900
rect 6188 60846 6302 60898
rect 6354 60846 6356 60898
rect 6188 60844 6356 60846
rect 2828 60786 2884 60798
rect 2828 60734 2830 60786
rect 2882 60734 2884 60786
rect 2828 60116 2884 60734
rect 1820 59106 1876 59118
rect 1820 59054 1822 59106
rect 1874 59054 1876 59106
rect 1708 58324 1764 58334
rect 1820 58324 1876 59054
rect 1764 58268 1876 58324
rect 2268 58434 2324 58446
rect 2268 58382 2270 58434
rect 2322 58382 2324 58434
rect 1708 58230 1764 58268
rect 1820 57764 1876 57774
rect 1820 57650 1876 57708
rect 1820 57598 1822 57650
rect 1874 57598 1876 57650
rect 1820 54514 1876 57598
rect 1820 54462 1822 54514
rect 1874 54462 1876 54514
rect 1820 54450 1876 54462
rect 1820 50594 1876 50606
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1820 47572 1876 50542
rect 1820 47458 1876 47516
rect 1820 47406 1822 47458
rect 1874 47406 1876 47458
rect 1820 47394 1876 47406
rect 2268 43708 2324 58382
rect 2492 58212 2548 58222
rect 2492 57762 2548 58156
rect 2492 57710 2494 57762
rect 2546 57710 2548 57762
rect 2492 57698 2548 57710
rect 2828 57764 2884 60060
rect 3500 60674 3556 60686
rect 3500 60622 3502 60674
rect 3554 60622 3556 60674
rect 3500 59444 3556 60622
rect 5628 60676 5684 60686
rect 5628 60582 5684 60620
rect 6300 60676 6356 60844
rect 6300 60610 6356 60620
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 6524 60002 6580 61068
rect 6524 59950 6526 60002
rect 6578 59950 6580 60002
rect 6524 59938 6580 59950
rect 6748 60786 6804 61404
rect 6860 61348 6916 61358
rect 6860 61254 6916 61292
rect 6748 60734 6750 60786
rect 6802 60734 6804 60786
rect 3500 59378 3556 59388
rect 5852 59780 5908 59790
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4060 58434 4116 58446
rect 4060 58382 4062 58434
rect 4114 58382 4116 58434
rect 2828 57698 2884 57708
rect 3836 58322 3892 58334
rect 3836 58270 3838 58322
rect 3890 58270 3892 58322
rect 3836 57764 3892 58270
rect 3948 58212 4004 58222
rect 3948 58118 4004 58156
rect 3836 57698 3892 57708
rect 4060 56868 4116 58382
rect 4284 58434 4340 58446
rect 4284 58382 4286 58434
rect 4338 58382 4340 58434
rect 4060 56802 4116 56812
rect 4172 57764 4228 57774
rect 4172 56756 4228 57708
rect 4284 56980 4340 58382
rect 5628 58322 5684 58334
rect 5628 58270 5630 58322
rect 5682 58270 5684 58322
rect 4844 58210 4900 58222
rect 4844 58158 4846 58210
rect 4898 58158 4900 58210
rect 4844 58100 4900 58158
rect 5516 58212 5572 58222
rect 5068 58100 5124 58110
rect 4844 58044 5068 58100
rect 4956 57764 5012 57774
rect 4956 57670 5012 57708
rect 4620 57540 4676 57550
rect 4620 57446 4676 57484
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4396 56980 4452 56990
rect 4284 56978 4452 56980
rect 4284 56926 4398 56978
rect 4450 56926 4452 56978
rect 4284 56924 4452 56926
rect 4396 56914 4452 56924
rect 4508 56868 4564 56878
rect 4508 56774 4564 56812
rect 4844 56868 4900 56878
rect 4284 56756 4340 56766
rect 4172 56754 4340 56756
rect 4172 56702 4286 56754
rect 4338 56702 4340 56754
rect 4172 56700 4340 56702
rect 4284 56690 4340 56700
rect 4508 55972 4564 55982
rect 4284 55970 4564 55972
rect 4284 55918 4510 55970
rect 4562 55918 4564 55970
rect 4284 55916 4564 55918
rect 4284 55524 4340 55916
rect 4508 55906 4564 55916
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4396 55524 4452 55534
rect 4284 55468 4396 55524
rect 3388 55300 3444 55310
rect 3836 55300 3892 55310
rect 3388 55298 3892 55300
rect 3388 55246 3390 55298
rect 3442 55246 3838 55298
rect 3890 55246 3892 55298
rect 3388 55244 3892 55246
rect 3388 55234 3444 55244
rect 3836 55234 3892 55244
rect 4396 55298 4452 55468
rect 4732 55524 4788 55534
rect 4844 55524 4900 56812
rect 4956 56866 5012 56878
rect 4956 56814 4958 56866
rect 5010 56814 5012 56866
rect 4956 55972 5012 56814
rect 5068 56756 5124 58044
rect 5516 57652 5572 58156
rect 5628 57876 5684 58270
rect 5740 58212 5796 58222
rect 5740 58118 5796 58156
rect 5852 58100 5908 59724
rect 5964 58212 6020 58222
rect 5964 58210 6356 58212
rect 5964 58158 5966 58210
rect 6018 58158 6356 58210
rect 5964 58156 6356 58158
rect 5964 58146 6020 58156
rect 5852 58034 5908 58044
rect 5628 57820 5908 57876
rect 5628 57652 5684 57662
rect 5516 57650 5684 57652
rect 5516 57598 5630 57650
rect 5682 57598 5684 57650
rect 5516 57596 5684 57598
rect 5628 57540 5684 57596
rect 5516 56868 5572 56878
rect 5628 56868 5684 57484
rect 5852 57538 5908 57820
rect 6300 57650 6356 58156
rect 6300 57598 6302 57650
rect 6354 57598 6356 57650
rect 6300 57586 6356 57598
rect 6748 57652 6804 60734
rect 6972 60226 7028 61628
rect 7084 61348 7140 61358
rect 7532 61348 7588 62132
rect 7084 61346 7476 61348
rect 7084 61294 7086 61346
rect 7138 61294 7476 61346
rect 7084 61292 7476 61294
rect 7084 61282 7140 61292
rect 6972 60174 6974 60226
rect 7026 60174 7028 60226
rect 6972 60162 7028 60174
rect 7084 60002 7140 60014
rect 7084 59950 7086 60002
rect 7138 59950 7140 60002
rect 7084 59780 7140 59950
rect 7420 60002 7476 61292
rect 7532 61346 7700 61348
rect 7532 61294 7534 61346
rect 7586 61294 7700 61346
rect 7532 61292 7700 61294
rect 7532 61282 7588 61292
rect 7420 59950 7422 60002
rect 7474 59950 7476 60002
rect 7420 59938 7476 59950
rect 7532 60786 7588 60798
rect 7532 60734 7534 60786
rect 7586 60734 7588 60786
rect 7532 59780 7588 60734
rect 6860 59724 7588 59780
rect 6860 57874 6916 59724
rect 7644 59668 7700 61292
rect 6860 57822 6862 57874
rect 6914 57822 6916 57874
rect 6860 57810 6916 57822
rect 7196 59612 7700 59668
rect 7868 61010 7924 61022
rect 7868 60958 7870 61010
rect 7922 60958 7924 61010
rect 6748 57596 6916 57652
rect 5852 57486 5854 57538
rect 5906 57486 5908 57538
rect 5852 57092 5908 57486
rect 6524 57428 6580 57438
rect 5852 57026 5908 57036
rect 6076 57426 6580 57428
rect 6076 57374 6526 57426
rect 6578 57374 6580 57426
rect 6076 57372 6580 57374
rect 6076 56978 6132 57372
rect 6524 57362 6580 57372
rect 6076 56926 6078 56978
rect 6130 56926 6132 56978
rect 6076 56914 6132 56926
rect 6188 57092 6244 57102
rect 5964 56868 6020 56878
rect 5628 56866 6020 56868
rect 5628 56814 5966 56866
rect 6018 56814 6020 56866
rect 5628 56812 6020 56814
rect 5516 56774 5572 56812
rect 5964 56802 6020 56812
rect 5292 56756 5348 56766
rect 5068 56700 5292 56756
rect 5068 55972 5124 55982
rect 4956 55970 5124 55972
rect 4956 55918 5070 55970
rect 5122 55918 5124 55970
rect 4956 55916 5124 55918
rect 5068 55636 5124 55916
rect 5068 55570 5124 55580
rect 4732 55522 4900 55524
rect 4732 55470 4734 55522
rect 4786 55470 4900 55522
rect 4732 55468 4900 55470
rect 4732 55458 4788 55468
rect 4396 55246 4398 55298
rect 4450 55246 4452 55298
rect 4396 55234 4452 55246
rect 2828 55186 2884 55198
rect 2828 55134 2830 55186
rect 2882 55134 2884 55186
rect 2828 55076 2884 55134
rect 3164 55186 3220 55198
rect 3164 55134 3166 55186
rect 3218 55134 3220 55186
rect 2828 55010 2884 55020
rect 2940 55074 2996 55086
rect 2940 55022 2942 55074
rect 2994 55022 2996 55074
rect 2940 54740 2996 55022
rect 2492 54684 2996 54740
rect 3052 55076 3108 55086
rect 2492 54626 2548 54684
rect 3052 54628 3108 55020
rect 2492 54574 2494 54626
rect 2546 54574 2548 54626
rect 2492 54562 2548 54574
rect 2940 54572 3108 54628
rect 3164 54628 3220 55134
rect 4844 55188 4900 55198
rect 4844 55186 5124 55188
rect 4844 55134 4846 55186
rect 4898 55134 5124 55186
rect 4844 55132 5124 55134
rect 4844 55122 4900 55132
rect 3724 55076 3780 55086
rect 3724 54982 3780 55020
rect 3948 55074 4004 55086
rect 3948 55022 3950 55074
rect 4002 55022 4004 55074
rect 2940 53842 2996 54572
rect 3164 54562 3220 54572
rect 3948 54628 4004 55022
rect 3948 54562 4004 54572
rect 4732 55074 4788 55086
rect 4732 55022 4734 55074
rect 4786 55022 4788 55074
rect 4620 54516 4676 54526
rect 4620 54404 4676 54460
rect 4284 54402 4676 54404
rect 4284 54350 4622 54402
rect 4674 54350 4676 54402
rect 4284 54348 4676 54350
rect 2940 53790 2942 53842
rect 2994 53790 2996 53842
rect 2940 53778 2996 53790
rect 3388 53956 3444 53966
rect 3388 53730 3444 53900
rect 4284 53956 4340 54348
rect 4620 54338 4676 54348
rect 4732 54292 4788 55022
rect 5068 54738 5124 55132
rect 5068 54686 5070 54738
rect 5122 54686 5124 54738
rect 5068 54674 5124 54686
rect 4956 54514 5012 54526
rect 4956 54462 4958 54514
rect 5010 54462 5012 54514
rect 4732 54236 4900 54292
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4844 53956 4900 54236
rect 4340 53900 4452 53956
rect 4284 53862 4340 53900
rect 3388 53678 3390 53730
rect 3442 53678 3444 53730
rect 3388 53666 3444 53678
rect 3836 53730 3892 53742
rect 3836 53678 3838 53730
rect 3890 53678 3892 53730
rect 3836 53620 3892 53678
rect 4284 53620 4340 53630
rect 3836 53618 4340 53620
rect 3836 53566 4286 53618
rect 4338 53566 4340 53618
rect 3836 53564 4340 53566
rect 4284 52724 4340 53564
rect 4396 53618 4452 53900
rect 4620 53900 4900 53956
rect 4620 53730 4676 53900
rect 4620 53678 4622 53730
rect 4674 53678 4676 53730
rect 4620 53666 4676 53678
rect 4396 53566 4398 53618
rect 4450 53566 4452 53618
rect 4396 53554 4452 53566
rect 4284 52658 4340 52668
rect 4956 52724 5012 54462
rect 5180 54516 5236 54526
rect 5180 54422 5236 54460
rect 5068 53844 5124 53854
rect 5292 53844 5348 56700
rect 6188 56642 6244 57036
rect 6748 56866 6804 56878
rect 6748 56814 6750 56866
rect 6802 56814 6804 56866
rect 6636 56756 6692 56766
rect 6748 56756 6804 56814
rect 6860 56868 6916 57596
rect 6860 56802 6916 56812
rect 6692 56700 6804 56756
rect 6636 56690 6692 56700
rect 6188 56590 6190 56642
rect 6242 56590 6244 56642
rect 6188 55524 6244 56590
rect 6188 55458 6244 55468
rect 6636 55636 6692 55646
rect 5068 53842 5348 53844
rect 5068 53790 5070 53842
rect 5122 53790 5348 53842
rect 5068 53788 5348 53790
rect 5404 54628 5460 54638
rect 5068 53778 5124 53788
rect 4956 52658 5012 52668
rect 5292 52946 5348 52958
rect 5292 52894 5294 52946
rect 5346 52894 5348 52946
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3948 52276 4004 52286
rect 3948 51604 4004 52220
rect 4620 52276 4676 52286
rect 4620 52182 4676 52220
rect 3836 51602 4004 51604
rect 3836 51550 3950 51602
rect 4002 51550 4004 51602
rect 3836 51548 4004 51550
rect 3388 51492 3444 51502
rect 3276 51378 3332 51390
rect 3276 51326 3278 51378
rect 3330 51326 3332 51378
rect 3276 51268 3332 51326
rect 3276 51202 3332 51212
rect 2492 50482 2548 50494
rect 2492 50430 2494 50482
rect 2546 50430 2548 50482
rect 2492 50036 2548 50430
rect 2492 49970 2548 49980
rect 3388 49810 3444 51436
rect 3612 51378 3668 51390
rect 3612 51326 3614 51378
rect 3666 51326 3668 51378
rect 3612 50596 3668 51326
rect 3612 50530 3668 50540
rect 3388 49758 3390 49810
rect 3442 49758 3444 49810
rect 3388 49746 3444 49758
rect 2492 47348 2548 47358
rect 2492 47346 2660 47348
rect 2492 47294 2494 47346
rect 2546 47294 2660 47346
rect 2492 47292 2660 47294
rect 2492 47282 2548 47292
rect 2604 46898 2660 47292
rect 2604 46846 2606 46898
rect 2658 46846 2660 46898
rect 2604 46834 2660 46846
rect 2492 46786 2548 46798
rect 2492 46734 2494 46786
rect 2546 46734 2548 46786
rect 2492 46116 2548 46734
rect 2716 46564 2772 46574
rect 2716 46470 2772 46508
rect 3388 46564 3444 46574
rect 3388 46470 3444 46508
rect 2492 46060 2996 46116
rect 2492 44324 2548 46060
rect 2940 46004 2996 46060
rect 2940 46002 3108 46004
rect 2940 45950 2942 46002
rect 2994 45950 3108 46002
rect 2940 45948 3108 45950
rect 2940 45938 2996 45948
rect 3052 45330 3108 45948
rect 3052 45278 3054 45330
rect 3106 45278 3108 45330
rect 3052 45266 3108 45278
rect 3500 44546 3556 44558
rect 3500 44494 3502 44546
rect 3554 44494 3556 44546
rect 2156 43652 2324 43708
rect 2380 44322 2548 44324
rect 2380 44270 2494 44322
rect 2546 44270 2548 44322
rect 2380 44268 2548 44270
rect 2380 43764 2436 44268
rect 2492 44258 2548 44268
rect 3388 44436 3444 44446
rect 3500 44436 3556 44494
rect 3500 44380 3780 44436
rect 2828 44210 2884 44222
rect 2828 44158 2830 44210
rect 2882 44158 2884 44210
rect 2716 44100 2772 44110
rect 2380 43698 2436 43708
rect 2492 44098 2772 44100
rect 2492 44046 2718 44098
rect 2770 44046 2772 44098
rect 2492 44044 2772 44046
rect 1820 43540 1876 43550
rect 1820 43446 1876 43484
rect 1820 39732 1876 39742
rect 1820 39618 1876 39676
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 36482 1876 39566
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 36418 1876 36430
rect 1820 35698 1876 35710
rect 1820 35646 1822 35698
rect 1874 35646 1876 35698
rect 1820 35028 1876 35646
rect 1820 34934 1876 34972
rect 2156 31948 2212 43652
rect 2492 43650 2548 44044
rect 2716 44034 2772 44044
rect 2492 43598 2494 43650
rect 2546 43598 2548 43650
rect 2492 43586 2548 43598
rect 2604 43764 2660 43774
rect 2604 41748 2660 43708
rect 2828 42868 2884 44158
rect 3388 44212 3444 44380
rect 3500 44212 3556 44222
rect 3388 44210 3556 44212
rect 3388 44158 3502 44210
rect 3554 44158 3556 44210
rect 3388 44156 3556 44158
rect 3500 44146 3556 44156
rect 3612 44210 3668 44222
rect 3612 44158 3614 44210
rect 3666 44158 3668 44210
rect 3612 43540 3668 44158
rect 3612 43474 3668 43484
rect 3612 42980 3668 42990
rect 2940 42868 2996 42878
rect 2828 42866 2996 42868
rect 2828 42814 2942 42866
rect 2994 42814 2996 42866
rect 2828 42812 2996 42814
rect 2940 42802 2996 42812
rect 3612 42754 3668 42924
rect 3724 42866 3780 44380
rect 3724 42814 3726 42866
rect 3778 42814 3780 42866
rect 3724 42802 3780 42814
rect 3612 42702 3614 42754
rect 3666 42702 3668 42754
rect 3276 41858 3332 41870
rect 3276 41806 3278 41858
rect 3330 41806 3332 41858
rect 2828 41748 2884 41758
rect 2604 41692 2828 41748
rect 2716 41300 2772 41310
rect 2492 41298 2772 41300
rect 2492 41246 2718 41298
rect 2770 41246 2772 41298
rect 2492 41244 2772 41246
rect 2492 39730 2548 41244
rect 2716 41234 2772 41244
rect 2828 41074 2884 41692
rect 3276 41748 3332 41806
rect 3276 41682 3332 41692
rect 3052 41076 3108 41086
rect 2828 41022 2830 41074
rect 2882 41022 2884 41074
rect 2828 41010 2884 41022
rect 2940 41074 3108 41076
rect 2940 41022 3054 41074
rect 3106 41022 3108 41074
rect 2940 41020 3108 41022
rect 3612 41076 3668 42702
rect 3836 42756 3892 51548
rect 3948 51538 4004 51548
rect 5068 51492 5124 51502
rect 4172 51378 4228 51390
rect 4172 51326 4174 51378
rect 4226 51326 4228 51378
rect 3948 51268 4004 51278
rect 3948 50708 4004 51212
rect 3948 49810 4004 50652
rect 4172 50484 4228 51326
rect 4396 51380 4452 51390
rect 4396 51286 4452 51324
rect 5068 51378 5124 51436
rect 5068 51326 5070 51378
rect 5122 51326 5124 51378
rect 4284 51266 4340 51278
rect 4284 51214 4286 51266
rect 4338 51214 4340 51266
rect 4284 50596 4340 51214
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5068 50818 5124 51326
rect 5068 50766 5070 50818
rect 5122 50766 5124 50818
rect 5068 50754 5124 50766
rect 4620 50708 4676 50718
rect 4620 50706 5012 50708
rect 4620 50654 4622 50706
rect 4674 50654 5012 50706
rect 4620 50652 5012 50654
rect 4620 50642 4676 50652
rect 4284 50540 4564 50596
rect 4172 50418 4228 50428
rect 4508 50428 4564 50540
rect 4956 50594 5012 50652
rect 4956 50542 4958 50594
rect 5010 50542 5012 50594
rect 4956 50530 5012 50542
rect 5292 50428 5348 52894
rect 5404 51490 5460 54572
rect 5964 53508 6020 53518
rect 5964 53058 6020 53452
rect 5964 53006 5966 53058
rect 6018 53006 6020 53058
rect 5964 52994 6020 53006
rect 5404 51438 5406 51490
rect 5458 51438 5460 51490
rect 5404 51426 5460 51438
rect 5740 51378 5796 51390
rect 5740 51326 5742 51378
rect 5794 51326 5796 51378
rect 5516 51266 5572 51278
rect 5516 51214 5518 51266
rect 5570 51214 5572 51266
rect 5516 50708 5572 51214
rect 5740 50818 5796 51326
rect 5740 50766 5742 50818
rect 5794 50766 5796 50818
rect 5740 50754 5796 50766
rect 5516 50642 5572 50652
rect 5628 50596 5684 50606
rect 5628 50502 5684 50540
rect 5740 50484 5796 50522
rect 4284 50372 4340 50382
rect 4508 50372 4900 50428
rect 5292 50372 5460 50428
rect 5740 50418 5796 50428
rect 4060 49924 4116 49934
rect 4284 49924 4340 50316
rect 4732 50260 4788 50270
rect 4508 50036 4564 50046
rect 4508 49942 4564 49980
rect 4060 49922 4340 49924
rect 4060 49870 4062 49922
rect 4114 49870 4340 49922
rect 4060 49868 4340 49870
rect 4060 49858 4116 49868
rect 3948 49758 3950 49810
rect 4002 49758 4004 49810
rect 3948 49746 4004 49758
rect 4284 49810 4340 49868
rect 4284 49758 4286 49810
rect 4338 49758 4340 49810
rect 4284 49746 4340 49758
rect 4732 49810 4788 50204
rect 4732 49758 4734 49810
rect 4786 49758 4788 49810
rect 4732 49588 4788 49758
rect 4844 49810 4900 50372
rect 4844 49758 4846 49810
rect 4898 49758 4900 49810
rect 4844 49746 4900 49758
rect 5404 49698 5460 50372
rect 5404 49646 5406 49698
rect 5458 49646 5460 49698
rect 4732 49532 4900 49588
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4844 48354 4900 49532
rect 5404 49028 5460 49646
rect 4844 48302 4846 48354
rect 4898 48302 4900 48354
rect 4844 48290 4900 48302
rect 5068 48972 5404 49028
rect 4620 48242 4676 48254
rect 4620 48190 4622 48242
rect 4674 48190 4676 48242
rect 4620 48020 4676 48190
rect 4956 48132 5012 48142
rect 4956 48038 5012 48076
rect 4284 47964 4676 48020
rect 4060 46676 4116 46686
rect 4284 46676 4340 47964
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4620 47570 4676 47582
rect 4620 47518 4622 47570
rect 4674 47518 4676 47570
rect 4620 47348 4676 47518
rect 5068 47572 5124 48972
rect 5404 48962 5460 48972
rect 6076 49028 6132 49038
rect 6076 48934 6132 48972
rect 5852 48356 5908 48366
rect 5516 48354 5908 48356
rect 5516 48302 5854 48354
rect 5906 48302 5908 48354
rect 5516 48300 5908 48302
rect 5516 48242 5572 48300
rect 5852 48290 5908 48300
rect 6076 48354 6132 48366
rect 6076 48302 6078 48354
rect 6130 48302 6132 48354
rect 5516 48190 5518 48242
rect 5570 48190 5572 48242
rect 5516 48178 5572 48190
rect 5628 48132 5684 48142
rect 5628 47682 5684 48076
rect 5628 47630 5630 47682
rect 5682 47630 5684 47682
rect 5628 47618 5684 47630
rect 6076 47572 6132 48302
rect 5124 47516 5572 47572
rect 5068 47478 5124 47516
rect 4620 47282 4676 47292
rect 5292 47348 5348 47358
rect 5292 46786 5348 47292
rect 5292 46734 5294 46786
rect 5346 46734 5348 46786
rect 5292 46722 5348 46734
rect 5404 47012 5460 47022
rect 4060 46674 4340 46676
rect 4060 46622 4062 46674
rect 4114 46622 4340 46674
rect 4060 46620 4340 46622
rect 4060 44434 4116 46620
rect 5404 46562 5460 46956
rect 5404 46510 5406 46562
rect 5458 46510 5460 46562
rect 5404 46498 5460 46510
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4956 45220 5012 45230
rect 4844 45218 5012 45220
rect 4844 45166 4958 45218
rect 5010 45166 5012 45218
rect 4844 45164 5012 45166
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4060 44382 4062 44434
rect 4114 44382 4116 44434
rect 4060 44370 4116 44382
rect 4508 44436 4564 44446
rect 4508 44322 4564 44380
rect 4508 44270 4510 44322
rect 4562 44270 4564 44322
rect 4508 44258 4564 44270
rect 4844 44324 4900 45164
rect 4956 45154 5012 45164
rect 5068 45108 5124 45118
rect 5068 45106 5236 45108
rect 5068 45054 5070 45106
rect 5122 45054 5236 45106
rect 5068 45052 5236 45054
rect 5068 45042 5124 45052
rect 4956 44882 5012 44894
rect 4956 44830 4958 44882
rect 5010 44830 5012 44882
rect 4956 44548 5012 44830
rect 5180 44548 5236 45052
rect 4956 44492 5124 44548
rect 3948 44210 4004 44222
rect 3948 44158 3950 44210
rect 4002 44158 4004 44210
rect 3948 42980 4004 44158
rect 4620 43428 4676 43438
rect 4844 43428 4900 44268
rect 4956 44322 5012 44334
rect 4956 44270 4958 44322
rect 5010 44270 5012 44322
rect 4956 43762 5012 44270
rect 4956 43710 4958 43762
rect 5010 43710 5012 43762
rect 4956 43698 5012 43710
rect 5068 43650 5124 44492
rect 5180 44482 5236 44492
rect 5516 43652 5572 47516
rect 5740 47516 6132 47572
rect 6188 48242 6244 48254
rect 6188 48190 6190 48242
rect 6242 48190 6244 48242
rect 5740 47348 5796 47516
rect 5740 47254 5796 47292
rect 5964 47348 6020 47358
rect 6188 47348 6244 48190
rect 5964 47346 6244 47348
rect 5964 47294 5966 47346
rect 6018 47294 6244 47346
rect 5964 47292 6244 47294
rect 5964 47282 6020 47292
rect 6188 47012 6244 47292
rect 6188 46946 6244 46956
rect 6076 45108 6132 45118
rect 6076 45014 6132 45052
rect 5628 44436 5684 44446
rect 5628 44342 5684 44380
rect 5964 44436 6020 44446
rect 5964 44342 6020 44380
rect 6188 44324 6244 44334
rect 6188 44230 6244 44268
rect 5068 43598 5070 43650
rect 5122 43598 5124 43650
rect 5068 43540 5124 43598
rect 5068 43474 5124 43484
rect 5404 43596 5516 43652
rect 4620 43426 4900 43428
rect 4620 43374 4622 43426
rect 4674 43374 4900 43426
rect 4620 43372 4900 43374
rect 4620 43362 4676 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 3948 42914 4004 42924
rect 3836 42700 4228 42756
rect 4060 41186 4116 41198
rect 4060 41134 4062 41186
rect 4114 41134 4116 41186
rect 3724 41076 3780 41086
rect 3612 41074 3780 41076
rect 3612 41022 3726 41074
rect 3778 41022 3780 41074
rect 3612 41020 3780 41022
rect 2716 40628 2772 40638
rect 2940 40628 2996 41020
rect 3052 41010 3108 41020
rect 3724 41010 3780 41020
rect 2716 40626 2996 40628
rect 2716 40574 2718 40626
rect 2770 40574 2996 40626
rect 2716 40572 2996 40574
rect 2716 40562 2772 40572
rect 3052 40516 3108 40526
rect 3052 40402 3108 40460
rect 4060 40516 4116 41134
rect 3052 40350 3054 40402
rect 3106 40350 3108 40402
rect 3052 40338 3108 40350
rect 3948 40404 4004 40414
rect 3948 40310 4004 40348
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 3948 38276 4004 38286
rect 4060 38276 4116 40460
rect 4172 38724 4228 42700
rect 5404 41970 5460 43596
rect 5516 43558 5572 43596
rect 5404 41918 5406 41970
rect 5458 41918 5460 41970
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4508 41300 4564 41310
rect 4508 41298 5012 41300
rect 4508 41246 4510 41298
rect 4562 41246 5012 41298
rect 4508 41244 5012 41246
rect 4508 41234 4564 41244
rect 4284 40964 4340 40974
rect 4284 40514 4340 40908
rect 4284 40462 4286 40514
rect 4338 40462 4340 40514
rect 4284 39844 4340 40462
rect 4956 40290 5012 41244
rect 5180 41188 5236 41198
rect 5180 41094 5236 41132
rect 5292 41076 5348 41086
rect 5068 40964 5124 40974
rect 5068 40626 5124 40908
rect 5068 40574 5070 40626
rect 5122 40574 5124 40626
rect 5068 40562 5124 40574
rect 5292 40514 5348 41020
rect 5292 40462 5294 40514
rect 5346 40462 5348 40514
rect 5292 40404 5348 40462
rect 5292 40338 5348 40348
rect 4956 40238 4958 40290
rect 5010 40238 5012 40290
rect 4956 40226 5012 40238
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 39788 4676 39844
rect 4620 39730 4676 39788
rect 4620 39678 4622 39730
rect 4674 39678 4676 39730
rect 4620 39666 4676 39678
rect 5068 39732 5124 39742
rect 5068 38668 5124 39676
rect 5404 39732 5460 41918
rect 6076 42532 6132 42542
rect 6076 41970 6132 42476
rect 6076 41918 6078 41970
rect 6130 41918 6132 41970
rect 6076 41906 6132 41918
rect 5516 41188 5572 41198
rect 5516 41094 5572 41132
rect 5852 41076 5908 41086
rect 5852 40982 5908 41020
rect 5740 40964 5796 40974
rect 5740 40870 5796 40908
rect 6636 39732 6692 55580
rect 7196 55636 7252 59612
rect 7644 59444 7700 59454
rect 7644 59350 7700 59388
rect 7532 59332 7588 59342
rect 7532 59238 7588 59276
rect 7756 59332 7812 59342
rect 7868 59332 7924 60958
rect 8428 60004 8484 60014
rect 8652 60004 8708 63868
rect 8764 63858 8820 63868
rect 8988 64482 9044 64494
rect 8988 64430 8990 64482
rect 9042 64430 9044 64482
rect 8988 63028 9044 64430
rect 11340 64146 11396 64540
rect 11340 64094 11342 64146
rect 11394 64094 11396 64146
rect 11340 64082 11396 64094
rect 11676 63922 11732 63934
rect 11676 63870 11678 63922
rect 11730 63870 11732 63922
rect 8988 62972 9604 63028
rect 8764 62356 8820 62366
rect 9436 62356 9492 62366
rect 8764 62354 9492 62356
rect 8764 62302 8766 62354
rect 8818 62302 9438 62354
rect 9490 62302 9492 62354
rect 8764 62300 9492 62302
rect 8764 62290 8820 62300
rect 9436 62290 9492 62300
rect 9548 62356 9604 62972
rect 10556 62468 10612 62478
rect 9548 62290 9604 62300
rect 10220 62356 10276 62366
rect 10220 62262 10276 62300
rect 10556 62242 10612 62412
rect 10892 62468 10948 62478
rect 10892 62374 10948 62412
rect 11676 62356 11732 63870
rect 12236 63924 12292 64766
rect 12684 64708 12740 65324
rect 13244 65378 13300 65390
rect 13244 65326 13246 65378
rect 13298 65326 13300 65378
rect 12796 64820 12852 64830
rect 12796 64726 12852 64764
rect 12684 64642 12740 64652
rect 12572 64596 12628 64606
rect 12572 64502 12628 64540
rect 12796 64484 12852 64494
rect 13244 64484 13300 65326
rect 17388 65378 17444 66220
rect 17612 66210 17668 66220
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 20188 65492 20244 65502
rect 17388 65326 17390 65378
rect 17442 65326 17444 65378
rect 17388 65314 17444 65326
rect 17612 65380 17668 65390
rect 16380 64818 16436 64830
rect 16380 64766 16382 64818
rect 16434 64766 16436 64818
rect 13580 64708 13636 64718
rect 13580 64614 13636 64652
rect 14252 64596 14308 64606
rect 14252 64594 14980 64596
rect 14252 64542 14254 64594
rect 14306 64542 14980 64594
rect 14252 64540 14980 64542
rect 14252 64530 14308 64540
rect 12684 64482 13300 64484
rect 12684 64430 12798 64482
rect 12850 64430 13300 64482
rect 12684 64428 13300 64430
rect 12236 63858 12292 63868
rect 12572 64148 12628 64158
rect 12572 63922 12628 64092
rect 12572 63870 12574 63922
rect 12626 63870 12628 63922
rect 12572 63026 12628 63870
rect 12572 62974 12574 63026
rect 12626 62974 12628 63026
rect 11900 62356 11956 62366
rect 11676 62300 11900 62356
rect 10556 62190 10558 62242
rect 10610 62190 10612 62242
rect 10220 60788 10276 60798
rect 8428 60002 8708 60004
rect 8428 59950 8430 60002
rect 8482 59950 8708 60002
rect 8428 59948 8708 59950
rect 9100 60004 9156 60014
rect 8428 59780 8484 59948
rect 9100 59910 9156 59948
rect 8428 59714 8484 59724
rect 7756 59330 7924 59332
rect 7756 59278 7758 59330
rect 7810 59278 7924 59330
rect 7756 59276 7924 59278
rect 8204 59332 8260 59342
rect 7756 59266 7812 59276
rect 8204 59238 8260 59276
rect 10220 58548 10276 60732
rect 10556 60116 10612 62190
rect 11788 61684 11844 61694
rect 11788 61012 11844 61628
rect 11676 60956 11844 61012
rect 11004 60900 11060 60910
rect 10780 60788 10836 60798
rect 10780 60694 10836 60732
rect 10556 60050 10612 60060
rect 11004 60004 11060 60844
rect 11564 60788 11620 60798
rect 11116 60786 11620 60788
rect 11116 60734 11566 60786
rect 11618 60734 11620 60786
rect 11116 60732 11620 60734
rect 11116 60674 11172 60732
rect 11564 60722 11620 60732
rect 11116 60622 11118 60674
rect 11170 60622 11172 60674
rect 11116 60610 11172 60622
rect 11228 60114 11284 60126
rect 11228 60062 11230 60114
rect 11282 60062 11284 60114
rect 11228 60004 11284 60062
rect 10668 59948 11284 60004
rect 11676 60002 11732 60956
rect 11900 60898 11956 62300
rect 12236 61684 12292 61694
rect 12236 61590 12292 61628
rect 11900 60846 11902 60898
rect 11954 60846 11956 60898
rect 11900 60834 11956 60846
rect 11788 60786 11844 60798
rect 11788 60734 11790 60786
rect 11842 60734 11844 60786
rect 11788 60340 11844 60734
rect 12572 60564 12628 62974
rect 12684 61684 12740 64428
rect 12796 64418 12852 64428
rect 13804 64148 13860 64158
rect 12796 64036 12852 64046
rect 12796 63026 12852 63980
rect 12908 64034 12964 64046
rect 12908 63982 12910 64034
rect 12962 63982 12964 64034
rect 12908 63924 12964 63982
rect 13692 64036 13748 64046
rect 13692 63942 13748 63980
rect 13804 64034 13860 64092
rect 13804 63982 13806 64034
rect 13858 63982 13860 64034
rect 13804 63970 13860 63982
rect 14140 64036 14196 64046
rect 14140 63942 14196 63980
rect 12908 63858 12964 63868
rect 14252 63924 14308 63934
rect 14252 63830 14308 63868
rect 13692 63698 13748 63710
rect 13692 63646 13694 63698
rect 13746 63646 13748 63698
rect 12796 62974 12798 63026
rect 12850 62974 12852 63026
rect 12796 62962 12852 62974
rect 12908 63250 12964 63262
rect 12908 63198 12910 63250
rect 12962 63198 12964 63250
rect 12908 62354 12964 63198
rect 13132 63140 13188 63150
rect 13132 62578 13188 63084
rect 13132 62526 13134 62578
rect 13186 62526 13188 62578
rect 13132 62514 13188 62526
rect 12908 62302 12910 62354
rect 12962 62302 12964 62354
rect 12908 62290 12964 62302
rect 13580 62466 13636 62478
rect 13580 62414 13582 62466
rect 13634 62414 13636 62466
rect 13580 62356 13636 62414
rect 13580 62290 13636 62300
rect 13692 62354 13748 63646
rect 14812 63026 14868 63038
rect 14812 62974 14814 63026
rect 14866 62974 14868 63026
rect 14812 62466 14868 62974
rect 14924 62578 14980 64540
rect 15484 63140 15540 63150
rect 15484 63046 15540 63084
rect 16268 63138 16324 63150
rect 16268 63086 16270 63138
rect 16322 63086 16324 63138
rect 14924 62526 14926 62578
rect 14978 62526 14980 62578
rect 14924 62514 14980 62526
rect 16268 62916 16324 63086
rect 16380 63028 16436 64766
rect 16828 64708 16884 64718
rect 16828 64614 16884 64652
rect 17612 64146 17668 65324
rect 19516 65380 19572 65390
rect 19516 65286 19572 65324
rect 17948 64708 18004 64718
rect 17948 64614 18004 64652
rect 20188 64708 20244 65436
rect 20860 65492 20916 65502
rect 20860 65378 20916 65436
rect 20860 65326 20862 65378
rect 20914 65326 20916 65378
rect 18620 64596 18676 64606
rect 18620 64594 19684 64596
rect 18620 64542 18622 64594
rect 18674 64542 19684 64594
rect 18620 64540 19684 64542
rect 18620 64530 18676 64540
rect 17612 64094 17614 64146
rect 17666 64094 17668 64146
rect 17612 64082 17668 64094
rect 16716 63924 16772 63934
rect 16492 63028 16548 63038
rect 16380 63026 16492 63028
rect 16380 62974 16382 63026
rect 16434 62974 16492 63026
rect 16380 62972 16492 62974
rect 16380 62962 16436 62972
rect 14812 62414 14814 62466
rect 14866 62414 14868 62466
rect 14812 62402 14868 62414
rect 13692 62302 13694 62354
rect 13746 62302 13748 62354
rect 13692 62290 13748 62302
rect 15148 62354 15204 62366
rect 15148 62302 15150 62354
rect 15202 62302 15204 62354
rect 15148 62244 15204 62302
rect 16268 62356 16324 62860
rect 16492 62578 16548 62972
rect 16492 62526 16494 62578
rect 16546 62526 16548 62578
rect 16492 62514 16548 62526
rect 16716 62578 16772 63868
rect 17276 63922 17332 63934
rect 17276 63870 17278 63922
rect 17330 63870 17332 63922
rect 17276 63140 17332 63870
rect 17612 63924 17668 63934
rect 17612 63830 17668 63868
rect 17836 63922 17892 63934
rect 17836 63870 17838 63922
rect 17890 63870 17892 63922
rect 17836 63476 17892 63870
rect 17500 63420 17892 63476
rect 17500 63250 17556 63420
rect 19628 63362 19684 64540
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 20188 63922 20244 64652
rect 20748 64818 20804 64830
rect 20748 64766 20750 64818
rect 20802 64766 20804 64818
rect 20748 64036 20804 64766
rect 20860 64484 20916 65326
rect 20860 64418 20916 64428
rect 20748 63980 21028 64036
rect 20188 63870 20190 63922
rect 20242 63870 20244 63922
rect 20188 63858 20244 63870
rect 19628 63310 19630 63362
rect 19682 63310 19684 63362
rect 19628 63298 19684 63310
rect 20860 63810 20916 63822
rect 20860 63758 20862 63810
rect 20914 63758 20916 63810
rect 17500 63198 17502 63250
rect 17554 63198 17556 63250
rect 17500 63186 17556 63198
rect 17276 63074 17332 63084
rect 18060 63140 18116 63150
rect 19628 63140 19684 63150
rect 18060 63138 18564 63140
rect 18060 63086 18062 63138
rect 18114 63086 18564 63138
rect 18060 63084 18564 63086
rect 18060 63074 18116 63084
rect 17612 63028 17668 63038
rect 17612 62934 17668 62972
rect 17388 62916 17444 62926
rect 17388 62822 17444 62860
rect 17948 62916 18004 62926
rect 16716 62526 16718 62578
rect 16770 62526 16772 62578
rect 16716 62514 16772 62526
rect 16380 62356 16436 62366
rect 16268 62354 16436 62356
rect 16268 62302 16382 62354
rect 16434 62302 16436 62354
rect 16268 62300 16436 62302
rect 15596 62244 15652 62254
rect 15148 62242 15652 62244
rect 15148 62190 15598 62242
rect 15650 62190 15652 62242
rect 15148 62188 15652 62190
rect 12684 61618 12740 61628
rect 15596 61684 15652 62188
rect 16380 61684 16436 62300
rect 13244 60900 13300 60910
rect 13244 60806 13300 60844
rect 12796 60788 12852 60798
rect 13020 60788 13076 60798
rect 12796 60786 13076 60788
rect 12796 60734 12798 60786
rect 12850 60734 13022 60786
rect 13074 60734 13076 60786
rect 12796 60732 13076 60734
rect 12796 60722 12852 60732
rect 13020 60722 13076 60732
rect 13356 60788 13412 60798
rect 13356 60694 13412 60732
rect 13916 60674 13972 60686
rect 14252 60676 14308 60686
rect 13916 60622 13918 60674
rect 13970 60622 13972 60674
rect 12572 60498 12628 60508
rect 13804 60564 13860 60574
rect 11788 60284 11956 60340
rect 11676 59950 11678 60002
rect 11730 59950 11732 60002
rect 10220 58546 10612 58548
rect 10220 58494 10222 58546
rect 10274 58494 10612 58546
rect 10220 58492 10612 58494
rect 10220 58482 10276 58492
rect 10556 58100 10612 58492
rect 10668 58322 10724 59948
rect 11676 59938 11732 59950
rect 11788 60114 11844 60126
rect 11788 60062 11790 60114
rect 11842 60062 11844 60114
rect 11788 60004 11844 60062
rect 11788 59938 11844 59948
rect 11340 59780 11396 59790
rect 11340 59442 11396 59724
rect 11340 59390 11342 59442
rect 11394 59390 11396 59442
rect 11340 59378 11396 59390
rect 11788 58436 11844 58446
rect 11900 58436 11956 60284
rect 12796 60116 12852 60126
rect 12796 60022 12852 60060
rect 12460 60004 12516 60014
rect 11788 58434 11956 58436
rect 11788 58382 11790 58434
rect 11842 58382 11956 58434
rect 11788 58380 11956 58382
rect 12012 59890 12068 59902
rect 12012 59838 12014 59890
rect 12066 59838 12068 59890
rect 10668 58270 10670 58322
rect 10722 58270 10724 58322
rect 10668 58258 10724 58270
rect 11004 58324 11060 58334
rect 10556 58044 10836 58100
rect 9884 57876 9940 57886
rect 10556 57876 10612 57886
rect 9548 57874 10612 57876
rect 9548 57822 9886 57874
rect 9938 57822 10558 57874
rect 10610 57822 10612 57874
rect 9548 57820 10612 57822
rect 7980 57764 8036 57774
rect 7980 57762 8260 57764
rect 7980 57710 7982 57762
rect 8034 57710 8260 57762
rect 7980 57708 8260 57710
rect 7980 57698 8036 57708
rect 8092 57538 8148 57550
rect 8092 57486 8094 57538
rect 8146 57486 8148 57538
rect 8092 57204 8148 57486
rect 7420 57148 8148 57204
rect 7420 56978 7476 57148
rect 7420 56926 7422 56978
rect 7474 56926 7476 56978
rect 7420 56914 7476 56926
rect 8204 56308 8260 57708
rect 8316 57652 8372 57662
rect 8428 57652 8484 57662
rect 8316 57650 8428 57652
rect 8316 57598 8318 57650
rect 8370 57598 8428 57650
rect 8316 57596 8428 57598
rect 8316 57586 8372 57596
rect 8204 56242 8260 56252
rect 8316 56196 8372 56206
rect 8316 56102 8372 56140
rect 8428 56084 8484 57596
rect 8540 57652 8596 57662
rect 9436 57652 9492 57662
rect 8540 57650 8708 57652
rect 8540 57598 8542 57650
rect 8594 57598 8708 57650
rect 8540 57596 8708 57598
rect 8540 57586 8596 57596
rect 8652 56306 8708 57596
rect 9436 57558 9492 57596
rect 9548 56978 9604 57820
rect 9884 57810 9940 57820
rect 10108 57652 10164 57662
rect 10332 57652 10388 57662
rect 10108 57558 10164 57596
rect 10220 57650 10388 57652
rect 10220 57598 10334 57650
rect 10386 57598 10388 57650
rect 10220 57596 10388 57598
rect 9996 57538 10052 57550
rect 9996 57486 9998 57538
rect 10050 57486 10052 57538
rect 9996 57092 10052 57486
rect 9996 57026 10052 57036
rect 9548 56926 9550 56978
rect 9602 56926 9604 56978
rect 9548 56914 9604 56926
rect 9772 56756 9828 56766
rect 8652 56254 8654 56306
rect 8706 56254 8708 56306
rect 8652 56242 8708 56254
rect 8764 56308 8820 56318
rect 8764 56214 8820 56252
rect 9772 56306 9828 56700
rect 9772 56254 9774 56306
rect 9826 56254 9828 56306
rect 9772 56242 9828 56254
rect 9884 56754 9940 56766
rect 9884 56702 9886 56754
rect 9938 56702 9940 56754
rect 9884 56308 9940 56702
rect 9884 56242 9940 56252
rect 8988 56196 9044 56206
rect 9044 56140 9156 56196
rect 8988 56130 9044 56140
rect 8540 56084 8596 56094
rect 8428 56082 8596 56084
rect 8428 56030 8542 56082
rect 8594 56030 8596 56082
rect 8428 56028 8596 56030
rect 7196 55570 7252 55580
rect 6860 54404 6916 54414
rect 6860 52276 6916 54348
rect 8540 53956 8596 56028
rect 8988 53956 9044 53966
rect 8540 53954 9044 53956
rect 8540 53902 8990 53954
rect 9042 53902 9044 53954
rect 8540 53900 9044 53902
rect 8988 53890 9044 53900
rect 8428 53732 8484 53742
rect 8876 53732 8932 53742
rect 8428 53730 8932 53732
rect 8428 53678 8430 53730
rect 8482 53678 8878 53730
rect 8930 53678 8932 53730
rect 8428 53676 8932 53678
rect 8428 53666 8484 53676
rect 8876 53666 8932 53676
rect 7084 53618 7140 53630
rect 7084 53566 7086 53618
rect 7138 53566 7140 53618
rect 7084 52836 7140 53566
rect 7420 53618 7476 53630
rect 7420 53566 7422 53618
rect 7474 53566 7476 53618
rect 7196 53508 7252 53518
rect 7196 53414 7252 53452
rect 7420 53508 7476 53566
rect 7420 53442 7476 53452
rect 7644 53618 7700 53630
rect 7644 53566 7646 53618
rect 7698 53566 7700 53618
rect 7644 53172 7700 53566
rect 8092 53508 8148 53518
rect 8316 53508 8372 53518
rect 8540 53508 8596 53518
rect 8092 53414 8148 53452
rect 8204 53506 8372 53508
rect 8204 53454 8318 53506
rect 8370 53454 8372 53506
rect 8204 53452 8372 53454
rect 7644 53106 7700 53116
rect 7308 52836 7364 52846
rect 8092 52836 8148 52846
rect 8204 52836 8260 53452
rect 8316 53442 8372 53452
rect 8428 53506 8596 53508
rect 8428 53454 8542 53506
rect 8594 53454 8596 53506
rect 8428 53452 8596 53454
rect 8428 53284 8484 53452
rect 8540 53442 8596 53452
rect 8652 53508 8708 53518
rect 7084 52780 7308 52836
rect 6860 52210 6916 52220
rect 7308 52274 7364 52780
rect 7308 52222 7310 52274
rect 7362 52222 7364 52274
rect 7308 52210 7364 52222
rect 7980 52834 8260 52836
rect 7980 52782 8094 52834
rect 8146 52782 8260 52834
rect 7980 52780 8260 52782
rect 8316 53228 8484 53284
rect 7980 52162 8036 52780
rect 8092 52770 8148 52780
rect 8204 52500 8260 52510
rect 8316 52500 8372 53228
rect 8540 53172 8596 53182
rect 8540 53078 8596 53116
rect 8428 52946 8484 52958
rect 8652 52948 8708 53452
rect 8988 53506 9044 53518
rect 8988 53454 8990 53506
rect 9042 53454 9044 53506
rect 8988 53172 9044 53454
rect 8428 52894 8430 52946
rect 8482 52894 8484 52946
rect 8428 52836 8484 52894
rect 8428 52770 8484 52780
rect 8540 52946 8708 52948
rect 8540 52894 8654 52946
rect 8706 52894 8708 52946
rect 8540 52892 8708 52894
rect 8260 52444 8372 52500
rect 8204 52274 8260 52444
rect 8204 52222 8206 52274
rect 8258 52222 8260 52274
rect 8204 52210 8260 52222
rect 7980 52110 7982 52162
rect 8034 52110 8036 52162
rect 7980 52052 8036 52110
rect 7980 51986 8036 51996
rect 8540 50484 8596 52892
rect 8652 52882 8708 52892
rect 8764 53116 9044 53172
rect 8652 52500 8708 52510
rect 8652 52162 8708 52444
rect 8764 52386 8820 53116
rect 9100 52948 9156 56140
rect 10220 56082 10276 57596
rect 10332 57586 10388 57596
rect 10220 56030 10222 56082
rect 10274 56030 10276 56082
rect 10220 56018 10276 56030
rect 10444 57092 10500 57102
rect 10444 56082 10500 57036
rect 10556 56866 10612 57820
rect 10556 56814 10558 56866
rect 10610 56814 10612 56866
rect 10556 56802 10612 56814
rect 10668 57652 10724 57662
rect 10668 56978 10724 57596
rect 10780 57092 10836 58044
rect 10780 57026 10836 57036
rect 10668 56926 10670 56978
rect 10722 56926 10724 56978
rect 10444 56030 10446 56082
rect 10498 56030 10500 56082
rect 10444 56018 10500 56030
rect 10332 55524 10388 55534
rect 10332 53618 10388 55468
rect 10668 54740 10724 56926
rect 10780 56308 10836 56318
rect 11004 56308 11060 58268
rect 11788 58324 11844 58380
rect 11788 58258 11844 58268
rect 12012 58210 12068 59838
rect 12236 59218 12292 59230
rect 12236 59166 12238 59218
rect 12290 59166 12292 59218
rect 12236 58884 12292 59166
rect 12236 58818 12292 58828
rect 12012 58158 12014 58210
rect 12066 58158 12068 58210
rect 12012 58146 12068 58158
rect 11900 57540 11956 57550
rect 10780 56306 11060 56308
rect 10780 56254 10782 56306
rect 10834 56254 11060 56306
rect 10780 56252 11060 56254
rect 11228 56756 11284 56766
rect 11228 56306 11284 56700
rect 11228 56254 11230 56306
rect 11282 56254 11284 56306
rect 10780 56242 10836 56252
rect 11228 56242 11284 56254
rect 11564 56082 11620 56094
rect 11564 56030 11566 56082
rect 11618 56030 11620 56082
rect 11004 55524 11060 55534
rect 11564 55524 11620 56030
rect 11788 55524 11844 55534
rect 11564 55468 11788 55524
rect 11004 55298 11060 55468
rect 11788 55410 11844 55468
rect 11788 55358 11790 55410
rect 11842 55358 11844 55410
rect 11788 55346 11844 55358
rect 11004 55246 11006 55298
rect 11058 55246 11060 55298
rect 11004 55234 11060 55246
rect 11340 55300 11396 55310
rect 11340 55206 11396 55244
rect 11116 55074 11172 55086
rect 11116 55022 11118 55074
rect 11170 55022 11172 55074
rect 11004 54740 11060 54750
rect 11116 54740 11172 55022
rect 10668 54738 11172 54740
rect 10668 54686 11006 54738
rect 11058 54686 11172 54738
rect 10668 54684 11172 54686
rect 11004 54674 11060 54684
rect 10332 53566 10334 53618
rect 10386 53566 10388 53618
rect 10332 53554 10388 53566
rect 11340 54514 11396 54526
rect 11340 54462 11342 54514
rect 11394 54462 11396 54514
rect 10668 53508 10724 53518
rect 10668 53506 10836 53508
rect 10668 53454 10670 53506
rect 10722 53454 10836 53506
rect 10668 53452 10836 53454
rect 10668 53442 10724 53452
rect 9100 52946 9268 52948
rect 9100 52894 9102 52946
rect 9154 52894 9268 52946
rect 9100 52892 9268 52894
rect 9100 52882 9156 52892
rect 8764 52334 8766 52386
rect 8818 52334 8820 52386
rect 8764 52322 8820 52334
rect 8652 52110 8654 52162
rect 8706 52110 8708 52162
rect 8652 52098 8708 52110
rect 8764 52052 8820 52062
rect 8764 51958 8820 51996
rect 9100 50594 9156 50606
rect 9100 50542 9102 50594
rect 9154 50542 9156 50594
rect 8764 50484 8820 50494
rect 8540 50482 8820 50484
rect 8540 50430 8766 50482
rect 8818 50430 8820 50482
rect 8540 50428 8820 50430
rect 9100 50428 9156 50542
rect 8764 50418 8820 50428
rect 8988 50372 9156 50428
rect 8988 49924 9044 50372
rect 8652 49810 8708 49822
rect 8652 49758 8654 49810
rect 8706 49758 8708 49810
rect 7980 49700 8036 49710
rect 7980 49698 8372 49700
rect 7980 49646 7982 49698
rect 8034 49646 8372 49698
rect 7980 49644 8372 49646
rect 7980 49634 8036 49644
rect 8316 49028 8372 49644
rect 8652 49476 8708 49758
rect 8876 49812 8932 49822
rect 8876 49718 8932 49756
rect 8988 49476 9044 49868
rect 8652 49420 9044 49476
rect 8540 49140 8596 49150
rect 8540 49028 8596 49084
rect 8316 48972 8596 49028
rect 6748 48916 6804 48926
rect 6748 48822 6804 48860
rect 8428 48804 8484 48814
rect 8316 48468 8372 48478
rect 8316 48374 8372 48412
rect 8428 48466 8484 48748
rect 8428 48414 8430 48466
rect 8482 48414 8484 48466
rect 8428 48402 8484 48414
rect 8540 48466 8596 48972
rect 8540 48414 8542 48466
rect 8594 48414 8596 48466
rect 8540 48402 8596 48414
rect 8876 49138 8932 49150
rect 8876 49086 8878 49138
rect 8930 49086 8932 49138
rect 8092 48356 8148 48366
rect 8092 46228 8148 48300
rect 8876 48354 8932 49086
rect 8988 48466 9044 49420
rect 9100 49140 9156 49150
rect 9100 49026 9156 49084
rect 9100 48974 9102 49026
rect 9154 48974 9156 49026
rect 9100 48962 9156 48974
rect 8988 48414 8990 48466
rect 9042 48414 9044 48466
rect 8988 48402 9044 48414
rect 8876 48302 8878 48354
rect 8930 48302 8932 48354
rect 8876 48290 8932 48302
rect 9212 48356 9268 52892
rect 9772 52836 9828 52846
rect 9772 52834 9940 52836
rect 9772 52782 9774 52834
rect 9826 52782 9940 52834
rect 9772 52780 9940 52782
rect 9772 52770 9828 52780
rect 9324 50706 9380 50718
rect 9324 50654 9326 50706
rect 9378 50654 9380 50706
rect 9324 49812 9380 50654
rect 9772 50594 9828 50606
rect 9772 50542 9774 50594
rect 9826 50542 9828 50594
rect 9772 50148 9828 50542
rect 9884 50428 9940 52780
rect 10108 52834 10164 52846
rect 10108 52782 10110 52834
rect 10162 52782 10164 52834
rect 10108 52500 10164 52782
rect 10668 52836 10724 52846
rect 10780 52836 10836 53452
rect 11340 52948 11396 54462
rect 11564 52948 11620 52958
rect 11340 52946 11620 52948
rect 11340 52894 11566 52946
rect 11618 52894 11620 52946
rect 11340 52892 11620 52894
rect 11116 52836 11172 52846
rect 10780 52834 11172 52836
rect 10780 52782 11118 52834
rect 11170 52782 11172 52834
rect 10780 52780 11172 52782
rect 10668 52742 10724 52780
rect 10108 52434 10164 52444
rect 10220 52724 10276 52734
rect 10332 52724 10388 52734
rect 10276 52722 10388 52724
rect 10276 52670 10334 52722
rect 10386 52670 10388 52722
rect 10276 52668 10388 52670
rect 10220 52276 10276 52668
rect 10332 52658 10388 52668
rect 9996 52220 10276 52276
rect 9996 52050 10052 52220
rect 10332 52164 10388 52174
rect 10780 52164 10836 52174
rect 10332 52162 10780 52164
rect 10332 52110 10334 52162
rect 10386 52110 10780 52162
rect 10332 52108 10780 52110
rect 10332 52098 10388 52108
rect 10780 52070 10836 52108
rect 9996 51998 9998 52050
rect 10050 51998 10052 52050
rect 9996 51986 10052 51998
rect 10780 50482 10836 50494
rect 10780 50430 10782 50482
rect 10834 50430 10836 50482
rect 10780 50428 10836 50430
rect 11004 50428 11060 52780
rect 11116 52770 11172 52780
rect 11452 52500 11508 52510
rect 11452 52050 11508 52444
rect 11452 51998 11454 52050
rect 11506 51998 11508 52050
rect 11452 51986 11508 51998
rect 9884 50372 10164 50428
rect 9436 50092 9828 50148
rect 9436 50034 9492 50092
rect 9436 49982 9438 50034
rect 9490 49982 9492 50034
rect 9436 49970 9492 49982
rect 9660 49924 9716 49934
rect 9324 49746 9380 49756
rect 9548 49922 9716 49924
rect 9548 49870 9662 49922
rect 9714 49870 9716 49922
rect 9548 49868 9716 49870
rect 9324 48916 9380 48926
rect 9324 48822 9380 48860
rect 9548 48914 9604 49868
rect 9660 49858 9716 49868
rect 9772 49812 9828 49822
rect 9996 49812 10052 49822
rect 9772 49810 10052 49812
rect 9772 49758 9774 49810
rect 9826 49758 9998 49810
rect 10050 49758 10052 49810
rect 9772 49756 10052 49758
rect 9772 49746 9828 49756
rect 9996 49746 10052 49756
rect 10108 49140 10164 50372
rect 10444 50372 10836 50428
rect 10220 49924 10276 49934
rect 10220 49830 10276 49868
rect 10332 49812 10388 49822
rect 10332 49718 10388 49756
rect 10220 49140 10276 49150
rect 10108 49138 10276 49140
rect 10108 49086 10222 49138
rect 10274 49086 10276 49138
rect 10108 49084 10276 49086
rect 9548 48862 9550 48914
rect 9602 48862 9604 48914
rect 9212 48290 9268 48300
rect 9548 48468 9604 48862
rect 9660 49026 9716 49038
rect 9660 48974 9662 49026
rect 9714 48974 9716 49026
rect 9660 48804 9716 48974
rect 9660 48738 9716 48748
rect 10108 49028 10164 49084
rect 10220 49074 10276 49084
rect 9548 47684 9604 48412
rect 9548 47618 9604 47628
rect 9660 47460 9716 47470
rect 8876 46786 8932 46798
rect 8876 46734 8878 46786
rect 8930 46734 8932 46786
rect 8764 46674 8820 46686
rect 8764 46622 8766 46674
rect 8818 46622 8820 46674
rect 8092 46172 8372 46228
rect 8092 45892 8148 45902
rect 7756 45890 8148 45892
rect 7756 45838 8094 45890
rect 8146 45838 8148 45890
rect 7756 45836 8148 45838
rect 7532 45220 7588 45230
rect 6748 44996 6804 45006
rect 6748 44994 7364 44996
rect 6748 44942 6750 44994
rect 6802 44942 7364 44994
rect 6748 44940 7364 44942
rect 6748 44930 6804 44940
rect 7308 44434 7364 44940
rect 7308 44382 7310 44434
rect 7362 44382 7364 44434
rect 7308 44370 7364 44382
rect 7532 44322 7588 45164
rect 7532 44270 7534 44322
rect 7586 44270 7588 44322
rect 7532 44258 7588 44270
rect 7756 44322 7812 45836
rect 8092 45826 8148 45836
rect 7756 44270 7758 44322
rect 7810 44270 7812 44322
rect 7756 44258 7812 44270
rect 7980 45666 8036 45678
rect 7980 45614 7982 45666
rect 8034 45614 8036 45666
rect 7980 44436 8036 45614
rect 8204 45666 8260 45678
rect 8204 45614 8206 45666
rect 8258 45614 8260 45666
rect 8204 45220 8260 45614
rect 8204 45154 8260 45164
rect 8316 45668 8372 46172
rect 8764 45780 8820 46622
rect 8764 45714 8820 45724
rect 8428 45668 8484 45678
rect 8316 45666 8484 45668
rect 8316 45614 8430 45666
rect 8482 45614 8484 45666
rect 8316 45612 8484 45614
rect 8092 44436 8148 44446
rect 7980 44434 8148 44436
rect 7980 44382 8094 44434
rect 8146 44382 8148 44434
rect 7980 44380 8148 44382
rect 7196 44210 7252 44222
rect 7196 44158 7198 44210
rect 7250 44158 7252 44210
rect 7196 43988 7252 44158
rect 7980 43988 8036 44380
rect 8092 44370 8148 44380
rect 8316 44100 8372 45612
rect 8428 45602 8484 45612
rect 8876 45332 8932 46734
rect 9100 46674 9156 46686
rect 9100 46622 9102 46674
rect 9154 46622 9156 46674
rect 9100 46002 9156 46622
rect 9660 46114 9716 47404
rect 10108 46564 10164 48972
rect 10108 46562 10276 46564
rect 10108 46510 10110 46562
rect 10162 46510 10276 46562
rect 10108 46508 10276 46510
rect 10108 46498 10164 46508
rect 9660 46062 9662 46114
rect 9714 46062 9716 46114
rect 9660 46050 9716 46062
rect 9100 45950 9102 46002
rect 9154 45950 9156 46002
rect 9100 45938 9156 45950
rect 9996 46004 10052 46014
rect 9996 45910 10052 45948
rect 9324 45892 9380 45902
rect 9324 45890 9604 45892
rect 9324 45838 9326 45890
rect 9378 45838 9604 45890
rect 9324 45836 9604 45838
rect 9324 45826 9380 45836
rect 8876 44996 8932 45276
rect 8764 44994 8932 44996
rect 8764 44942 8878 44994
rect 8930 44942 8932 44994
rect 8764 44940 8932 44942
rect 8764 44322 8820 44940
rect 8876 44930 8932 44940
rect 9436 45444 9492 45454
rect 9436 45108 9492 45388
rect 9548 45332 9604 45836
rect 9996 45780 10052 45790
rect 9884 45724 9996 45780
rect 9660 45332 9716 45342
rect 9548 45330 9716 45332
rect 9548 45278 9662 45330
rect 9714 45278 9716 45330
rect 9548 45276 9716 45278
rect 9660 45266 9716 45276
rect 9772 45332 9828 45342
rect 9772 45238 9828 45276
rect 9324 44548 9380 44558
rect 8988 44546 9380 44548
rect 8988 44494 9326 44546
rect 9378 44494 9380 44546
rect 8988 44492 9380 44494
rect 8988 44434 9044 44492
rect 9324 44482 9380 44492
rect 8988 44382 8990 44434
rect 9042 44382 9044 44434
rect 8988 44370 9044 44382
rect 9436 44436 9492 45052
rect 9548 45108 9604 45118
rect 9884 45108 9940 45724
rect 9996 45714 10052 45724
rect 9548 45106 9940 45108
rect 9548 45054 9550 45106
rect 9602 45054 9940 45106
rect 9548 45052 9940 45054
rect 10108 45220 10164 45230
rect 10108 45106 10164 45164
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 9548 45042 9604 45052
rect 9660 44546 9716 45052
rect 9660 44494 9662 44546
rect 9714 44494 9716 44546
rect 9660 44482 9716 44494
rect 9548 44436 9604 44446
rect 9436 44434 9604 44436
rect 9436 44382 9550 44434
rect 9602 44382 9604 44434
rect 9436 44380 9604 44382
rect 9548 44370 9604 44380
rect 8764 44270 8766 44322
rect 8818 44270 8820 44322
rect 8764 44258 8820 44270
rect 7196 43932 8036 43988
rect 8092 44044 8372 44100
rect 8092 40626 8148 44044
rect 10108 42978 10164 45054
rect 10108 42926 10110 42978
rect 10162 42926 10164 42978
rect 10108 42914 10164 42926
rect 8428 42756 8484 42766
rect 8764 42756 8820 42766
rect 8428 42754 8764 42756
rect 8428 42702 8430 42754
rect 8482 42702 8764 42754
rect 8428 42700 8764 42702
rect 8428 42690 8484 42700
rect 8764 42662 8820 42700
rect 9660 42754 9716 42766
rect 9660 42702 9662 42754
rect 9714 42702 9716 42754
rect 8316 42644 8372 42654
rect 8204 41972 8260 41982
rect 8204 41858 8260 41916
rect 8204 41806 8206 41858
rect 8258 41806 8260 41858
rect 8204 41794 8260 41806
rect 8092 40574 8094 40626
rect 8146 40574 8148 40626
rect 8092 40562 8148 40574
rect 8204 41188 8260 41198
rect 7756 40404 7812 40414
rect 7084 40402 7812 40404
rect 7084 40350 7758 40402
rect 7810 40350 7812 40402
rect 7084 40348 7812 40350
rect 6860 39732 6916 39742
rect 6636 39730 6916 39732
rect 6636 39678 6862 39730
rect 6914 39678 6916 39730
rect 6636 39676 6916 39678
rect 5404 39666 5460 39676
rect 6188 39060 6244 39070
rect 6748 39060 6804 39676
rect 6860 39666 6916 39676
rect 6188 39058 6804 39060
rect 6188 39006 6190 39058
rect 6242 39006 6804 39058
rect 6188 39004 6804 39006
rect 6188 38994 6244 39004
rect 5852 38836 5908 38846
rect 4172 38612 4340 38668
rect 5068 38612 5236 38668
rect 3948 38274 4116 38276
rect 3948 38222 3950 38274
rect 4002 38222 4116 38274
rect 3948 38220 4116 38222
rect 4284 38276 4340 38612
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4284 38220 4564 38276
rect 3948 38210 4004 38220
rect 4060 38052 4116 38062
rect 3612 37996 4060 38052
rect 2716 37492 2772 37502
rect 2716 37378 2772 37436
rect 3612 37492 3668 37996
rect 4060 37958 4116 37996
rect 3612 37398 3668 37436
rect 3948 37826 4004 37838
rect 3948 37774 3950 37826
rect 4002 37774 4004 37826
rect 2716 37326 2718 37378
rect 2770 37326 2772 37378
rect 2716 37314 2772 37326
rect 3052 37380 3108 37390
rect 3052 37286 3108 37324
rect 3948 37380 4004 37774
rect 3164 37268 3220 37278
rect 3164 37174 3220 37212
rect 3724 37268 3780 37278
rect 3724 37174 3780 37212
rect 3836 37268 3892 37278
rect 3948 37268 4004 37324
rect 3836 37266 4004 37268
rect 3836 37214 3838 37266
rect 3890 37214 4004 37266
rect 3836 37212 4004 37214
rect 4284 37266 4340 38220
rect 4508 38162 4564 38220
rect 4508 38110 4510 38162
rect 4562 38110 4564 38162
rect 4508 38098 4564 38110
rect 4284 37214 4286 37266
rect 4338 37214 4340 37266
rect 2828 37154 2884 37166
rect 2828 37102 2830 37154
rect 2882 37102 2884 37154
rect 2828 36820 2884 37102
rect 2492 36764 2884 36820
rect 2492 36594 2548 36764
rect 2492 36542 2494 36594
rect 2546 36542 2548 36594
rect 2492 36530 2548 36542
rect 3836 36596 3892 37212
rect 4284 37202 4340 37214
rect 4620 37268 4676 37278
rect 4620 37174 4676 37212
rect 5180 37268 5236 38612
rect 5852 38050 5908 38780
rect 6412 38834 6468 38846
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6412 38612 6468 38782
rect 6636 38836 6692 38846
rect 6636 38742 6692 38780
rect 5852 37998 5854 38050
rect 5906 37998 5908 38050
rect 5852 37986 5908 37998
rect 6188 38556 6412 38612
rect 6188 38050 6244 38556
rect 6412 38546 6468 38556
rect 6524 38722 6580 38734
rect 6524 38670 6526 38722
rect 6578 38670 6580 38722
rect 6188 37998 6190 38050
rect 6242 37998 6244 38050
rect 6188 37986 6244 37998
rect 6412 38052 6468 38062
rect 6524 38052 6580 38670
rect 6748 38162 6804 39004
rect 7084 38834 7140 40348
rect 7756 40338 7812 40348
rect 7084 38782 7086 38834
rect 7138 38782 7140 38834
rect 7084 38500 7140 38782
rect 7868 39060 7924 39070
rect 7868 38946 7924 39004
rect 8204 39058 8260 41132
rect 8316 40962 8372 42588
rect 9100 42644 9156 42654
rect 9100 42550 9156 42588
rect 8988 42532 9044 42542
rect 8988 42438 9044 42476
rect 8876 42308 8932 42318
rect 8764 42082 8820 42094
rect 8764 42030 8766 42082
rect 8818 42030 8820 42082
rect 8764 41972 8820 42030
rect 8764 41906 8820 41916
rect 8876 41970 8932 42252
rect 9660 42308 9716 42702
rect 9660 42242 9716 42252
rect 10108 42754 10164 42766
rect 10108 42702 10110 42754
rect 10162 42702 10164 42754
rect 9884 42196 9940 42206
rect 9660 42082 9716 42094
rect 9660 42030 9662 42082
rect 9714 42030 9716 42082
rect 8876 41918 8878 41970
rect 8930 41918 8932 41970
rect 8876 41906 8932 41918
rect 9548 41970 9604 41982
rect 9548 41918 9550 41970
rect 9602 41918 9604 41970
rect 8988 41748 9044 41758
rect 9548 41748 9604 41918
rect 8988 41746 9604 41748
rect 8988 41694 8990 41746
rect 9042 41694 9604 41746
rect 8988 41692 9604 41694
rect 8988 41682 9044 41692
rect 9548 41300 9604 41692
rect 9548 41234 9604 41244
rect 9660 41972 9716 42030
rect 8652 41188 8708 41198
rect 8652 41094 8708 41132
rect 9660 41074 9716 41916
rect 9884 41970 9940 42140
rect 9884 41918 9886 41970
rect 9938 41918 9940 41970
rect 9884 41906 9940 41918
rect 9996 41300 10052 41310
rect 9996 41206 10052 41244
rect 10108 41188 10164 42702
rect 10220 41970 10276 46508
rect 10220 41918 10222 41970
rect 10274 41918 10276 41970
rect 10220 41906 10276 41918
rect 10108 41122 10164 41132
rect 9660 41022 9662 41074
rect 9714 41022 9716 41074
rect 9660 41010 9716 41022
rect 8316 40910 8318 40962
rect 8370 40910 8372 40962
rect 8316 40898 8372 40910
rect 8204 39006 8206 39058
rect 8258 39006 8260 39058
rect 8204 38994 8260 39006
rect 7868 38894 7870 38946
rect 7922 38894 7924 38946
rect 7868 38836 7924 38894
rect 7868 38770 7924 38780
rect 7980 38946 8036 38958
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7532 38724 7588 38762
rect 7532 38658 7588 38668
rect 7420 38612 7476 38622
rect 7140 38444 7252 38500
rect 7084 38434 7140 38444
rect 6748 38110 6750 38162
rect 6802 38110 6804 38162
rect 6748 38098 6804 38110
rect 6412 38050 6580 38052
rect 6412 37998 6414 38050
rect 6466 37998 6580 38050
rect 6412 37996 6580 37998
rect 7196 38050 7252 38444
rect 7196 37998 7198 38050
rect 7250 37998 7252 38050
rect 6412 37986 6468 37996
rect 7196 37986 7252 37998
rect 5964 37828 6020 37838
rect 5292 37826 6020 37828
rect 5292 37774 5966 37826
rect 6018 37774 6020 37826
rect 5292 37772 6020 37774
rect 5292 37378 5348 37772
rect 5964 37762 6020 37772
rect 5292 37326 5294 37378
rect 5346 37326 5348 37378
rect 5292 37314 5348 37326
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36596 4676 36606
rect 3836 36594 4676 36596
rect 3836 36542 4622 36594
rect 4674 36542 4676 36594
rect 3836 36540 4676 36542
rect 4620 36530 4676 36540
rect 5180 36594 5236 37212
rect 7420 37154 7476 38556
rect 7980 38612 8036 38894
rect 7980 38546 8036 38556
rect 9884 38276 9940 38286
rect 9884 38182 9940 38220
rect 8876 38050 8932 38062
rect 8876 37998 8878 38050
rect 8930 37998 8932 38050
rect 8764 37940 8820 37950
rect 8652 37938 8820 37940
rect 8652 37886 8766 37938
rect 8818 37886 8820 37938
rect 8652 37884 8820 37886
rect 8428 37380 8484 37390
rect 7868 37268 7924 37278
rect 7868 37174 7924 37212
rect 7420 37102 7422 37154
rect 7474 37102 7476 37154
rect 7420 37090 7476 37102
rect 5180 36542 5182 36594
rect 5234 36542 5236 36594
rect 5180 36530 5236 36542
rect 8428 36036 8484 37324
rect 8540 37378 8596 37390
rect 8540 37326 8542 37378
rect 8594 37326 8596 37378
rect 8540 37268 8596 37326
rect 8540 37202 8596 37212
rect 8652 37378 8708 37884
rect 8764 37874 8820 37884
rect 8652 37326 8654 37378
rect 8706 37326 8708 37378
rect 8652 36596 8708 37326
rect 8764 37380 8820 37390
rect 8764 37286 8820 37324
rect 8764 37156 8820 37166
rect 8764 37062 8820 37100
rect 8876 36706 8932 37998
rect 9548 38050 9604 38062
rect 9548 37998 9550 38050
rect 9602 37998 9604 38050
rect 8988 37268 9044 37278
rect 9324 37268 9380 37278
rect 8988 37266 9156 37268
rect 8988 37214 8990 37266
rect 9042 37214 9156 37266
rect 8988 37212 9156 37214
rect 8988 37202 9044 37212
rect 8876 36654 8878 36706
rect 8930 36654 8932 36706
rect 8876 36642 8932 36654
rect 9100 37044 9156 37212
rect 8764 36596 8820 36606
rect 8652 36540 8764 36596
rect 8764 36530 8820 36540
rect 8204 35980 8484 36036
rect 8764 36370 8820 36382
rect 8764 36318 8766 36370
rect 8818 36318 8820 36370
rect 2268 35588 2324 35598
rect 2268 35494 2324 35532
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 7868 34916 7924 34926
rect 7868 34822 7924 34860
rect 8204 34914 8260 35980
rect 8652 35700 8708 35710
rect 8652 35026 8708 35644
rect 8764 35364 8820 36318
rect 8764 35298 8820 35308
rect 8876 36372 8932 36382
rect 8876 36258 8932 36316
rect 8876 36206 8878 36258
rect 8930 36206 8932 36258
rect 8652 34974 8654 35026
rect 8706 34974 8708 35026
rect 8652 34962 8708 34974
rect 8204 34862 8206 34914
rect 8258 34862 8260 34914
rect 8204 34850 8260 34862
rect 8428 34916 8484 34926
rect 8484 34860 8596 34916
rect 8428 34822 8484 34860
rect 7980 34690 8036 34702
rect 7980 34638 7982 34690
rect 8034 34638 8036 34690
rect 5852 34020 5908 34030
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 2156 31892 2324 31948
rect 2268 26516 2324 31892
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4396 29428 4452 29438
rect 4396 29426 4900 29428
rect 4396 29374 4398 29426
rect 4450 29374 4900 29426
rect 4396 29372 4900 29374
rect 4396 29362 4452 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 27860 4900 29372
rect 5068 29316 5124 29326
rect 5068 29222 5124 29260
rect 5516 28420 5572 28430
rect 5516 27970 5572 28364
rect 5516 27918 5518 27970
rect 5570 27918 5572 27970
rect 5516 27906 5572 27918
rect 4844 27766 4900 27804
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2268 26450 2324 26460
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5852 11732 5908 33964
rect 7980 31892 8036 34638
rect 8540 34356 8596 34860
rect 8764 34802 8820 34814
rect 8764 34750 8766 34802
rect 8818 34750 8820 34802
rect 8540 34300 8708 34356
rect 7980 31826 8036 31836
rect 8540 34130 8596 34142
rect 8540 34078 8542 34130
rect 8594 34078 8596 34130
rect 8540 32676 8596 34078
rect 8540 31890 8596 32620
rect 8540 31838 8542 31890
rect 8594 31838 8596 31890
rect 8540 31826 8596 31838
rect 8652 31892 8708 34300
rect 8764 34244 8820 34750
rect 8764 34178 8820 34188
rect 8876 34018 8932 36206
rect 8876 33966 8878 34018
rect 8930 33966 8932 34018
rect 8876 33954 8932 33966
rect 8988 32788 9044 32798
rect 9100 32788 9156 36988
rect 9324 36594 9380 37212
rect 9436 37266 9492 37278
rect 9436 37214 9438 37266
rect 9490 37214 9492 37266
rect 9436 37156 9492 37214
rect 9436 37090 9492 37100
rect 9548 37044 9604 37998
rect 9884 37380 9940 37390
rect 9884 37286 9940 37324
rect 9548 36978 9604 36988
rect 10220 37266 10276 37278
rect 10220 37214 10222 37266
rect 10274 37214 10276 37266
rect 10220 37044 10276 37214
rect 10220 36978 10276 36988
rect 9324 36542 9326 36594
rect 9378 36542 9380 36594
rect 9324 36530 9380 36542
rect 9772 36596 9828 36606
rect 9436 35364 9492 35374
rect 9492 35308 9716 35364
rect 9436 35298 9492 35308
rect 9548 34916 9604 34926
rect 9548 33908 9604 34860
rect 9660 34354 9716 35308
rect 9660 34302 9662 34354
rect 9714 34302 9716 34354
rect 9660 34290 9716 34302
rect 9548 33906 9716 33908
rect 9548 33854 9550 33906
rect 9602 33854 9716 33906
rect 9548 33852 9716 33854
rect 9548 33842 9604 33852
rect 8988 32786 9156 32788
rect 8988 32734 8990 32786
rect 9042 32734 9156 32786
rect 8988 32732 9156 32734
rect 8988 32722 9044 32732
rect 8764 32562 8820 32574
rect 9548 32564 9604 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 32452 8820 32510
rect 8764 32386 8820 32396
rect 9324 32562 9604 32564
rect 9324 32510 9550 32562
rect 9602 32510 9604 32562
rect 9324 32508 9604 32510
rect 9324 32002 9380 32508
rect 9548 32498 9604 32508
rect 9324 31950 9326 32002
rect 9378 31950 9380 32002
rect 9324 31938 9380 31950
rect 8876 31892 8932 31902
rect 8652 31836 8820 31892
rect 8428 31778 8484 31790
rect 8428 31726 8430 31778
rect 8482 31726 8484 31778
rect 8092 31668 8148 31678
rect 7980 31612 8092 31668
rect 7644 30996 7700 31006
rect 7196 29316 7252 29326
rect 7644 29316 7700 30940
rect 7980 30100 8036 31612
rect 8092 31574 8148 31612
rect 8204 30882 8260 30894
rect 8204 30830 8206 30882
rect 8258 30830 8260 30882
rect 8204 30436 8260 30830
rect 8204 30370 8260 30380
rect 7196 29314 7700 29316
rect 7196 29262 7198 29314
rect 7250 29262 7700 29314
rect 7196 29260 7700 29262
rect 7868 30098 8036 30100
rect 7868 30046 7982 30098
rect 8034 30046 8036 30098
rect 7868 30044 8036 30046
rect 7868 29314 7924 30044
rect 7980 30034 8036 30044
rect 8092 30324 8148 30334
rect 7868 29262 7870 29314
rect 7922 29262 7924 29314
rect 7196 29250 7252 29260
rect 7868 29250 7924 29262
rect 8092 28754 8148 30268
rect 8428 30324 8484 31726
rect 8652 31666 8708 31678
rect 8652 31614 8654 31666
rect 8706 31614 8708 31666
rect 8540 30996 8596 31006
rect 8652 30996 8708 31614
rect 8596 30940 8708 30996
rect 8540 30902 8596 30940
rect 8428 30258 8484 30268
rect 8764 30100 8820 31836
rect 8876 30996 8932 31836
rect 8988 31668 9044 31678
rect 8988 31574 9044 31612
rect 9212 31556 9268 31566
rect 8876 30902 8932 30940
rect 9100 31554 9268 31556
rect 9100 31502 9214 31554
rect 9266 31502 9268 31554
rect 9100 31500 9268 31502
rect 8988 30436 9044 30446
rect 9100 30436 9156 31500
rect 9212 31490 9268 31500
rect 9044 30380 9156 30436
rect 9324 30772 9380 30782
rect 8988 30210 9044 30380
rect 9212 30324 9268 30334
rect 9212 30230 9268 30268
rect 8988 30158 8990 30210
rect 9042 30158 9044 30210
rect 8988 30146 9044 30158
rect 8540 30044 8820 30100
rect 8092 28702 8094 28754
rect 8146 28702 8148 28754
rect 8092 28690 8148 28702
rect 8316 29426 8372 29438
rect 8316 29374 8318 29426
rect 8370 29374 8372 29426
rect 7644 28642 7700 28654
rect 7644 28590 7646 28642
rect 7698 28590 7700 28642
rect 7196 28418 7252 28430
rect 7196 28366 7198 28418
rect 7250 28366 7252 28418
rect 6076 27860 6132 27870
rect 6076 26290 6132 27804
rect 7196 27860 7252 28366
rect 7196 27794 7252 27804
rect 7644 27748 7700 28590
rect 8316 28084 8372 29374
rect 8316 28018 8372 28028
rect 8092 27860 8148 27870
rect 8092 27766 8148 27804
rect 7644 27654 7700 27692
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 6076 26226 6132 26238
rect 8540 27188 8596 30044
rect 8988 29652 9044 29662
rect 8988 29538 9044 29596
rect 8988 29486 8990 29538
rect 9042 29486 9044 29538
rect 8988 29474 9044 29486
rect 8764 29426 8820 29438
rect 8764 29374 8766 29426
rect 8818 29374 8820 29426
rect 8652 27748 8708 27758
rect 8764 27748 8820 29374
rect 9324 28642 9380 30716
rect 9660 30100 9716 33852
rect 9772 33460 9828 36540
rect 9884 36258 9940 36270
rect 9884 36206 9886 36258
rect 9938 36206 9940 36258
rect 9884 36148 9940 36206
rect 9884 34132 9940 36092
rect 10444 35138 10500 50372
rect 10780 50036 10836 50372
rect 10780 49970 10836 49980
rect 10892 50372 11060 50428
rect 11116 50482 11172 50494
rect 11116 50430 11118 50482
rect 11170 50430 11172 50482
rect 10556 48356 10612 48366
rect 10556 46788 10612 48300
rect 10556 46004 10612 46732
rect 10556 45938 10612 45948
rect 10556 42754 10612 42766
rect 10556 42702 10558 42754
rect 10610 42702 10612 42754
rect 10556 42196 10612 42702
rect 10556 42130 10612 42140
rect 10780 38724 10836 38734
rect 10668 37940 10724 37950
rect 10556 37938 10724 37940
rect 10556 37886 10670 37938
rect 10722 37886 10724 37938
rect 10556 37884 10724 37886
rect 10556 37044 10612 37884
rect 10668 37874 10724 37884
rect 10780 37268 10836 38668
rect 10892 37380 10948 50372
rect 11116 50036 11172 50430
rect 11564 50428 11620 52892
rect 11788 51938 11844 51950
rect 11788 51886 11790 51938
rect 11842 51886 11844 51938
rect 11788 51604 11844 51886
rect 11788 51538 11844 51548
rect 11676 50708 11732 50718
rect 11676 50614 11732 50652
rect 11564 50372 11732 50428
rect 11116 49970 11172 49980
rect 11116 48914 11172 48926
rect 11116 48862 11118 48914
rect 11170 48862 11172 48914
rect 11116 48242 11172 48862
rect 11116 48190 11118 48242
rect 11170 48190 11172 48242
rect 11116 48132 11172 48190
rect 11116 48066 11172 48076
rect 11228 48802 11284 48814
rect 11228 48750 11230 48802
rect 11282 48750 11284 48802
rect 11116 47684 11172 47694
rect 11116 47590 11172 47628
rect 11228 47570 11284 48750
rect 11340 48802 11396 48814
rect 11340 48750 11342 48802
rect 11394 48750 11396 48802
rect 11340 48356 11396 48750
rect 11340 48290 11396 48300
rect 11228 47518 11230 47570
rect 11282 47518 11284 47570
rect 11228 47506 11284 47518
rect 11116 47460 11172 47470
rect 11116 47366 11172 47404
rect 11676 45332 11732 50372
rect 11788 48242 11844 48254
rect 11788 48190 11790 48242
rect 11842 48190 11844 48242
rect 11788 47460 11844 48190
rect 11788 47394 11844 47404
rect 11676 45266 11732 45276
rect 11788 47236 11844 47246
rect 11788 42756 11844 47180
rect 11900 43988 11956 57484
rect 12460 57540 12516 59948
rect 13804 59892 13860 60508
rect 13916 60004 13972 60622
rect 14140 60674 14308 60676
rect 14140 60622 14254 60674
rect 14306 60622 14308 60674
rect 14140 60620 14308 60622
rect 14140 60004 14196 60620
rect 14252 60610 14308 60620
rect 13916 59948 14140 60004
rect 14140 59910 14196 59948
rect 15148 60004 15204 60014
rect 13468 59890 13860 59892
rect 13468 59838 13806 59890
rect 13858 59838 13860 59890
rect 13468 59836 13860 59838
rect 12796 59780 12852 59790
rect 12796 59108 12852 59724
rect 12796 59014 12852 59052
rect 13468 58322 13524 59836
rect 13804 59826 13860 59836
rect 15036 59780 15092 59790
rect 15036 59442 15092 59724
rect 15036 59390 15038 59442
rect 15090 59390 15092 59442
rect 15036 59378 15092 59390
rect 15148 59442 15204 59948
rect 15148 59390 15150 59442
rect 15202 59390 15204 59442
rect 15148 59378 15204 59390
rect 15260 60002 15316 60014
rect 15260 59950 15262 60002
rect 15314 59950 15316 60002
rect 14476 59220 14532 59230
rect 14140 59218 14532 59220
rect 14140 59166 14478 59218
rect 14530 59166 14532 59218
rect 14140 59164 14532 59166
rect 13468 58270 13470 58322
rect 13522 58270 13524 58322
rect 13468 58258 13524 58270
rect 13804 58436 13860 58446
rect 13804 57874 13860 58380
rect 13804 57822 13806 57874
rect 13858 57822 13860 57874
rect 13804 57810 13860 57822
rect 13916 57650 13972 57662
rect 13916 57598 13918 57650
rect 13970 57598 13972 57650
rect 12460 57474 12516 57484
rect 13356 57540 13412 57550
rect 13356 57446 13412 57484
rect 13916 57540 13972 57598
rect 13916 57474 13972 57484
rect 13804 57426 13860 57438
rect 13804 57374 13806 57426
rect 13858 57374 13860 57426
rect 12236 57092 12292 57102
rect 12012 56756 12068 56766
rect 12012 56662 12068 56700
rect 12124 56308 12180 56318
rect 12236 56308 12292 57036
rect 13692 56756 13748 56766
rect 12572 56644 12628 56654
rect 12572 56550 12628 56588
rect 12124 56306 12292 56308
rect 12124 56254 12126 56306
rect 12178 56254 12292 56306
rect 12124 56252 12292 56254
rect 12908 56308 12964 56318
rect 12124 56242 12180 56252
rect 12908 56194 12964 56252
rect 13692 56306 13748 56700
rect 13804 56754 13860 57374
rect 14140 56978 14196 59164
rect 14476 59154 14532 59164
rect 14924 59218 14980 59230
rect 14924 59166 14926 59218
rect 14978 59166 14980 59218
rect 14140 56926 14142 56978
rect 14194 56926 14196 56978
rect 14140 56914 14196 56926
rect 14364 58884 14420 58894
rect 14364 58212 14420 58828
rect 14924 58436 14980 59166
rect 14476 58212 14532 58222
rect 14364 58210 14532 58212
rect 14364 58158 14478 58210
rect 14530 58158 14532 58210
rect 14364 58156 14532 58158
rect 13804 56702 13806 56754
rect 13858 56702 13860 56754
rect 13804 56690 13860 56702
rect 13916 56754 13972 56766
rect 13916 56702 13918 56754
rect 13970 56702 13972 56754
rect 13692 56254 13694 56306
rect 13746 56254 13748 56306
rect 13692 56242 13748 56254
rect 13916 56644 13972 56702
rect 14252 56756 14308 56766
rect 14252 56662 14308 56700
rect 12908 56142 12910 56194
rect 12962 56142 12964 56194
rect 12460 56084 12516 56094
rect 12796 56084 12852 56094
rect 12460 56082 12852 56084
rect 12460 56030 12462 56082
rect 12514 56030 12798 56082
rect 12850 56030 12852 56082
rect 12460 56028 12852 56030
rect 12460 56018 12516 56028
rect 12684 55076 12740 55086
rect 12796 55076 12852 56028
rect 12908 55524 12964 56142
rect 13132 56196 13188 56206
rect 13356 56196 13412 56206
rect 13132 56194 13356 56196
rect 13132 56142 13134 56194
rect 13186 56142 13356 56194
rect 13132 56140 13356 56142
rect 13132 56130 13188 56140
rect 13356 56102 13412 56140
rect 13468 56194 13524 56206
rect 13468 56142 13470 56194
rect 13522 56142 13524 56194
rect 13020 55524 13076 55534
rect 12908 55468 13020 55524
rect 12740 55020 12852 55076
rect 12684 54982 12740 55020
rect 12572 54516 12628 54526
rect 12572 53172 12628 54460
rect 12012 53116 12628 53172
rect 12012 53058 12068 53116
rect 12012 53006 12014 53058
rect 12066 53006 12068 53058
rect 12012 52994 12068 53006
rect 12572 53058 12628 53116
rect 12572 53006 12574 53058
rect 12626 53006 12628 53058
rect 12572 52994 12628 53006
rect 12908 53060 12964 53070
rect 12348 52946 12404 52958
rect 12348 52894 12350 52946
rect 12402 52894 12404 52946
rect 12348 52836 12404 52894
rect 12348 52770 12404 52780
rect 12684 52946 12740 52958
rect 12684 52894 12686 52946
rect 12738 52894 12740 52946
rect 12348 52276 12404 52286
rect 12684 52276 12740 52894
rect 12348 52274 12740 52276
rect 12348 52222 12350 52274
rect 12402 52222 12740 52274
rect 12348 52220 12740 52222
rect 12348 52210 12404 52220
rect 12796 52164 12852 52174
rect 12236 51938 12292 51950
rect 12236 51886 12238 51938
rect 12290 51886 12292 51938
rect 12236 50708 12292 51886
rect 12236 50642 12292 50652
rect 12460 51938 12516 51950
rect 12460 51886 12462 51938
rect 12514 51886 12516 51938
rect 12460 50428 12516 51886
rect 12796 51602 12852 52108
rect 12908 52164 12964 53004
rect 13020 52948 13076 55468
rect 13132 55412 13188 55422
rect 13132 53170 13188 55356
rect 13468 55300 13524 56142
rect 13916 56194 13972 56588
rect 14028 56644 14084 56654
rect 14028 56642 14196 56644
rect 14028 56590 14030 56642
rect 14082 56590 14196 56642
rect 14028 56588 14196 56590
rect 14028 56578 14084 56588
rect 13916 56142 13918 56194
rect 13970 56142 13972 56194
rect 13916 56130 13972 56142
rect 14028 56196 14084 56206
rect 14028 56102 14084 56140
rect 14028 55412 14084 55422
rect 14140 55412 14196 56588
rect 14252 56084 14308 56094
rect 14252 55990 14308 56028
rect 14084 55356 14196 55412
rect 14028 55346 14084 55356
rect 14364 55300 14420 58156
rect 14476 58146 14532 58156
rect 14924 57764 14980 58380
rect 15260 58212 15316 59950
rect 15596 60004 15652 61628
rect 16044 61628 16436 61684
rect 15708 60788 15764 60798
rect 15708 60114 15764 60732
rect 15708 60062 15710 60114
rect 15762 60062 15764 60114
rect 15708 60050 15764 60062
rect 15596 59938 15652 59948
rect 15708 59444 15764 59454
rect 16044 59444 16100 61628
rect 16268 60900 16324 60910
rect 16156 59892 16212 59902
rect 16156 59798 16212 59836
rect 16268 59892 16324 60844
rect 17500 60900 17556 60910
rect 17500 60806 17556 60844
rect 17948 60898 18004 62860
rect 18508 62914 18564 63084
rect 18508 62862 18510 62914
rect 18562 62862 18564 62914
rect 18172 62356 18228 62366
rect 17948 60846 17950 60898
rect 18002 60846 18004 60898
rect 17948 60834 18004 60846
rect 18060 60900 18116 60910
rect 18172 60900 18228 62300
rect 18060 60898 18228 60900
rect 18060 60846 18062 60898
rect 18114 60846 18228 60898
rect 18060 60844 18228 60846
rect 18060 60834 18116 60844
rect 17388 60786 17444 60798
rect 17388 60734 17390 60786
rect 17442 60734 17444 60786
rect 17052 60116 17108 60126
rect 17388 60116 17444 60734
rect 17724 60786 17780 60798
rect 17724 60734 17726 60786
rect 17778 60734 17780 60786
rect 17612 60228 17668 60238
rect 17612 60134 17668 60172
rect 17052 60114 17444 60116
rect 17052 60062 17054 60114
rect 17106 60062 17444 60114
rect 17052 60060 17444 60062
rect 16492 60004 16548 60014
rect 16940 60004 16996 60014
rect 16492 60002 16996 60004
rect 16492 59950 16494 60002
rect 16546 59950 16942 60002
rect 16994 59950 16996 60002
rect 16492 59948 16996 59950
rect 16492 59938 16548 59948
rect 16940 59938 16996 59948
rect 16268 59890 16436 59892
rect 16268 59838 16270 59890
rect 16322 59838 16436 59890
rect 16268 59836 16436 59838
rect 16268 59826 16324 59836
rect 15708 59442 16100 59444
rect 15708 59390 15710 59442
rect 15762 59390 16100 59442
rect 15708 59388 16100 59390
rect 16380 59444 16436 59836
rect 16940 59780 16996 59790
rect 17052 59780 17108 60060
rect 16996 59724 17108 59780
rect 16940 59714 16996 59724
rect 16716 59444 16772 59454
rect 16380 59388 16660 59444
rect 15708 59378 15764 59388
rect 15932 59220 15988 59230
rect 14924 57698 14980 57708
rect 15036 58156 15316 58212
rect 15372 58212 15428 58222
rect 15820 58212 15876 58222
rect 15932 58212 15988 59164
rect 16044 59218 16100 59230
rect 16044 59166 16046 59218
rect 16098 59166 16100 59218
rect 16044 58548 16100 59166
rect 16380 59220 16436 59230
rect 16380 59126 16436 59164
rect 16492 59108 16548 59118
rect 16044 58492 16324 58548
rect 16268 58436 16324 58492
rect 16380 58436 16436 58446
rect 16268 58380 16380 58436
rect 16380 58342 16436 58380
rect 16156 58322 16212 58334
rect 16156 58270 16158 58322
rect 16210 58270 16212 58322
rect 16156 58212 16212 58270
rect 15372 58210 16212 58212
rect 15372 58158 15374 58210
rect 15426 58158 15822 58210
rect 15874 58158 16212 58210
rect 15372 58156 16212 58158
rect 15036 56978 15092 58156
rect 15372 58146 15428 58156
rect 15036 56926 15038 56978
rect 15090 56926 15092 56978
rect 15036 56914 15092 56926
rect 15484 57764 15540 57774
rect 14588 56866 14644 56878
rect 14588 56814 14590 56866
rect 14642 56814 14644 56866
rect 14588 56644 14644 56814
rect 15148 56756 15204 56766
rect 15148 56662 15204 56700
rect 14588 56578 14644 56588
rect 14924 56642 14980 56654
rect 14924 56590 14926 56642
rect 14978 56590 14980 56642
rect 14588 56308 14644 56318
rect 14588 56214 14644 56252
rect 14924 55412 14980 56590
rect 15148 56084 15204 56094
rect 15148 55990 15204 56028
rect 15260 55970 15316 55982
rect 15260 55918 15262 55970
rect 15314 55918 15316 55970
rect 15260 55468 15316 55918
rect 14924 55346 14980 55356
rect 15036 55412 15316 55468
rect 13468 55234 13524 55244
rect 14140 55244 14420 55300
rect 14476 55300 14532 55310
rect 13132 53118 13134 53170
rect 13186 53118 13188 53170
rect 13132 53106 13188 53118
rect 13580 55076 13636 55086
rect 13020 52892 13188 52948
rect 12908 52162 13076 52164
rect 12908 52110 12910 52162
rect 12962 52110 13076 52162
rect 12908 52108 13076 52110
rect 12908 52098 12964 52108
rect 12796 51550 12798 51602
rect 12850 51550 12852 51602
rect 12460 50372 12740 50428
rect 12348 50036 12404 50046
rect 12348 49942 12404 49980
rect 12684 49812 12740 50372
rect 12684 49718 12740 49756
rect 12460 48130 12516 48142
rect 12460 48078 12462 48130
rect 12514 48078 12516 48130
rect 12124 47628 12404 47684
rect 12124 46002 12180 47628
rect 12236 47458 12292 47470
rect 12236 47406 12238 47458
rect 12290 47406 12292 47458
rect 12236 47348 12292 47406
rect 12348 47460 12404 47628
rect 12460 47682 12516 48078
rect 12460 47630 12462 47682
rect 12514 47630 12516 47682
rect 12460 47618 12516 47630
rect 12572 47460 12628 47470
rect 12348 47458 12628 47460
rect 12348 47406 12574 47458
rect 12626 47406 12628 47458
rect 12348 47404 12628 47406
rect 12572 47394 12628 47404
rect 12236 47292 12404 47348
rect 12348 47124 12404 47292
rect 12684 47236 12740 47246
rect 12684 47142 12740 47180
rect 12348 47068 12628 47124
rect 12348 46900 12404 46910
rect 12348 46674 12404 46844
rect 12572 46898 12628 47068
rect 12796 47012 12852 51550
rect 13020 51602 13076 52108
rect 13020 51550 13022 51602
rect 13074 51550 13076 51602
rect 13020 51538 13076 51550
rect 13132 51268 13188 52892
rect 13356 52164 13412 52174
rect 13244 51604 13300 51614
rect 13244 51510 13300 51548
rect 13356 51378 13412 52108
rect 13356 51326 13358 51378
rect 13410 51326 13412 51378
rect 13356 51314 13412 51326
rect 13468 51604 13524 51614
rect 13132 51212 13300 51268
rect 13244 50428 13300 51212
rect 13244 50372 13412 50428
rect 13244 49812 13300 49822
rect 13244 49718 13300 49756
rect 12572 46846 12574 46898
rect 12626 46846 12628 46898
rect 12572 46834 12628 46846
rect 12684 46956 12852 47012
rect 12908 48132 12964 48142
rect 12348 46622 12350 46674
rect 12402 46622 12404 46674
rect 12348 46610 12404 46622
rect 12124 45950 12126 46002
rect 12178 45950 12180 46002
rect 12124 45938 12180 45950
rect 12684 44660 12740 46956
rect 12796 46788 12852 46798
rect 12796 46694 12852 46732
rect 12908 46786 12964 48076
rect 13020 48130 13076 48142
rect 13020 48078 13022 48130
rect 13074 48078 13076 48130
rect 13020 47236 13076 48078
rect 13020 47170 13076 47180
rect 13356 47124 13412 50372
rect 12908 46734 12910 46786
rect 12962 46734 12964 46786
rect 12908 46722 12964 46734
rect 13244 47068 13412 47124
rect 12796 45890 12852 45902
rect 12796 45838 12798 45890
rect 12850 45838 12852 45890
rect 12796 45444 12852 45838
rect 12796 45378 12852 45388
rect 12236 44604 12740 44660
rect 12124 43988 12180 43998
rect 11900 43932 12124 43988
rect 12124 43922 12180 43932
rect 11788 42690 11844 42700
rect 11564 42084 11620 42094
rect 11564 42082 11844 42084
rect 11564 42030 11566 42082
rect 11618 42030 11844 42082
rect 11564 42028 11844 42030
rect 11564 42018 11620 42028
rect 11004 41858 11060 41870
rect 11004 41806 11006 41858
rect 11058 41806 11060 41858
rect 11004 41076 11060 41806
rect 11788 41300 11844 42028
rect 11788 41188 11844 41244
rect 12124 41188 12180 41198
rect 11788 41186 12180 41188
rect 11788 41134 12126 41186
rect 12178 41134 12180 41186
rect 11788 41132 12180 41134
rect 12124 41122 12180 41132
rect 11004 40404 11060 41020
rect 12236 40964 12292 44604
rect 12572 44100 12628 44110
rect 12348 41076 12404 41086
rect 12348 40982 12404 41020
rect 12460 41074 12516 41086
rect 12460 41022 12462 41074
rect 12514 41022 12516 41074
rect 11004 40338 11060 40348
rect 11900 40908 12292 40964
rect 12460 40964 12516 41022
rect 11452 39618 11508 39630
rect 11452 39566 11454 39618
rect 11506 39566 11508 39618
rect 11452 38836 11508 39566
rect 11452 38742 11508 38780
rect 11676 39394 11732 39406
rect 11676 39342 11678 39394
rect 11730 39342 11732 39394
rect 11676 38724 11732 39342
rect 11676 38658 11732 38668
rect 11116 38610 11172 38622
rect 11116 38558 11118 38610
rect 11170 38558 11172 38610
rect 11116 38052 11172 38558
rect 11788 38388 11844 38398
rect 11788 38274 11844 38332
rect 11788 38222 11790 38274
rect 11842 38222 11844 38274
rect 11788 38210 11844 38222
rect 11900 38276 11956 40908
rect 12460 40898 12516 40908
rect 12572 40628 12628 44044
rect 12124 40572 12628 40628
rect 12684 43988 12740 43998
rect 12012 38948 12068 38958
rect 12012 38854 12068 38892
rect 11900 38210 11956 38220
rect 11116 37986 11172 37996
rect 11452 38052 11508 38062
rect 11452 38050 11732 38052
rect 11452 37998 11454 38050
rect 11506 37998 11732 38050
rect 11452 37996 11732 37998
rect 11452 37986 11508 37996
rect 11228 37938 11284 37950
rect 11228 37886 11230 37938
rect 11282 37886 11284 37938
rect 11228 37380 11284 37886
rect 11340 37380 11396 37390
rect 11228 37324 11340 37380
rect 10892 37314 10948 37324
rect 11340 37286 11396 37324
rect 10556 36978 10612 36988
rect 10668 37212 10836 37268
rect 10668 35252 10724 37212
rect 11004 37044 11060 37054
rect 11004 36484 11060 36988
rect 11116 37044 11172 37054
rect 11116 37042 11284 37044
rect 11116 36990 11118 37042
rect 11170 36990 11284 37042
rect 11116 36988 11284 36990
rect 11116 36978 11172 36988
rect 11116 36484 11172 36494
rect 11004 36482 11172 36484
rect 11004 36430 11118 36482
rect 11170 36430 11172 36482
rect 11004 36428 11172 36430
rect 11228 36484 11284 36988
rect 11452 36484 11508 36494
rect 11228 36482 11508 36484
rect 11228 36430 11454 36482
rect 11506 36430 11508 36482
rect 11228 36428 11508 36430
rect 10780 36260 10836 36270
rect 10780 36166 10836 36204
rect 11004 36258 11060 36270
rect 11004 36206 11006 36258
rect 11058 36206 11060 36258
rect 11004 36148 11060 36206
rect 11004 36082 11060 36092
rect 10668 35196 10948 35252
rect 10444 35086 10446 35138
rect 10498 35086 10500 35138
rect 10444 35074 10500 35086
rect 9996 34916 10052 34926
rect 9996 34822 10052 34860
rect 10556 34914 10612 34926
rect 10556 34862 10558 34914
rect 10610 34862 10612 34914
rect 10556 34692 10612 34862
rect 10892 34916 10948 35196
rect 11116 34916 11172 36428
rect 11340 35700 11396 36428
rect 11452 36418 11508 36428
rect 11564 36372 11620 36382
rect 11564 35700 11620 36316
rect 11676 35922 11732 37996
rect 12012 37378 12068 37390
rect 12012 37326 12014 37378
rect 12066 37326 12068 37378
rect 11900 37266 11956 37278
rect 11900 37214 11902 37266
rect 11954 37214 11956 37266
rect 11900 37044 11956 37214
rect 11900 36978 11956 36988
rect 12012 36820 12068 37326
rect 11900 36764 12068 36820
rect 11900 36372 11956 36764
rect 12012 36596 12068 36606
rect 12124 36596 12180 40572
rect 12348 39620 12404 39630
rect 12236 39618 12404 39620
rect 12236 39566 12350 39618
rect 12402 39566 12404 39618
rect 12236 39564 12404 39566
rect 12236 38946 12292 39564
rect 12348 39554 12404 39564
rect 12572 39396 12628 39406
rect 12572 39302 12628 39340
rect 12236 38894 12238 38946
rect 12290 38894 12292 38946
rect 12236 38612 12292 38894
rect 12236 38546 12292 38556
rect 12348 39060 12404 39070
rect 12236 38276 12292 38286
rect 12348 38276 12404 39004
rect 12460 38834 12516 38846
rect 12460 38782 12462 38834
rect 12514 38782 12516 38834
rect 12460 38724 12516 38782
rect 12572 38836 12628 38874
rect 12572 38770 12628 38780
rect 12460 38658 12516 38668
rect 12236 38274 12404 38276
rect 12236 38222 12238 38274
rect 12290 38222 12404 38274
rect 12236 38220 12404 38222
rect 12572 38612 12628 38622
rect 12572 38274 12628 38556
rect 12572 38222 12574 38274
rect 12626 38222 12628 38274
rect 12236 38210 12292 38220
rect 12572 38210 12628 38222
rect 12684 37490 12740 43932
rect 13020 43092 13076 43102
rect 13020 42868 13076 43036
rect 12796 42866 13076 42868
rect 12796 42814 13022 42866
rect 13074 42814 13076 42866
rect 12796 42812 13076 42814
rect 12796 41970 12852 42812
rect 13020 42802 13076 42812
rect 12796 41918 12798 41970
rect 12850 41918 12852 41970
rect 12796 40628 12852 41918
rect 12852 40572 13076 40628
rect 12796 40562 12852 40572
rect 12908 39620 12964 39630
rect 12908 39506 12964 39564
rect 12908 39454 12910 39506
rect 12962 39454 12964 39506
rect 12908 38948 12964 39454
rect 13020 39058 13076 40572
rect 13020 39006 13022 39058
rect 13074 39006 13076 39058
rect 13020 38994 13076 39006
rect 12908 38668 12964 38892
rect 13132 38836 13188 38846
rect 13132 38668 13188 38780
rect 12796 38612 12964 38668
rect 13020 38612 13188 38668
rect 12796 38162 12852 38612
rect 12796 38110 12798 38162
rect 12850 38110 12852 38162
rect 12796 38098 12852 38110
rect 12684 37438 12686 37490
rect 12738 37438 12740 37490
rect 12684 37426 12740 37438
rect 12460 37380 12516 37390
rect 12460 37286 12516 37324
rect 12012 36594 12180 36596
rect 12012 36542 12014 36594
rect 12066 36542 12180 36594
rect 12012 36540 12180 36542
rect 12012 36530 12068 36540
rect 12348 36484 12404 36494
rect 11900 36306 11956 36316
rect 12124 36482 12404 36484
rect 12124 36430 12350 36482
rect 12402 36430 12404 36482
rect 12124 36428 12404 36430
rect 11676 35870 11678 35922
rect 11730 35870 11732 35922
rect 11676 35858 11732 35870
rect 11676 35700 11732 35710
rect 11564 35698 11732 35700
rect 11564 35646 11678 35698
rect 11730 35646 11732 35698
rect 11564 35644 11732 35646
rect 11340 35606 11396 35644
rect 11676 35634 11732 35644
rect 12012 35698 12068 35710
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 11452 34916 11508 34926
rect 10892 34914 11060 34916
rect 10892 34862 10894 34914
rect 10946 34862 11060 34914
rect 10892 34860 11060 34862
rect 10892 34850 10948 34860
rect 10556 34626 10612 34636
rect 9884 34038 9940 34076
rect 10556 34242 10612 34254
rect 10556 34190 10558 34242
rect 10610 34190 10612 34242
rect 10556 33684 10612 34190
rect 10556 33618 10612 33628
rect 10780 34244 10836 34254
rect 9772 33404 10052 33460
rect 9884 32452 9940 32462
rect 9772 31668 9828 31678
rect 9772 30882 9828 31612
rect 9884 31218 9940 32396
rect 9884 31166 9886 31218
rect 9938 31166 9940 31218
rect 9884 31154 9940 31166
rect 9772 30830 9774 30882
rect 9826 30830 9828 30882
rect 9772 30818 9828 30830
rect 9884 30994 9940 31006
rect 9884 30942 9886 30994
rect 9938 30942 9940 30994
rect 9772 30324 9828 30334
rect 9884 30324 9940 30942
rect 9828 30268 9940 30324
rect 9772 30258 9828 30268
rect 9772 30100 9828 30110
rect 9660 30098 9828 30100
rect 9660 30046 9774 30098
rect 9826 30046 9828 30098
rect 9660 30044 9828 30046
rect 9772 30034 9828 30044
rect 9996 29428 10052 33404
rect 10780 32676 10836 34188
rect 10444 32620 10836 32676
rect 10892 33348 10948 33358
rect 10332 31890 10388 31902
rect 10332 31838 10334 31890
rect 10386 31838 10388 31890
rect 10220 30994 10276 31006
rect 10220 30942 10222 30994
rect 10274 30942 10276 30994
rect 10220 30884 10276 30942
rect 10220 30818 10276 30828
rect 10332 29652 10388 31838
rect 10444 31778 10500 32620
rect 10892 32564 10948 33292
rect 11004 32674 11060 34860
rect 11116 34354 11172 34860
rect 11116 34302 11118 34354
rect 11170 34302 11172 34354
rect 11116 34290 11172 34302
rect 11340 34914 11508 34916
rect 11340 34862 11454 34914
rect 11506 34862 11508 34914
rect 11340 34860 11508 34862
rect 12012 34916 12068 35646
rect 12124 35140 12180 36428
rect 12348 36418 12404 36428
rect 12684 36260 12740 36270
rect 12684 36166 12740 36204
rect 13020 35924 13076 38612
rect 13244 38388 13300 47068
rect 13356 46900 13412 46910
rect 13356 46806 13412 46844
rect 13468 44548 13524 51548
rect 13580 46228 13636 55020
rect 13692 52834 13748 52846
rect 13692 52782 13694 52834
rect 13746 52782 13748 52834
rect 13692 52274 13748 52782
rect 13692 52222 13694 52274
rect 13746 52222 13748 52274
rect 13692 52164 13748 52222
rect 13692 52098 13748 52108
rect 13804 52162 13860 52174
rect 13804 52110 13806 52162
rect 13858 52110 13860 52162
rect 13804 51604 13860 52110
rect 13804 51538 13860 51548
rect 14028 50594 14084 50606
rect 14028 50542 14030 50594
rect 14082 50542 14084 50594
rect 13692 50372 13748 50382
rect 14028 50372 14084 50542
rect 14140 50596 14196 55244
rect 14476 55206 14532 55244
rect 14588 55076 14644 55086
rect 14252 55074 14644 55076
rect 14252 55022 14590 55074
rect 14642 55022 14644 55074
rect 14252 55020 14644 55022
rect 14252 54514 14308 55020
rect 14588 55010 14644 55020
rect 15036 54852 15092 55412
rect 14700 54796 15092 54852
rect 14588 54740 14644 54750
rect 14700 54740 14756 54796
rect 14588 54738 14756 54740
rect 14588 54686 14590 54738
rect 14642 54686 14756 54738
rect 14588 54684 14756 54686
rect 14588 54674 14644 54684
rect 14252 54462 14254 54514
rect 14306 54462 14308 54514
rect 14252 54450 14308 54462
rect 14476 54516 14532 54526
rect 14812 54516 14868 54526
rect 15148 54516 15204 54526
rect 14476 54422 14532 54460
rect 14700 54514 15204 54516
rect 14700 54462 14814 54514
rect 14866 54462 15150 54514
rect 15202 54462 15204 54514
rect 14700 54460 15204 54462
rect 14588 53172 14644 53182
rect 14700 53172 14756 54460
rect 14812 54450 14868 54460
rect 15148 54450 15204 54460
rect 15372 54516 15428 54526
rect 15372 54422 15428 54460
rect 14588 53170 14756 53172
rect 14588 53118 14590 53170
rect 14642 53118 14756 53170
rect 14588 53116 14756 53118
rect 14588 53106 14644 53116
rect 14812 53060 14868 53070
rect 14812 52966 14868 53004
rect 14924 52946 14980 52958
rect 14924 52894 14926 52946
rect 14978 52894 14980 52946
rect 14924 52276 14980 52894
rect 14476 52164 14532 52174
rect 14476 51380 14532 52108
rect 14812 52162 14868 52174
rect 14812 52110 14814 52162
rect 14866 52110 14868 52162
rect 14588 51380 14644 51390
rect 14476 51378 14644 51380
rect 14476 51326 14590 51378
rect 14642 51326 14644 51378
rect 14476 51324 14644 51326
rect 14588 51314 14644 51324
rect 14364 50820 14420 50830
rect 14812 50820 14868 52110
rect 14924 51716 14980 52220
rect 15036 52162 15092 52174
rect 15036 52110 15038 52162
rect 15090 52110 15092 52162
rect 15036 51828 15092 52110
rect 15260 52164 15316 52174
rect 15260 52070 15316 52108
rect 15036 51772 15316 51828
rect 14924 51660 15204 51716
rect 15148 51602 15204 51660
rect 15148 51550 15150 51602
rect 15202 51550 15204 51602
rect 15148 51538 15204 51550
rect 15036 51378 15092 51390
rect 15036 51326 15038 51378
rect 15090 51326 15092 51378
rect 15036 50820 15092 51326
rect 14364 50818 15092 50820
rect 14364 50766 14366 50818
rect 14418 50766 15092 50818
rect 14364 50764 15092 50766
rect 15260 51378 15316 51772
rect 15260 51326 15262 51378
rect 15314 51326 15316 51378
rect 14364 50754 14420 50764
rect 14140 50540 14420 50596
rect 14364 50428 14420 50540
rect 13692 50370 14084 50372
rect 13692 50318 13694 50370
rect 13746 50318 14084 50370
rect 13692 50316 14084 50318
rect 13692 50306 13748 50316
rect 14028 50036 14084 50316
rect 14028 49698 14084 49980
rect 14028 49646 14030 49698
rect 14082 49646 14084 49698
rect 14028 49634 14084 49646
rect 14252 50370 14308 50382
rect 14364 50372 14868 50428
rect 14252 50318 14254 50370
rect 14306 50318 14308 50370
rect 14252 49812 14308 50318
rect 13916 48356 13972 48366
rect 13692 48354 13972 48356
rect 13692 48302 13918 48354
rect 13970 48302 13972 48354
rect 13692 48300 13972 48302
rect 13692 47012 13748 48300
rect 13916 48290 13972 48300
rect 14028 48244 14084 48254
rect 14028 48150 14084 48188
rect 13804 48132 13860 48142
rect 13804 47346 13860 48076
rect 14140 48132 14196 48142
rect 14140 48038 14196 48076
rect 14252 47460 14308 49756
rect 14700 49588 14756 49598
rect 14700 49494 14756 49532
rect 14028 47404 14308 47460
rect 14588 48354 14644 48366
rect 14588 48302 14590 48354
rect 14642 48302 14644 48354
rect 14028 47348 14084 47404
rect 13804 47294 13806 47346
rect 13858 47294 13860 47346
rect 13804 47282 13860 47294
rect 13916 47292 14084 47348
rect 13692 46898 13748 46956
rect 13692 46846 13694 46898
rect 13746 46846 13748 46898
rect 13692 46834 13748 46846
rect 13580 46172 13748 46228
rect 13580 46004 13636 46014
rect 13580 45666 13636 45948
rect 13580 45614 13582 45666
rect 13634 45614 13636 45666
rect 13580 45444 13636 45614
rect 13580 45378 13636 45388
rect 13468 44492 13636 44548
rect 13468 44324 13524 44334
rect 13468 44210 13524 44268
rect 13468 44158 13470 44210
rect 13522 44158 13524 44210
rect 13468 44146 13524 44158
rect 13244 38322 13300 38332
rect 13468 41972 13524 41982
rect 13468 41074 13524 41916
rect 13468 41022 13470 41074
rect 13522 41022 13524 41074
rect 12796 35868 13076 35924
rect 12124 35138 12628 35140
rect 12124 35086 12126 35138
rect 12178 35086 12628 35138
rect 12124 35084 12628 35086
rect 12124 35074 12180 35084
rect 12012 34860 12292 34916
rect 11004 32622 11006 32674
rect 11058 32622 11060 32674
rect 11004 32610 11060 32622
rect 11340 34130 11396 34860
rect 11452 34850 11508 34860
rect 11340 34078 11342 34130
rect 11394 34078 11396 34130
rect 10780 32562 10948 32564
rect 10780 32510 10894 32562
rect 10946 32510 10948 32562
rect 10780 32508 10948 32510
rect 10780 32002 10836 32508
rect 10892 32498 10948 32508
rect 10780 31950 10782 32002
rect 10834 31950 10836 32002
rect 10780 31938 10836 31950
rect 11340 31780 11396 34078
rect 10444 31726 10446 31778
rect 10498 31726 10500 31778
rect 10444 30772 10500 31726
rect 10444 30706 10500 30716
rect 10556 31778 11396 31780
rect 10556 31726 11342 31778
rect 11394 31726 11396 31778
rect 10556 31724 11396 31726
rect 10332 29428 10388 29596
rect 10332 29372 10500 29428
rect 9996 28754 10052 29372
rect 10444 29314 10500 29372
rect 10444 29262 10446 29314
rect 10498 29262 10500 29314
rect 10444 29250 10500 29262
rect 9996 28702 9998 28754
rect 10050 28702 10052 28754
rect 9996 28690 10052 28702
rect 9324 28590 9326 28642
rect 9378 28590 9380 28642
rect 9324 28578 9380 28590
rect 10444 28532 10500 28542
rect 10556 28532 10612 31724
rect 11340 31714 11396 31724
rect 11452 34692 11508 34702
rect 11452 32562 11508 34636
rect 11788 34690 11844 34702
rect 11788 34638 11790 34690
rect 11842 34638 11844 34690
rect 11788 34356 11844 34638
rect 11676 34300 11844 34356
rect 12012 34690 12068 34702
rect 12012 34638 12014 34690
rect 12066 34638 12068 34690
rect 11676 33908 11732 34300
rect 11788 34130 11844 34142
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 11788 34020 11844 34078
rect 11788 33964 11956 34020
rect 11676 33852 11844 33908
rect 11676 33348 11732 33358
rect 11676 33254 11732 33292
rect 11452 32510 11454 32562
rect 11506 32510 11508 32562
rect 11452 31556 11508 32510
rect 11228 31500 11508 31556
rect 11116 30882 11172 30894
rect 11116 30830 11118 30882
rect 11170 30830 11172 30882
rect 11116 30772 11172 30830
rect 11116 30706 11172 30716
rect 11004 30436 11060 30446
rect 10444 28530 10612 28532
rect 10444 28478 10446 28530
rect 10498 28478 10612 28530
rect 10444 28476 10612 28478
rect 10668 29764 10724 29774
rect 10444 27970 10500 28476
rect 10444 27918 10446 27970
rect 10498 27918 10500 27970
rect 10444 27906 10500 27918
rect 8708 27692 8820 27748
rect 9548 27858 9604 27870
rect 9548 27806 9550 27858
rect 9602 27806 9604 27858
rect 9548 27748 9604 27806
rect 8652 27682 8708 27692
rect 9548 27682 9604 27692
rect 9660 27860 9716 27870
rect 9660 27188 9716 27804
rect 9996 27748 10052 27758
rect 9996 27654 10052 27692
rect 8540 27132 9268 27188
rect 6748 26180 6804 26190
rect 6748 26178 8372 26180
rect 6748 26126 6750 26178
rect 6802 26126 8372 26178
rect 6748 26124 8372 26126
rect 6748 26114 6804 26124
rect 8316 25618 8372 26124
rect 8316 25566 8318 25618
rect 8370 25566 8372 25618
rect 8316 25554 8372 25566
rect 8540 25506 8596 27132
rect 9212 26962 9268 27132
rect 9660 27186 10052 27188
rect 9660 27134 9662 27186
rect 9714 27134 10052 27186
rect 9660 27132 10052 27134
rect 9660 27122 9716 27132
rect 8876 26908 8932 26918
rect 9212 26910 9214 26962
rect 9266 26910 9268 26962
rect 9212 26908 9268 26910
rect 9212 26852 9828 26908
rect 8876 26850 8932 26852
rect 8876 26798 8878 26850
rect 8930 26798 8932 26850
rect 8876 26178 8932 26798
rect 9772 26514 9828 26852
rect 9772 26462 9774 26514
rect 9826 26462 9828 26514
rect 9772 26450 9828 26462
rect 9548 26290 9604 26302
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 8876 26126 8878 26178
rect 8930 26126 8932 26178
rect 8876 26114 8932 26126
rect 8988 26180 9044 26190
rect 8876 25956 8932 25966
rect 8540 25454 8542 25506
rect 8594 25454 8596 25506
rect 8540 25442 8596 25454
rect 8764 25900 8876 25956
rect 8764 25506 8820 25900
rect 8876 25890 8932 25900
rect 8764 25454 8766 25506
rect 8818 25454 8820 25506
rect 8764 25442 8820 25454
rect 8204 25396 8260 25406
rect 8204 25302 8260 25340
rect 8988 25396 9044 26124
rect 9548 26180 9604 26238
rect 9548 26114 9604 26124
rect 9660 26178 9716 26190
rect 9660 26126 9662 26178
rect 9714 26126 9716 26178
rect 9660 25956 9716 26126
rect 9660 25890 9716 25900
rect 9436 25620 9492 25630
rect 9436 25526 9492 25564
rect 8988 24946 9044 25340
rect 9996 25508 10052 27132
rect 10668 26516 10724 29708
rect 11004 28642 11060 30380
rect 11116 30324 11172 30334
rect 11116 30230 11172 30268
rect 11228 29426 11284 31500
rect 11452 30994 11508 31006
rect 11452 30942 11454 30994
rect 11506 30942 11508 30994
rect 11452 30884 11508 30942
rect 11788 30996 11844 33852
rect 11900 32228 11956 33964
rect 12012 33684 12068 34638
rect 12012 33618 12068 33628
rect 12236 34130 12292 34860
rect 12572 34914 12628 35084
rect 12572 34862 12574 34914
rect 12626 34862 12628 34914
rect 12572 34850 12628 34862
rect 12684 34692 12740 34702
rect 12684 34598 12740 34636
rect 12236 34078 12238 34130
rect 12290 34078 12292 34130
rect 12236 33346 12292 34078
rect 12796 33570 12852 35868
rect 13468 35140 13524 41022
rect 13580 38668 13636 44492
rect 13692 41300 13748 46172
rect 13916 45556 13972 47292
rect 14140 47236 14196 47246
rect 14588 47236 14644 48302
rect 14700 47236 14756 47246
rect 14140 47234 14420 47236
rect 14140 47182 14142 47234
rect 14194 47182 14420 47234
rect 14140 47180 14420 47182
rect 14140 47170 14196 47180
rect 14028 46676 14084 46686
rect 14252 46676 14308 46686
rect 14028 46674 14252 46676
rect 14028 46622 14030 46674
rect 14082 46622 14252 46674
rect 14028 46620 14252 46622
rect 14028 46610 14084 46620
rect 14252 46610 14308 46620
rect 14364 46564 14420 47180
rect 14588 47234 14756 47236
rect 14588 47182 14702 47234
rect 14754 47182 14756 47234
rect 14588 47180 14756 47182
rect 14476 46564 14532 46574
rect 14364 46508 14476 46564
rect 14476 46498 14532 46508
rect 14588 46340 14644 47180
rect 14700 47170 14756 47180
rect 14812 46900 14868 50372
rect 15260 48354 15316 51326
rect 15484 49812 15540 57708
rect 15596 49924 15652 58156
rect 15820 58146 15876 58156
rect 16156 56980 16212 56990
rect 16492 56980 16548 59052
rect 16604 58660 16660 59388
rect 16716 59350 16772 59388
rect 17612 59332 17668 59342
rect 17612 59238 17668 59276
rect 17724 59218 17780 60734
rect 18060 60562 18116 60574
rect 18060 60510 18062 60562
rect 18114 60510 18116 60562
rect 18060 59892 18116 60510
rect 18060 59332 18116 59836
rect 18172 60116 18228 60844
rect 18172 59444 18228 60060
rect 18508 59780 18564 62862
rect 19404 63138 19684 63140
rect 19404 63086 19630 63138
rect 19682 63086 19684 63138
rect 19404 63084 19684 63086
rect 19404 62578 19460 63084
rect 19628 63074 19684 63084
rect 19964 63026 20020 63038
rect 19964 62974 19966 63026
rect 20018 62974 20020 63026
rect 19964 62916 20020 62974
rect 19404 62526 19406 62578
rect 19458 62526 19460 62578
rect 19404 62514 19460 62526
rect 19628 62860 20020 62916
rect 19628 62580 19684 62860
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 20860 62692 20916 63758
rect 20972 63140 21028 63980
rect 21084 63364 21140 67172
rect 22876 66386 22932 69200
rect 24892 66500 24948 69200
rect 26908 67228 26964 69200
rect 28924 67228 28980 69200
rect 30940 67228 30996 69200
rect 32956 67228 33012 69200
rect 34972 67228 35028 69200
rect 26908 67172 27412 67228
rect 28924 67172 29204 67228
rect 30940 67172 31220 67228
rect 32956 67172 33236 67228
rect 34972 67172 35140 67228
rect 24892 66434 24948 66444
rect 26124 66500 26180 66510
rect 26124 66406 26180 66444
rect 22876 66334 22878 66386
rect 22930 66334 22932 66386
rect 22876 66322 22932 66334
rect 23548 66274 23604 66286
rect 25116 66276 25172 66286
rect 23548 66222 23550 66274
rect 23602 66222 23604 66274
rect 21868 65490 21924 65502
rect 23548 65492 23604 66222
rect 21868 65438 21870 65490
rect 21922 65438 21924 65490
rect 21420 64484 21476 64494
rect 21420 64390 21476 64428
rect 21868 64484 21924 65438
rect 22988 65436 23604 65492
rect 24668 66274 25172 66276
rect 24668 66222 25118 66274
rect 25170 66222 25172 66274
rect 24668 66220 25172 66222
rect 22540 65378 22596 65390
rect 22540 65326 22542 65378
rect 22594 65326 22596 65378
rect 22540 64932 22596 65326
rect 22540 64866 22596 64876
rect 21868 64418 21924 64428
rect 22988 63810 23044 65436
rect 24668 65378 24724 66220
rect 25116 66210 25172 66220
rect 24668 65326 24670 65378
rect 24722 65326 24724 65378
rect 24668 65314 24724 65326
rect 25452 65378 25508 65390
rect 25452 65326 25454 65378
rect 25506 65326 25508 65378
rect 23548 64932 23604 64942
rect 23548 64838 23604 64876
rect 23996 64706 24052 64718
rect 23996 64654 23998 64706
rect 24050 64654 24052 64706
rect 23660 64594 23716 64606
rect 23660 64542 23662 64594
rect 23714 64542 23716 64594
rect 23212 64484 23268 64494
rect 23212 63924 23268 64428
rect 23436 63924 23492 63934
rect 23212 63922 23604 63924
rect 23212 63870 23438 63922
rect 23490 63870 23604 63922
rect 23212 63868 23604 63870
rect 23436 63858 23492 63868
rect 22988 63758 22990 63810
rect 23042 63758 23044 63810
rect 22988 63746 23044 63758
rect 21084 63298 21140 63308
rect 22316 63364 22372 63374
rect 22316 63270 22372 63308
rect 21308 63140 21364 63150
rect 20972 63138 21364 63140
rect 20972 63086 21310 63138
rect 21362 63086 21364 63138
rect 20972 63084 21364 63086
rect 21308 63074 21364 63084
rect 20860 62636 21140 62692
rect 19964 62580 20020 62590
rect 19628 62578 20020 62580
rect 19628 62526 19966 62578
rect 20018 62526 20020 62578
rect 19628 62524 20020 62526
rect 19964 62514 20020 62524
rect 18956 62468 19012 62478
rect 18732 62412 18956 62468
rect 18732 60004 18788 62412
rect 18956 62374 19012 62412
rect 20412 62468 20468 62478
rect 19180 62354 19236 62366
rect 19180 62302 19182 62354
rect 19234 62302 19236 62354
rect 19180 62132 19236 62302
rect 19516 62356 19572 62366
rect 19852 62356 19908 62366
rect 19572 62354 19908 62356
rect 19572 62302 19854 62354
rect 19906 62302 19908 62354
rect 19572 62300 19908 62302
rect 19516 62262 19572 62300
rect 19852 62290 19908 62300
rect 20076 62354 20132 62366
rect 20076 62302 20078 62354
rect 20130 62302 20132 62354
rect 20076 62132 20132 62302
rect 20412 62354 20468 62412
rect 20860 62468 20916 62478
rect 20860 62374 20916 62412
rect 20412 62302 20414 62354
rect 20466 62302 20468 62354
rect 20412 62290 20468 62302
rect 19180 62076 20132 62132
rect 19180 61572 19236 62076
rect 20300 61796 20356 61806
rect 20300 61794 21028 61796
rect 20300 61742 20302 61794
rect 20354 61742 21028 61794
rect 20300 61740 21028 61742
rect 20300 61730 20356 61740
rect 18844 61516 19236 61572
rect 18844 60674 18900 61516
rect 19964 61460 20020 61470
rect 18844 60622 18846 60674
rect 18898 60622 18900 60674
rect 18844 60340 18900 60622
rect 18844 60274 18900 60284
rect 18956 61458 20020 61460
rect 18956 61406 19966 61458
rect 20018 61406 20020 61458
rect 18956 61404 20020 61406
rect 18956 60226 19012 61404
rect 19964 61394 20020 61404
rect 20412 61458 20468 61470
rect 20412 61406 20414 61458
rect 20466 61406 20468 61458
rect 20188 61348 20244 61358
rect 20412 61348 20468 61406
rect 20188 61346 20468 61348
rect 20188 61294 20190 61346
rect 20242 61294 20468 61346
rect 20188 61292 20468 61294
rect 20636 61458 20692 61470
rect 20636 61406 20638 61458
rect 20690 61406 20692 61458
rect 20636 61348 20692 61406
rect 20748 61348 20804 61358
rect 20636 61346 20804 61348
rect 20636 61294 20750 61346
rect 20802 61294 20804 61346
rect 20636 61292 20804 61294
rect 20188 61282 20244 61292
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 18956 60174 18958 60226
rect 19010 60174 19012 60226
rect 18956 60162 19012 60174
rect 20188 60340 20244 60350
rect 19852 60116 19908 60126
rect 18844 60004 18900 60014
rect 18732 60002 18900 60004
rect 18732 59950 18846 60002
rect 18898 59950 18900 60002
rect 18732 59948 18900 59950
rect 18844 59938 18900 59948
rect 19852 60002 19908 60060
rect 19852 59950 19854 60002
rect 19906 59950 19908 60002
rect 19852 59938 19908 59950
rect 20188 60002 20244 60284
rect 20188 59950 20190 60002
rect 20242 59950 20244 60002
rect 20188 59938 20244 59950
rect 18508 59724 18900 59780
rect 18172 59378 18228 59388
rect 18060 59266 18116 59276
rect 17724 59166 17726 59218
rect 17778 59166 17780 59218
rect 17724 59154 17780 59166
rect 18060 59108 18116 59118
rect 18060 59014 18116 59052
rect 16716 58660 16772 58670
rect 16604 58658 16772 58660
rect 16604 58606 16718 58658
rect 16770 58606 16772 58658
rect 16604 58604 16772 58606
rect 16716 58594 16772 58604
rect 16156 56978 16548 56980
rect 16156 56926 16158 56978
rect 16210 56926 16548 56978
rect 16156 56924 16548 56926
rect 16156 56914 16212 56924
rect 16492 56866 16548 56924
rect 16492 56814 16494 56866
rect 16546 56814 16548 56866
rect 16492 56802 16548 56814
rect 16604 58324 16660 58334
rect 15932 55860 15988 55870
rect 15932 55766 15988 55804
rect 16044 54404 16100 54414
rect 16044 54310 16100 54348
rect 15708 52388 15764 52398
rect 16156 52388 16212 52398
rect 15708 52386 16212 52388
rect 15708 52334 15710 52386
rect 15762 52334 16158 52386
rect 16210 52334 16212 52386
rect 15708 52332 16212 52334
rect 15708 52322 15764 52332
rect 16156 52322 16212 52332
rect 16492 52388 16548 52398
rect 16492 52294 16548 52332
rect 15932 52164 15988 52174
rect 15932 52070 15988 52108
rect 15596 49868 16100 49924
rect 15484 49756 15764 49812
rect 15596 49588 15652 49598
rect 15596 49028 15652 49532
rect 15260 48302 15262 48354
rect 15314 48302 15316 48354
rect 15260 48290 15316 48302
rect 15372 49026 15652 49028
rect 15372 48974 15598 49026
rect 15650 48974 15652 49026
rect 15372 48972 15652 48974
rect 14924 48242 14980 48254
rect 14924 48190 14926 48242
rect 14978 48190 14980 48242
rect 14924 47460 14980 48190
rect 15372 48130 15428 48972
rect 15596 48962 15652 48972
rect 15484 48244 15540 48254
rect 15484 48150 15540 48188
rect 15372 48078 15374 48130
rect 15426 48078 15428 48130
rect 15372 48066 15428 48078
rect 15708 47908 15764 49756
rect 14924 47394 14980 47404
rect 15260 47852 15764 47908
rect 15820 49138 15876 49150
rect 15820 49086 15822 49138
rect 15874 49086 15876 49138
rect 15036 47348 15092 47358
rect 15036 47254 15092 47292
rect 14812 46834 14868 46844
rect 14476 46284 14644 46340
rect 14700 46676 14756 46686
rect 14028 45556 14084 45566
rect 13916 45500 14028 45556
rect 14028 45490 14084 45500
rect 14476 44884 14532 46284
rect 14364 44828 14532 44884
rect 14588 45220 14644 45230
rect 14700 45220 14756 46620
rect 14924 46564 14980 46574
rect 14812 45780 14868 45790
rect 14812 45686 14868 45724
rect 14588 45218 14756 45220
rect 14588 45166 14590 45218
rect 14642 45166 14756 45218
rect 14588 45164 14756 45166
rect 14812 45556 14868 45566
rect 13804 44100 13860 44110
rect 13804 44006 13860 44044
rect 13916 43092 13972 43102
rect 13916 42642 13972 43036
rect 13916 42590 13918 42642
rect 13970 42590 13972 42642
rect 13916 42578 13972 42590
rect 14028 42754 14084 42766
rect 14028 42702 14030 42754
rect 14082 42702 14084 42754
rect 13804 41746 13860 41758
rect 13804 41694 13806 41746
rect 13858 41694 13860 41746
rect 13804 41524 13860 41694
rect 13804 41458 13860 41468
rect 14028 41410 14084 42702
rect 14364 42530 14420 44828
rect 14364 42478 14366 42530
rect 14418 42478 14420 42530
rect 14364 42466 14420 42478
rect 14476 42754 14532 42766
rect 14476 42702 14478 42754
rect 14530 42702 14532 42754
rect 14476 42194 14532 42702
rect 14476 42142 14478 42194
rect 14530 42142 14532 42194
rect 14476 42130 14532 42142
rect 14140 41972 14196 41982
rect 14476 41972 14532 41982
rect 14140 41878 14196 41916
rect 14364 41916 14476 41972
rect 14028 41358 14030 41410
rect 14082 41358 14084 41410
rect 14028 41346 14084 41358
rect 13692 41244 13860 41300
rect 13692 40964 13748 40974
rect 13692 40870 13748 40908
rect 13804 40180 13860 41244
rect 14364 41188 14420 41916
rect 14476 41878 14532 41916
rect 14028 41132 14420 41188
rect 13916 41076 13972 41086
rect 14028 41076 14084 41132
rect 13972 41020 14084 41076
rect 13916 40982 13972 41020
rect 14588 40852 14644 45164
rect 14812 42644 14868 45500
rect 14924 45106 14980 46508
rect 14924 45054 14926 45106
rect 14978 45054 14980 45106
rect 14924 42868 14980 45054
rect 15036 45890 15092 45902
rect 15036 45838 15038 45890
rect 15090 45838 15092 45890
rect 15036 45108 15092 45838
rect 15260 45444 15316 47852
rect 15484 47572 15540 47582
rect 15820 47572 15876 49086
rect 15484 47570 15876 47572
rect 15484 47518 15486 47570
rect 15538 47518 15876 47570
rect 15484 47516 15876 47518
rect 15932 48244 15988 48254
rect 15484 47506 15540 47516
rect 15372 47460 15428 47470
rect 15372 47346 15428 47404
rect 15932 47458 15988 48188
rect 15932 47406 15934 47458
rect 15986 47406 15988 47458
rect 15932 47394 15988 47406
rect 15372 47294 15374 47346
rect 15426 47294 15428 47346
rect 15372 46900 15428 47294
rect 15708 47348 15764 47358
rect 15708 47254 15764 47292
rect 15372 46844 15764 46900
rect 15372 46564 15428 46574
rect 15372 46470 15428 46508
rect 15484 45780 15540 45790
rect 15484 45686 15540 45724
rect 15596 45666 15652 45678
rect 15596 45614 15598 45666
rect 15650 45614 15652 45666
rect 15260 45388 15540 45444
rect 15148 45108 15204 45118
rect 15036 45052 15148 45108
rect 15148 45042 15204 45052
rect 15484 44996 15540 45388
rect 15372 44940 15540 44996
rect 15596 45218 15652 45614
rect 15596 45166 15598 45218
rect 15650 45166 15652 45218
rect 15372 43650 15428 44940
rect 15596 44436 15652 45166
rect 15708 44994 15764 46844
rect 15820 45892 15876 45902
rect 15820 45798 15876 45836
rect 15708 44942 15710 44994
rect 15762 44942 15764 44994
rect 15708 44930 15764 44942
rect 15820 45108 15876 45118
rect 15596 44370 15652 44380
rect 15484 44324 15540 44334
rect 15484 44230 15540 44268
rect 15820 44324 15876 45052
rect 15820 44258 15876 44268
rect 15372 43598 15374 43650
rect 15426 43598 15428 43650
rect 15372 43586 15428 43598
rect 15596 43650 15652 43662
rect 15596 43598 15598 43650
rect 15650 43598 15652 43650
rect 14924 42802 14980 42812
rect 15372 42754 15428 42766
rect 15372 42702 15374 42754
rect 15426 42702 15428 42754
rect 14812 42588 14980 42644
rect 14812 41970 14868 41982
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 41860 14868 41918
rect 14364 40796 14644 40852
rect 14700 41298 14756 41310
rect 14700 41246 14702 41298
rect 14754 41246 14756 41298
rect 14700 41188 14756 41246
rect 14028 40628 14084 40638
rect 14028 40534 14084 40572
rect 13804 40114 13860 40124
rect 14140 39620 14196 39630
rect 14140 39526 14196 39564
rect 13580 38612 13748 38668
rect 13692 38274 13748 38612
rect 13692 38222 13694 38274
rect 13746 38222 13748 38274
rect 13692 38210 13748 38222
rect 14028 38052 14084 38062
rect 14028 37958 14084 37996
rect 14252 35140 14308 35150
rect 14364 35140 14420 40796
rect 13468 35084 13636 35140
rect 13468 34916 13524 34926
rect 13468 34822 13524 34860
rect 12908 34804 12964 34814
rect 12908 34710 12964 34748
rect 12796 33518 12798 33570
rect 12850 33518 12852 33570
rect 12796 33506 12852 33518
rect 13132 33908 13188 33918
rect 12236 33294 12238 33346
rect 12290 33294 12292 33346
rect 12236 32340 12292 33294
rect 12796 33346 12852 33358
rect 12796 33294 12798 33346
rect 12850 33294 12852 33346
rect 12796 33124 12852 33294
rect 12460 32676 12516 32686
rect 12460 32562 12516 32620
rect 12460 32510 12462 32562
rect 12514 32510 12516 32562
rect 12460 32498 12516 32510
rect 12796 32562 12852 33068
rect 13132 32786 13188 33852
rect 13468 33124 13524 33134
rect 13468 33030 13524 33068
rect 13132 32734 13134 32786
rect 13186 32734 13188 32786
rect 13132 32722 13188 32734
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12236 32284 12516 32340
rect 11900 32172 12292 32228
rect 12236 32002 12292 32172
rect 12236 31950 12238 32002
rect 12290 31950 12292 32002
rect 12236 31938 12292 31950
rect 11788 30930 11844 30940
rect 12348 31554 12404 31566
rect 12348 31502 12350 31554
rect 12402 31502 12404 31554
rect 11452 30324 11508 30828
rect 11452 30268 11844 30324
rect 11228 29374 11230 29426
rect 11282 29374 11284 29426
rect 11228 28868 11284 29374
rect 11228 28802 11284 28812
rect 11004 28590 11006 28642
rect 11058 28590 11060 28642
rect 11004 28308 11060 28590
rect 11788 28308 11844 30268
rect 11004 28242 11060 28252
rect 11676 28252 11844 28308
rect 11900 30212 11956 30222
rect 11900 30098 11956 30156
rect 11900 30046 11902 30098
rect 11954 30046 11956 30098
rect 11452 28084 11508 28094
rect 11452 27990 11508 28028
rect 10892 27860 10948 27870
rect 11340 27860 11396 27870
rect 10892 27858 11396 27860
rect 10892 27806 10894 27858
rect 10946 27806 11342 27858
rect 11394 27806 11396 27858
rect 10892 27804 11396 27806
rect 11676 27860 11732 28252
rect 11788 28084 11844 28094
rect 11788 27990 11844 28028
rect 11676 27804 11844 27860
rect 10892 26964 10948 27804
rect 11340 27794 11396 27804
rect 10892 26898 10948 26908
rect 11788 26908 11844 27804
rect 11900 27748 11956 30046
rect 12348 29988 12404 31502
rect 12460 31218 12516 32284
rect 12572 31668 12628 31678
rect 12796 31668 12852 32510
rect 13020 32674 13076 32686
rect 13020 32622 13022 32674
rect 13074 32622 13076 32674
rect 13020 31892 13076 32622
rect 13020 31826 13076 31836
rect 13468 31778 13524 31790
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 12796 31612 13188 31668
rect 12572 31574 12628 31612
rect 12460 31166 12462 31218
rect 12514 31166 12516 31218
rect 12460 31154 12516 31166
rect 12908 30996 12964 31006
rect 12684 30884 12740 30894
rect 12684 30790 12740 30828
rect 12908 30210 12964 30940
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30146 12964 30158
rect 12796 29988 12852 29998
rect 12348 29986 12852 29988
rect 12348 29934 12798 29986
rect 12850 29934 12852 29986
rect 12348 29932 12852 29934
rect 12012 29428 12068 29438
rect 12796 29428 12852 29932
rect 13020 29428 13076 29438
rect 12796 29426 13076 29428
rect 12796 29374 13022 29426
rect 13074 29374 13076 29426
rect 12796 29372 13076 29374
rect 12012 29334 12068 29372
rect 13020 29362 13076 29372
rect 12012 28868 12068 28878
rect 12012 28774 12068 28812
rect 12348 28642 12404 28654
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 12348 28084 12404 28590
rect 12348 28018 12404 28028
rect 12572 28532 12628 28542
rect 12348 27748 12404 27758
rect 11900 27746 12404 27748
rect 11900 27694 12350 27746
rect 12402 27694 12404 27746
rect 11900 27692 12404 27694
rect 12348 27682 12404 27692
rect 12460 27188 12516 27198
rect 12572 27188 12628 28476
rect 12684 28084 12740 28094
rect 12684 27858 12740 28028
rect 12796 28084 12852 28094
rect 13132 28084 13188 31612
rect 13468 31106 13524 31726
rect 13468 31054 13470 31106
rect 13522 31054 13524 31106
rect 13468 30212 13524 31054
rect 13580 30436 13636 35084
rect 14252 35138 14420 35140
rect 14252 35086 14254 35138
rect 14306 35086 14420 35138
rect 14252 35084 14420 35086
rect 14476 40404 14532 40414
rect 14252 35074 14308 35084
rect 13692 34802 13748 34814
rect 13692 34750 13694 34802
rect 13746 34750 13748 34802
rect 13692 33908 13748 34750
rect 13804 34804 13860 34814
rect 13804 34710 13860 34748
rect 13692 33842 13748 33852
rect 13916 34132 13972 34142
rect 13580 30370 13636 30380
rect 13692 33684 13748 33694
rect 13580 30212 13636 30222
rect 13468 30156 13580 30212
rect 13580 30118 13636 30156
rect 13692 29988 13748 33628
rect 13916 33458 13972 34076
rect 14476 34018 14532 40348
rect 14588 39620 14644 39630
rect 14700 39620 14756 41132
rect 14812 40964 14868 41804
rect 14812 40898 14868 40908
rect 14924 39842 14980 42588
rect 15372 42196 15428 42702
rect 15596 42308 15652 43598
rect 15708 43540 15764 43550
rect 15708 43538 15876 43540
rect 15708 43486 15710 43538
rect 15762 43486 15876 43538
rect 15708 43484 15876 43486
rect 15708 43474 15764 43484
rect 15708 42754 15764 42766
rect 15708 42702 15710 42754
rect 15762 42702 15764 42754
rect 15708 42420 15764 42702
rect 15820 42756 15876 43484
rect 15932 42756 15988 42794
rect 15820 42700 15932 42756
rect 15932 42690 15988 42700
rect 15932 42532 15988 42542
rect 15820 42420 15876 42430
rect 15708 42364 15820 42420
rect 15820 42354 15876 42364
rect 15596 42252 15764 42308
rect 15372 42140 15652 42196
rect 15260 41972 15316 41982
rect 15260 41878 15316 41916
rect 15148 40964 15204 40974
rect 15372 40964 15428 42140
rect 15596 42082 15652 42140
rect 15596 42030 15598 42082
rect 15650 42030 15652 42082
rect 15596 42018 15652 42030
rect 15484 41972 15540 41982
rect 15484 41878 15540 41916
rect 15708 41748 15764 42252
rect 15708 41682 15764 41692
rect 15932 41970 15988 42476
rect 15932 41918 15934 41970
rect 15986 41918 15988 41970
rect 15148 40962 15428 40964
rect 15148 40910 15150 40962
rect 15202 40910 15428 40962
rect 15148 40908 15428 40910
rect 15820 41188 15876 41198
rect 15148 40898 15204 40908
rect 14924 39790 14926 39842
rect 14978 39790 14980 39842
rect 14924 39778 14980 39790
rect 15036 40402 15092 40414
rect 15036 40350 15038 40402
rect 15090 40350 15092 40402
rect 14924 39620 14980 39630
rect 14700 39618 14980 39620
rect 14700 39566 14926 39618
rect 14978 39566 14980 39618
rect 14700 39564 14980 39566
rect 14588 38276 14644 39564
rect 14924 39554 14980 39564
rect 14588 38210 14644 38220
rect 14812 38052 14868 38062
rect 14812 37958 14868 37996
rect 14700 37938 14756 37950
rect 14700 37886 14702 37938
rect 14754 37886 14756 37938
rect 14700 37380 14756 37886
rect 15036 37492 15092 40350
rect 15148 40180 15204 40190
rect 15148 40086 15204 40124
rect 15148 38500 15204 38510
rect 15148 37828 15204 38444
rect 15260 38052 15316 40908
rect 15820 40402 15876 41132
rect 15820 40350 15822 40402
rect 15874 40350 15876 40402
rect 15820 40338 15876 40350
rect 15932 40180 15988 41918
rect 15596 40124 15988 40180
rect 15484 39618 15540 39630
rect 15484 39566 15486 39618
rect 15538 39566 15540 39618
rect 15484 39508 15540 39566
rect 15484 39442 15540 39452
rect 15596 39284 15652 40124
rect 16044 39732 16100 49868
rect 16268 49252 16324 49262
rect 16268 49138 16324 49196
rect 16268 49086 16270 49138
rect 16322 49086 16324 49138
rect 16268 49074 16324 49086
rect 16268 45780 16324 45790
rect 16268 44546 16324 45724
rect 16268 44494 16270 44546
rect 16322 44494 16324 44546
rect 16268 44482 16324 44494
rect 16156 44324 16212 44334
rect 16156 44230 16212 44268
rect 16604 43708 16660 58268
rect 17276 56756 17332 56766
rect 17276 56754 17892 56756
rect 17276 56702 17278 56754
rect 17330 56702 17892 56754
rect 17276 56700 17892 56702
rect 17276 56690 17332 56700
rect 17836 55970 17892 56700
rect 17836 55918 17838 55970
rect 17890 55918 17892 55970
rect 17836 55906 17892 55918
rect 17948 56194 18004 56206
rect 17948 56142 17950 56194
rect 18002 56142 18004 56194
rect 17948 55468 18004 56142
rect 18172 55972 18228 55982
rect 18732 55972 18788 55982
rect 18172 55970 18788 55972
rect 18172 55918 18174 55970
rect 18226 55918 18734 55970
rect 18786 55918 18788 55970
rect 18172 55916 18788 55918
rect 18172 55906 18228 55916
rect 18732 55906 18788 55916
rect 18844 55468 18900 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 20300 59220 20356 61292
rect 20748 61282 20804 61292
rect 20972 60898 21028 61740
rect 20972 60846 20974 60898
rect 21026 60846 21028 60898
rect 20972 60834 21028 60846
rect 21084 60676 21140 62636
rect 20300 59154 20356 59164
rect 20524 60620 21140 60676
rect 21756 61570 21812 61582
rect 21756 61518 21758 61570
rect 21810 61518 21812 61570
rect 21756 60786 21812 61518
rect 22428 61460 22484 61470
rect 22428 61458 22596 61460
rect 22428 61406 22430 61458
rect 22482 61406 22596 61458
rect 22428 61404 22596 61406
rect 22428 61394 22484 61404
rect 21756 60734 21758 60786
rect 21810 60734 21812 60786
rect 21756 60676 21812 60734
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19740 57876 19796 57886
rect 19628 57764 19684 57774
rect 19516 57762 19684 57764
rect 19516 57710 19630 57762
rect 19682 57710 19684 57762
rect 19516 57708 19684 57710
rect 19404 57652 19460 57662
rect 19404 57558 19460 57596
rect 19068 57540 19124 57550
rect 19068 56194 19124 57484
rect 19516 57092 19572 57708
rect 19628 57698 19684 57708
rect 19740 57762 19796 57820
rect 20300 57876 20356 57886
rect 20356 57820 20468 57876
rect 20300 57810 20356 57820
rect 19740 57710 19742 57762
rect 19794 57710 19796 57762
rect 19740 57698 19796 57710
rect 20076 57650 20132 57662
rect 20076 57598 20078 57650
rect 20130 57598 20132 57650
rect 19516 57036 20020 57092
rect 19404 56980 19460 56990
rect 19516 56980 19572 57036
rect 19404 56978 19572 56980
rect 19404 56926 19406 56978
rect 19458 56926 19572 56978
rect 19404 56924 19572 56926
rect 19404 56914 19460 56924
rect 19852 56868 19908 56878
rect 19852 56756 19908 56812
rect 19068 56142 19070 56194
rect 19122 56142 19124 56194
rect 19068 56130 19124 56142
rect 19628 56754 19908 56756
rect 19628 56702 19854 56754
rect 19906 56702 19908 56754
rect 19628 56700 19908 56702
rect 17948 55412 18116 55468
rect 18844 55412 19572 55468
rect 18060 55076 18116 55412
rect 18396 55076 18452 55086
rect 18060 55074 18452 55076
rect 18060 55022 18398 55074
rect 18450 55022 18452 55074
rect 18060 55020 18452 55022
rect 17836 53844 17892 53854
rect 17836 53730 17892 53788
rect 17836 53678 17838 53730
rect 17890 53678 17892 53730
rect 17836 53666 17892 53678
rect 17948 53620 18004 53630
rect 17948 53526 18004 53564
rect 18060 53396 18116 55020
rect 18396 55010 18452 55020
rect 18284 54516 18340 54526
rect 18284 54422 18340 54460
rect 19068 54516 19124 54526
rect 18732 53844 18788 53854
rect 18732 53750 18788 53788
rect 18396 53730 18452 53742
rect 18396 53678 18398 53730
rect 18450 53678 18452 53730
rect 17948 53340 18116 53396
rect 18172 53506 18228 53518
rect 18172 53454 18174 53506
rect 18226 53454 18228 53506
rect 17500 52948 17556 52958
rect 17500 52854 17556 52892
rect 17388 49140 17444 49150
rect 17388 49046 17444 49084
rect 16716 49028 16772 49038
rect 16716 48934 16772 48972
rect 17500 47570 17556 47582
rect 17500 47518 17502 47570
rect 17554 47518 17556 47570
rect 17500 46564 17556 47518
rect 17836 47458 17892 47470
rect 17836 47406 17838 47458
rect 17890 47406 17892 47458
rect 17836 47348 17892 47406
rect 17836 46674 17892 47292
rect 17836 46622 17838 46674
rect 17890 46622 17892 46674
rect 17724 46564 17780 46574
rect 17500 46562 17780 46564
rect 17500 46510 17726 46562
rect 17778 46510 17780 46562
rect 17500 46508 17780 46510
rect 17724 46002 17780 46508
rect 17724 45950 17726 46002
rect 17778 45950 17780 46002
rect 17052 45892 17108 45902
rect 17052 45798 17108 45836
rect 17724 45780 17780 45950
rect 17836 45890 17892 46622
rect 17836 45838 17838 45890
rect 17890 45838 17892 45890
rect 17836 45826 17892 45838
rect 17724 45714 17780 45724
rect 16828 45332 16884 45342
rect 16828 44434 16884 45276
rect 16828 44382 16830 44434
rect 16882 44382 16884 44434
rect 16828 44370 16884 44382
rect 17276 44322 17332 44334
rect 17276 44270 17278 44322
rect 17330 44270 17332 44322
rect 16380 43652 16436 43662
rect 16380 43558 16436 43596
rect 16492 43652 16660 43708
rect 16940 44210 16996 44222
rect 16940 44158 16942 44210
rect 16994 44158 16996 44210
rect 16492 43426 16548 43652
rect 16492 43374 16494 43426
rect 16546 43374 16548 43426
rect 16492 43362 16548 43374
rect 16940 43540 16996 44158
rect 16156 43314 16212 43326
rect 16156 43262 16158 43314
rect 16210 43262 16212 43314
rect 16156 41188 16212 43262
rect 16828 42868 16884 42878
rect 16828 42774 16884 42812
rect 16492 42756 16548 42766
rect 16492 42662 16548 42700
rect 16828 42642 16884 42654
rect 16828 42590 16830 42642
rect 16882 42590 16884 42642
rect 16828 42532 16884 42590
rect 16828 42466 16884 42476
rect 16156 41122 16212 41132
rect 16268 42420 16324 42430
rect 16268 40404 16324 42364
rect 16716 41970 16772 41982
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16380 41748 16436 41758
rect 16380 41074 16436 41692
rect 16716 41300 16772 41918
rect 16716 41234 16772 41244
rect 16940 41636 16996 43484
rect 17276 42980 17332 44270
rect 17500 44324 17556 44334
rect 17276 42914 17332 42924
rect 17388 43426 17444 43438
rect 17388 43374 17390 43426
rect 17442 43374 17444 43426
rect 17388 41860 17444 43374
rect 17388 41794 17444 41804
rect 16380 41022 16382 41074
rect 16434 41022 16436 41074
rect 16380 41010 16436 41022
rect 16940 40740 16996 41580
rect 16604 40684 16996 40740
rect 17388 41186 17444 41198
rect 17388 41134 17390 41186
rect 17442 41134 17444 41186
rect 15484 39228 15652 39284
rect 15708 39676 16100 39732
rect 16156 40348 16436 40404
rect 15372 38612 15428 38622
rect 15372 38518 15428 38556
rect 15484 38500 15540 39228
rect 15484 38434 15540 38444
rect 15596 38834 15652 38846
rect 15596 38782 15598 38834
rect 15650 38782 15652 38834
rect 15372 38276 15428 38286
rect 15372 38182 15428 38220
rect 15596 38164 15652 38782
rect 15596 38098 15652 38108
rect 15372 38052 15428 38062
rect 15260 38050 15428 38052
rect 15260 37998 15374 38050
rect 15426 37998 15428 38050
rect 15260 37996 15428 37998
rect 15260 37828 15316 37838
rect 15148 37772 15260 37828
rect 15260 37762 15316 37772
rect 15148 37492 15204 37502
rect 15036 37490 15204 37492
rect 15036 37438 15150 37490
rect 15202 37438 15204 37490
rect 15036 37436 15204 37438
rect 15148 37426 15204 37436
rect 14812 37380 14868 37390
rect 14700 37324 14812 37380
rect 14812 37286 14868 37324
rect 14924 37378 14980 37390
rect 14924 37326 14926 37378
rect 14978 37326 14980 37378
rect 14924 35700 14980 37326
rect 15372 35924 15428 37996
rect 15484 38052 15540 38062
rect 15484 37490 15540 37996
rect 15484 37438 15486 37490
rect 15538 37438 15540 37490
rect 15484 37426 15540 37438
rect 15596 37716 15652 37726
rect 15484 37268 15540 37278
rect 15484 37174 15540 37212
rect 15596 37266 15652 37660
rect 15596 37214 15598 37266
rect 15650 37214 15652 37266
rect 15596 37202 15652 37214
rect 15708 36708 15764 39676
rect 16156 39508 16212 40348
rect 16380 39620 16436 40348
rect 16492 40180 16548 40190
rect 16492 40086 16548 40124
rect 16380 39554 16436 39564
rect 15932 39452 16212 39508
rect 16492 39508 16548 39518
rect 15820 38836 15876 38846
rect 15820 38722 15876 38780
rect 15820 38670 15822 38722
rect 15874 38670 15876 38722
rect 15820 38658 15876 38670
rect 15932 37716 15988 39452
rect 16492 39284 16548 39452
rect 16156 39228 16548 39284
rect 16156 38668 16212 39228
rect 16604 39172 16660 40684
rect 15932 37650 15988 37660
rect 16044 38612 16212 38668
rect 16268 39116 16660 39172
rect 16716 40514 16772 40526
rect 16716 40462 16718 40514
rect 16770 40462 16772 40514
rect 16044 38276 16100 38612
rect 16044 37268 16100 38220
rect 16044 37202 16100 37212
rect 16156 38164 16212 38174
rect 15820 37156 15876 37166
rect 15820 37062 15876 37100
rect 15708 36652 15876 36708
rect 15708 36482 15764 36494
rect 15708 36430 15710 36482
rect 15762 36430 15764 36482
rect 15708 36372 15764 36430
rect 15708 36306 15764 36316
rect 15596 35924 15652 35934
rect 15372 35922 15652 35924
rect 15372 35870 15598 35922
rect 15650 35870 15652 35922
rect 15372 35868 15652 35870
rect 15596 35858 15652 35868
rect 14924 35634 14980 35644
rect 15820 35252 15876 36652
rect 16156 36706 16212 38108
rect 16268 37156 16324 39116
rect 16380 38834 16436 38846
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 16380 37268 16436 38782
rect 16716 38836 16772 40462
rect 17388 40180 17444 41134
rect 17500 41074 17556 44268
rect 17836 44322 17892 44334
rect 17836 44270 17838 44322
rect 17890 44270 17892 44322
rect 17724 43650 17780 43662
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 17612 43540 17668 43550
rect 17612 43446 17668 43484
rect 17724 42532 17780 43598
rect 17500 41022 17502 41074
rect 17554 41022 17556 41074
rect 17500 41010 17556 41022
rect 17612 42476 17780 42532
rect 17500 40404 17556 40414
rect 17612 40404 17668 42476
rect 17836 42196 17892 44270
rect 17948 42420 18004 53340
rect 18172 53058 18228 53454
rect 18396 53508 18452 53678
rect 19068 53618 19124 54460
rect 19068 53566 19070 53618
rect 19122 53566 19124 53618
rect 19068 53554 19124 53566
rect 19404 53620 19460 53630
rect 18620 53508 18676 53518
rect 18396 53506 18676 53508
rect 18396 53454 18622 53506
rect 18674 53454 18676 53506
rect 18396 53452 18676 53454
rect 18172 53006 18174 53058
rect 18226 53006 18228 53058
rect 18172 52994 18228 53006
rect 18508 52274 18564 53452
rect 18620 53442 18676 53452
rect 18844 53508 18900 53518
rect 18844 53414 18900 53452
rect 18508 52222 18510 52274
rect 18562 52222 18564 52274
rect 18508 52210 18564 52222
rect 19180 52276 19236 52286
rect 19180 52162 19236 52220
rect 19404 52274 19460 53564
rect 19404 52222 19406 52274
rect 19458 52222 19460 52274
rect 19404 52210 19460 52222
rect 19180 52110 19182 52162
rect 19234 52110 19236 52162
rect 19180 52098 19236 52110
rect 19516 50036 19572 55412
rect 19628 54516 19684 56700
rect 19852 56690 19908 56700
rect 19964 56644 20020 57036
rect 20076 56980 20132 57598
rect 20300 57652 20356 57662
rect 20300 57558 20356 57596
rect 20188 56980 20244 56990
rect 20076 56978 20244 56980
rect 20076 56926 20190 56978
rect 20242 56926 20244 56978
rect 20076 56924 20244 56926
rect 20188 56914 20244 56924
rect 20300 56868 20356 56878
rect 20412 56868 20468 57820
rect 20524 57874 20580 60620
rect 21756 59668 21812 60620
rect 22540 60228 22596 61404
rect 22652 61348 22708 61358
rect 22652 60786 22708 61292
rect 22652 60734 22654 60786
rect 22706 60734 22708 60786
rect 22652 60722 22708 60734
rect 23212 60676 23268 60686
rect 23212 60582 23268 60620
rect 23548 60676 23604 63868
rect 23660 63812 23716 64542
rect 23996 64484 24052 64654
rect 23996 64418 24052 64428
rect 24780 64594 24836 64606
rect 24780 64542 24782 64594
rect 24834 64542 24836 64594
rect 23660 63746 23716 63756
rect 24780 63252 24836 64542
rect 25452 64484 25508 65326
rect 27356 65378 27412 67172
rect 29148 66162 29204 67172
rect 29148 66110 29150 66162
rect 29202 66110 29204 66162
rect 29148 66098 29204 66110
rect 31164 66162 31220 67172
rect 31164 66110 31166 66162
rect 31218 66110 31220 66162
rect 31164 66098 31220 66110
rect 33180 66162 33236 67172
rect 33180 66110 33182 66162
rect 33234 66110 33236 66162
rect 33180 66098 33236 66110
rect 35084 66164 35140 67172
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 36988 66386 37044 69200
rect 39004 66500 39060 69200
rect 39004 66434 39060 66444
rect 40796 66500 40852 66510
rect 40796 66406 40852 66444
rect 36988 66334 36990 66386
rect 37042 66334 37044 66386
rect 36988 66322 37044 66334
rect 39228 66276 39284 66286
rect 39788 66276 39844 66286
rect 39228 66274 39396 66276
rect 39228 66222 39230 66274
rect 39282 66222 39396 66274
rect 39228 66220 39396 66222
rect 39228 66210 39284 66220
rect 35196 66164 35252 66174
rect 35084 66162 35252 66164
rect 35084 66110 35198 66162
rect 35250 66110 35252 66162
rect 35084 66108 35252 66110
rect 35196 66098 35252 66108
rect 34860 65602 34916 65614
rect 34860 65550 34862 65602
rect 34914 65550 34916 65602
rect 27356 65326 27358 65378
rect 27410 65326 27412 65378
rect 27356 65314 27412 65326
rect 29708 65490 29764 65502
rect 29708 65438 29710 65490
rect 29762 65438 29764 65490
rect 29708 65380 29764 65438
rect 33740 65492 33796 65502
rect 30268 65380 30324 65390
rect 29708 65378 30324 65380
rect 29708 65326 30270 65378
rect 30322 65326 30324 65378
rect 29708 65324 30324 65326
rect 30268 64932 30324 65324
rect 30268 64866 30324 64876
rect 25452 64418 25508 64428
rect 26908 64818 26964 64830
rect 33516 64820 33572 64830
rect 26908 64766 26910 64818
rect 26962 64766 26964 64818
rect 26684 64260 26740 64270
rect 26908 64260 26964 64766
rect 32508 64818 33572 64820
rect 32508 64766 33518 64818
rect 33570 64766 33572 64818
rect 32508 64764 33572 64766
rect 27804 64708 27860 64718
rect 26740 64204 26964 64260
rect 27244 64482 27300 64494
rect 27244 64430 27246 64482
rect 27298 64430 27300 64482
rect 26684 63922 26740 64204
rect 26684 63870 26686 63922
rect 26738 63870 26740 63922
rect 26684 63858 26740 63870
rect 26348 63810 26404 63822
rect 27132 63812 27188 63822
rect 26348 63758 26350 63810
rect 26402 63758 26404 63810
rect 26348 63700 26404 63758
rect 24780 63186 24836 63196
rect 26236 63252 26292 63262
rect 26236 63158 26292 63196
rect 26124 63026 26180 63038
rect 26124 62974 26126 63026
rect 26178 62974 26180 63026
rect 26124 62916 26180 62974
rect 26124 62850 26180 62860
rect 25900 62132 25956 62142
rect 24556 61682 24612 61694
rect 24556 61630 24558 61682
rect 24610 61630 24612 61682
rect 24556 61460 24612 61630
rect 24892 61460 24948 61470
rect 24556 61458 24948 61460
rect 24556 61406 24894 61458
rect 24946 61406 24948 61458
rect 24556 61404 24948 61406
rect 23548 60610 23604 60620
rect 22652 60228 22708 60238
rect 22540 60226 22708 60228
rect 22540 60174 22654 60226
rect 22706 60174 22708 60226
rect 22540 60172 22708 60174
rect 22652 60162 22708 60172
rect 23996 60002 24052 60014
rect 23996 59950 23998 60002
rect 24050 59950 24052 60002
rect 22988 59892 23044 59902
rect 23324 59892 23380 59902
rect 22988 59890 23380 59892
rect 22988 59838 22990 59890
rect 23042 59838 23326 59890
rect 23378 59838 23380 59890
rect 22988 59836 23380 59838
rect 22988 59826 23044 59836
rect 23324 59826 23380 59836
rect 23996 59892 24052 59950
rect 21980 59778 22036 59790
rect 21980 59726 21982 59778
rect 22034 59726 22036 59778
rect 21980 59668 22036 59726
rect 22764 59780 22820 59790
rect 22764 59778 22932 59780
rect 22764 59726 22766 59778
rect 22818 59726 22932 59778
rect 22764 59724 22932 59726
rect 22764 59714 22820 59724
rect 21756 59612 22036 59668
rect 20524 57822 20526 57874
rect 20578 57822 20580 57874
rect 20524 57810 20580 57822
rect 21084 59220 21140 59230
rect 20748 57764 20804 57774
rect 20748 57650 20804 57708
rect 20748 57598 20750 57650
rect 20802 57598 20804 57650
rect 20748 57586 20804 57598
rect 20748 56868 20804 56878
rect 20300 56866 20692 56868
rect 20300 56814 20302 56866
rect 20354 56814 20692 56866
rect 20300 56812 20692 56814
rect 20300 56802 20356 56812
rect 20076 56644 20132 56682
rect 19964 56642 20244 56644
rect 19964 56590 20078 56642
rect 20130 56590 20244 56642
rect 19964 56588 20244 56590
rect 20076 56578 20132 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 56196 20244 56588
rect 20300 56196 20356 56206
rect 20188 56194 20356 56196
rect 20188 56142 20302 56194
rect 20354 56142 20356 56194
rect 20188 56140 20356 56142
rect 20300 56130 20356 56140
rect 20636 55972 20692 56812
rect 20748 56774 20804 56812
rect 20748 55972 20804 55982
rect 20636 55970 20804 55972
rect 20636 55918 20750 55970
rect 20802 55918 20804 55970
rect 20636 55916 20804 55918
rect 20748 55906 20804 55916
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19628 54450 19684 54460
rect 20524 53844 20580 53854
rect 19852 53732 19908 53742
rect 19852 53638 19908 53676
rect 19964 53732 20020 53742
rect 19964 53730 20468 53732
rect 19964 53678 19966 53730
rect 20018 53678 20468 53730
rect 19964 53676 20468 53678
rect 19964 53666 20020 53676
rect 19628 53508 19684 53518
rect 19628 53172 19684 53452
rect 20076 53508 20132 53546
rect 20300 53508 20356 53518
rect 20076 53442 20132 53452
rect 20188 53506 20356 53508
rect 20188 53454 20302 53506
rect 20354 53454 20356 53506
rect 20188 53452 20356 53454
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19628 53116 20132 53172
rect 20076 52052 20132 53116
rect 20188 52274 20244 53452
rect 20300 53442 20356 53452
rect 20188 52222 20190 52274
rect 20242 52222 20244 52274
rect 20188 52210 20244 52222
rect 20300 52836 20356 52846
rect 20300 52276 20356 52780
rect 20412 52386 20468 53676
rect 20524 53506 20580 53788
rect 20636 53620 20692 53630
rect 20636 53526 20692 53564
rect 20524 53454 20526 53506
rect 20578 53454 20580 53506
rect 20524 52836 20580 53454
rect 20636 53284 20692 53294
rect 20636 52948 20692 53228
rect 20636 52854 20692 52892
rect 20524 52770 20580 52780
rect 20412 52334 20414 52386
rect 20466 52334 20468 52386
rect 20412 52322 20468 52334
rect 20300 52210 20356 52220
rect 20748 52276 20804 52286
rect 20748 52182 20804 52220
rect 20076 51996 20356 52052
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19516 49970 19572 49980
rect 19628 50482 19684 50494
rect 19628 50430 19630 50482
rect 19682 50430 19684 50482
rect 19292 49924 19348 49934
rect 19292 49830 19348 49868
rect 19180 49810 19236 49822
rect 19180 49758 19182 49810
rect 19234 49758 19236 49810
rect 19180 49700 19236 49758
rect 19516 49812 19572 49822
rect 19516 49718 19572 49756
rect 19180 49364 19236 49644
rect 19180 49308 19348 49364
rect 19068 49028 19124 49038
rect 19068 48466 19124 48972
rect 19068 48414 19070 48466
rect 19122 48414 19124 48466
rect 18284 47348 18340 47358
rect 18284 47254 18340 47292
rect 18508 46900 18564 46910
rect 18396 45780 18452 45790
rect 18396 45686 18452 45724
rect 18508 44324 18564 46844
rect 18508 44230 18564 44268
rect 19068 46004 19124 48414
rect 19292 48244 19348 49308
rect 19516 49140 19572 49150
rect 19628 49140 19684 50430
rect 19740 50372 19796 50382
rect 19740 50370 20244 50372
rect 19740 50318 19742 50370
rect 19794 50318 20244 50370
rect 19740 50316 20244 50318
rect 19740 50306 19796 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20188 49924 20244 50316
rect 20188 49810 20244 49868
rect 20300 49922 20356 51996
rect 20300 49870 20302 49922
rect 20354 49870 20356 49922
rect 20300 49858 20356 49870
rect 20188 49758 20190 49810
rect 20242 49758 20244 49810
rect 19516 49138 19684 49140
rect 19516 49086 19518 49138
rect 19570 49086 19684 49138
rect 19516 49084 19684 49086
rect 20076 49140 20132 49150
rect 19516 49074 19572 49084
rect 20076 49046 20132 49084
rect 19964 48916 20020 48926
rect 19964 48822 20020 48860
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48468 20244 49758
rect 20524 49700 20580 49710
rect 20524 49606 20580 49644
rect 20300 48914 20356 48926
rect 20300 48862 20302 48914
rect 20354 48862 20356 48914
rect 20300 48692 20356 48862
rect 20524 48916 20580 48926
rect 20524 48822 20580 48860
rect 20300 48626 20356 48636
rect 20412 48804 20468 48814
rect 19964 48412 20244 48468
rect 19516 48244 19572 48254
rect 19292 48242 19572 48244
rect 19292 48190 19518 48242
rect 19570 48190 19572 48242
rect 19292 48188 19572 48190
rect 19516 48178 19572 48188
rect 19964 48242 20020 48412
rect 20412 48354 20468 48748
rect 20972 48468 21028 48478
rect 20972 48374 21028 48412
rect 20412 48302 20414 48354
rect 20466 48302 20468 48354
rect 20412 48290 20468 48302
rect 19964 48190 19966 48242
rect 20018 48190 20020 48242
rect 19964 48178 20020 48190
rect 21084 47236 21140 59164
rect 21308 56868 21364 56878
rect 21756 56868 21812 59612
rect 22876 57762 22932 59724
rect 22876 57710 22878 57762
rect 22930 57710 22932 57762
rect 22764 57652 22820 57662
rect 22092 57650 22820 57652
rect 22092 57598 22766 57650
rect 22818 57598 22820 57650
rect 22092 57596 22820 57598
rect 22092 56978 22148 57596
rect 22764 57586 22820 57596
rect 22092 56926 22094 56978
rect 22146 56926 22148 56978
rect 22092 56914 22148 56926
rect 22652 57426 22708 57438
rect 22652 57374 22654 57426
rect 22706 57374 22708 57426
rect 21308 56866 21812 56868
rect 21308 56814 21310 56866
rect 21362 56814 21812 56866
rect 21308 56812 21812 56814
rect 21308 55636 21364 56812
rect 22652 56306 22708 57374
rect 22652 56254 22654 56306
rect 22706 56254 22708 56306
rect 22652 56242 22708 56254
rect 21196 53844 21252 53854
rect 21196 53060 21252 53788
rect 21308 53284 21364 55580
rect 22876 55468 22932 57710
rect 23996 57762 24052 59836
rect 24892 59890 24948 61404
rect 25004 61348 25060 61358
rect 25564 61348 25620 61358
rect 25900 61348 25956 62076
rect 26348 61348 26404 63644
rect 27020 63810 27188 63812
rect 27020 63758 27134 63810
rect 27186 63758 27188 63810
rect 27020 63756 27188 63758
rect 26684 63140 26740 63150
rect 26684 63046 26740 63084
rect 26460 63028 26516 63038
rect 26460 62934 26516 62972
rect 27020 62916 27076 63756
rect 27132 63746 27188 63756
rect 27244 63700 27300 64430
rect 27356 64482 27412 64494
rect 27356 64430 27358 64482
rect 27410 64430 27412 64482
rect 27356 64036 27412 64430
rect 27468 64482 27524 64494
rect 27468 64430 27470 64482
rect 27522 64430 27524 64482
rect 27468 64260 27524 64430
rect 27468 64194 27524 64204
rect 27804 64146 27860 64652
rect 27916 64706 27972 64718
rect 27916 64654 27918 64706
rect 27970 64654 27972 64706
rect 27916 64484 27972 64654
rect 29036 64706 29092 64718
rect 29036 64654 29038 64706
rect 29090 64654 29092 64706
rect 28700 64484 28756 64494
rect 29036 64484 29092 64654
rect 27916 64428 28420 64484
rect 27804 64094 27806 64146
rect 27858 64094 27860 64146
rect 27804 64082 27860 64094
rect 28140 64260 28196 64270
rect 27468 64036 27524 64046
rect 27356 64034 27524 64036
rect 27356 63982 27470 64034
rect 27522 63982 27524 64034
rect 27356 63980 27524 63982
rect 27468 63970 27524 63980
rect 27580 64034 27636 64046
rect 27580 63982 27582 64034
rect 27634 63982 27636 64034
rect 27580 63812 27636 63982
rect 28028 63924 28084 63934
rect 27916 63922 28084 63924
rect 27916 63870 28030 63922
rect 28082 63870 28084 63922
rect 27916 63868 28084 63870
rect 27580 63756 27860 63812
rect 27244 63634 27300 63644
rect 27132 63140 27188 63150
rect 27132 63046 27188 63084
rect 27580 63138 27636 63150
rect 27580 63086 27582 63138
rect 27634 63086 27636 63138
rect 27020 62822 27076 62860
rect 27244 63028 27300 63038
rect 27244 62914 27300 62972
rect 27244 62862 27246 62914
rect 27298 62862 27300 62914
rect 27244 62244 27300 62862
rect 27580 62916 27636 63086
rect 27804 63138 27860 63756
rect 27804 63086 27806 63138
rect 27858 63086 27860 63138
rect 27804 63074 27860 63086
rect 27580 62850 27636 62860
rect 27244 62178 27300 62188
rect 27692 62244 27748 62254
rect 27916 62244 27972 63868
rect 28028 63858 28084 63868
rect 28140 63700 28196 64204
rect 28028 63644 28196 63700
rect 28252 63700 28308 63710
rect 28028 63026 28084 63644
rect 28140 63140 28196 63150
rect 28252 63140 28308 63644
rect 28140 63138 28308 63140
rect 28140 63086 28142 63138
rect 28194 63086 28308 63138
rect 28140 63084 28308 63086
rect 28140 63074 28196 63084
rect 28028 62974 28030 63026
rect 28082 62974 28084 63026
rect 28028 62962 28084 62974
rect 27692 62242 27972 62244
rect 27692 62190 27694 62242
rect 27746 62190 27972 62242
rect 27692 62188 27972 62190
rect 28364 62244 28420 64428
rect 28588 64482 29092 64484
rect 28588 64430 28702 64482
rect 28754 64430 29092 64482
rect 28588 64428 29092 64430
rect 29148 64708 29204 64718
rect 27692 62132 27748 62188
rect 28364 62178 28420 62188
rect 28476 62916 28532 62926
rect 28588 62916 28644 64428
rect 28700 64418 28756 64428
rect 28812 63812 28868 63822
rect 28812 63810 29092 63812
rect 28812 63758 28814 63810
rect 28866 63758 29092 63810
rect 28812 63756 29092 63758
rect 28812 63746 28868 63756
rect 28532 62914 28644 62916
rect 28532 62862 28590 62914
rect 28642 62862 28644 62914
rect 28532 62860 28644 62862
rect 27692 62066 27748 62076
rect 25004 61346 25508 61348
rect 25004 61294 25006 61346
rect 25058 61294 25508 61346
rect 25004 61292 25508 61294
rect 25004 61282 25060 61292
rect 25452 61012 25508 61292
rect 25564 61254 25620 61292
rect 25788 61346 25956 61348
rect 25788 61294 25902 61346
rect 25954 61294 25956 61346
rect 25788 61292 25956 61294
rect 25452 60918 25508 60956
rect 25676 60676 25732 60686
rect 25788 60676 25844 61292
rect 25900 61282 25956 61292
rect 26124 61292 26404 61348
rect 26012 61012 26068 61022
rect 26012 60918 26068 60956
rect 25732 60620 25844 60676
rect 25900 60786 25956 60798
rect 25900 60734 25902 60786
rect 25954 60734 25956 60786
rect 25900 60676 25956 60734
rect 25676 60610 25732 60620
rect 25900 60610 25956 60620
rect 25228 60564 25284 60574
rect 25452 60564 25508 60574
rect 25228 60562 25452 60564
rect 25228 60510 25230 60562
rect 25282 60510 25452 60562
rect 25228 60508 25452 60510
rect 25228 60498 25284 60508
rect 25452 60114 25508 60508
rect 25564 60562 25620 60574
rect 25564 60510 25566 60562
rect 25618 60510 25620 60562
rect 25564 60228 25620 60510
rect 25564 60172 25956 60228
rect 25452 60062 25454 60114
rect 25506 60062 25508 60114
rect 25452 60050 25508 60062
rect 25900 60002 25956 60172
rect 25900 59950 25902 60002
rect 25954 59950 25956 60002
rect 25900 59938 25956 59950
rect 24892 59838 24894 59890
rect 24946 59838 24948 59890
rect 24892 59826 24948 59838
rect 26012 59778 26068 59790
rect 26012 59726 26014 59778
rect 26066 59726 26068 59778
rect 25228 58436 25284 58446
rect 25228 57874 25284 58380
rect 25228 57822 25230 57874
rect 25282 57822 25284 57874
rect 25228 57810 25284 57822
rect 25452 57764 25508 57774
rect 23996 57710 23998 57762
rect 24050 57710 24052 57762
rect 23996 57698 24052 57710
rect 25340 57762 25508 57764
rect 25340 57710 25454 57762
rect 25506 57710 25508 57762
rect 25340 57708 25508 57710
rect 23660 57650 23716 57662
rect 23660 57598 23662 57650
rect 23714 57598 23716 57650
rect 22988 56196 23044 56206
rect 22988 56082 23044 56140
rect 23660 56196 23716 57598
rect 24668 57650 24724 57662
rect 24668 57598 24670 57650
rect 24722 57598 24724 57650
rect 23660 56130 23716 56140
rect 23772 57538 23828 57550
rect 23772 57486 23774 57538
rect 23826 57486 23828 57538
rect 22988 56030 22990 56082
rect 23042 56030 23044 56082
rect 22988 56018 23044 56030
rect 22428 55412 22932 55468
rect 23548 55524 23604 55534
rect 23660 55524 23716 55534
rect 23548 55522 23660 55524
rect 23548 55470 23550 55522
rect 23602 55470 23660 55522
rect 23548 55468 23660 55470
rect 23548 55458 23604 55468
rect 23660 55458 23716 55468
rect 22316 53844 22372 53854
rect 22316 53750 22372 53788
rect 22428 53506 22484 55412
rect 23772 55410 23828 57486
rect 24668 57090 24724 57598
rect 25340 57204 25396 57708
rect 25452 57698 25508 57708
rect 25564 57764 25620 57774
rect 25900 57764 25956 57774
rect 25564 57762 25956 57764
rect 25564 57710 25566 57762
rect 25618 57710 25902 57762
rect 25954 57710 25956 57762
rect 25564 57708 25956 57710
rect 25564 57698 25620 57708
rect 25900 57540 25956 57708
rect 26012 57764 26068 59726
rect 26012 57698 26068 57708
rect 26124 57540 26180 61292
rect 28140 61236 28196 61246
rect 27244 60898 27300 60910
rect 27244 60846 27246 60898
rect 27298 60846 27300 60898
rect 26236 60786 26292 60798
rect 26236 60734 26238 60786
rect 26290 60734 26292 60786
rect 26236 60004 26292 60734
rect 27132 60786 27188 60798
rect 27132 60734 27134 60786
rect 27186 60734 27188 60786
rect 27132 60676 27188 60734
rect 26460 60004 26516 60014
rect 26236 60002 26516 60004
rect 26236 59950 26462 60002
rect 26514 59950 26516 60002
rect 26236 59948 26516 59950
rect 26460 59938 26516 59948
rect 26572 59892 26628 59902
rect 26572 59798 26628 59836
rect 27020 59444 27076 59454
rect 27132 59444 27188 60620
rect 27244 60564 27300 60846
rect 27804 60900 27860 60910
rect 27804 60806 27860 60844
rect 27244 60498 27300 60508
rect 27468 60786 27524 60798
rect 27468 60734 27470 60786
rect 27522 60734 27524 60786
rect 27468 60004 27524 60734
rect 27692 60786 27748 60798
rect 27692 60734 27694 60786
rect 27746 60734 27748 60786
rect 27692 60676 27748 60734
rect 27916 60788 27972 60798
rect 27916 60694 27972 60732
rect 27692 60610 27748 60620
rect 28028 60564 28084 60574
rect 27916 60508 28028 60564
rect 27804 60116 27860 60126
rect 27916 60116 27972 60508
rect 28028 60498 28084 60508
rect 27804 60114 27972 60116
rect 27804 60062 27806 60114
rect 27858 60062 27972 60114
rect 27804 60060 27972 60062
rect 27804 60050 27860 60060
rect 27468 59938 27524 59948
rect 28028 60002 28084 60014
rect 28028 59950 28030 60002
rect 28082 59950 28084 60002
rect 27020 59442 27188 59444
rect 27020 59390 27022 59442
rect 27074 59390 27188 59442
rect 27020 59388 27188 59390
rect 27468 59778 27524 59790
rect 27468 59726 27470 59778
rect 27522 59726 27524 59778
rect 27020 59378 27076 59388
rect 27244 59218 27300 59230
rect 27244 59166 27246 59218
rect 27298 59166 27300 59218
rect 27244 59108 27300 59166
rect 27468 59108 27524 59726
rect 27804 59108 27860 59118
rect 28028 59108 28084 59950
rect 27244 59106 28084 59108
rect 27244 59054 27806 59106
rect 27858 59054 28084 59106
rect 27244 59052 28084 59054
rect 26684 58436 26740 58446
rect 26684 58342 26740 58380
rect 26572 58210 26628 58222
rect 26572 58158 26574 58210
rect 26626 58158 26628 58210
rect 25900 57484 26180 57540
rect 26236 57650 26292 57662
rect 26236 57598 26238 57650
rect 26290 57598 26292 57650
rect 24668 57038 24670 57090
rect 24722 57038 24724 57090
rect 24668 57026 24724 57038
rect 25116 57148 25396 57204
rect 24220 56978 24276 56990
rect 24220 56926 24222 56978
rect 24274 56926 24276 56978
rect 24220 56644 24276 56926
rect 24780 56756 24836 56766
rect 25116 56756 25172 57148
rect 25452 56868 25508 56878
rect 26124 56868 26180 56878
rect 25452 56866 26180 56868
rect 25452 56814 25454 56866
rect 25506 56814 26126 56866
rect 26178 56814 26180 56866
rect 25452 56812 26180 56814
rect 26236 56868 26292 57598
rect 26572 56868 26628 58158
rect 27244 57876 27300 59052
rect 27804 59042 27860 59052
rect 27580 58546 27636 58558
rect 27580 58494 27582 58546
rect 27634 58494 27636 58546
rect 26908 57820 27300 57876
rect 27468 58434 27524 58446
rect 27468 58382 27470 58434
rect 27522 58382 27524 58434
rect 26684 56868 26740 56878
rect 26236 56812 26684 56868
rect 25452 56802 25508 56812
rect 24780 56754 25172 56756
rect 24780 56702 24782 56754
rect 24834 56702 25118 56754
rect 25170 56702 25172 56754
rect 24780 56700 25172 56702
rect 24668 56644 24724 56654
rect 24220 56642 24724 56644
rect 24220 56590 24670 56642
rect 24722 56590 24724 56642
rect 24220 56588 24724 56590
rect 23772 55358 23774 55410
rect 23826 55358 23828 55410
rect 23772 55346 23828 55358
rect 23884 56196 23940 56206
rect 24220 56196 24276 56588
rect 24668 56578 24724 56588
rect 24780 56420 24836 56700
rect 25116 56690 25172 56700
rect 23884 56194 24276 56196
rect 23884 56142 23886 56194
rect 23938 56142 24276 56194
rect 23884 56140 24276 56142
rect 24444 56364 24836 56420
rect 23884 55298 23940 56140
rect 23884 55246 23886 55298
rect 23938 55246 23940 55298
rect 23884 55234 23940 55246
rect 24108 55972 24164 55982
rect 23324 53956 23380 53966
rect 23324 53862 23380 53900
rect 24108 53842 24164 55916
rect 24444 55970 24500 56364
rect 24444 55918 24446 55970
rect 24498 55918 24500 55970
rect 24444 55524 24500 55918
rect 24444 55458 24500 55468
rect 25340 55970 25396 55982
rect 25340 55918 25342 55970
rect 25394 55918 25396 55970
rect 25340 55636 25396 55918
rect 24108 53790 24110 53842
rect 24162 53790 24164 53842
rect 24108 53778 24164 53790
rect 24780 53956 24836 53966
rect 23884 53732 23940 53742
rect 24780 53732 24836 53900
rect 23884 53730 24052 53732
rect 23884 53678 23886 53730
rect 23938 53678 24052 53730
rect 23884 53676 24052 53678
rect 23884 53666 23940 53676
rect 22652 53620 22708 53630
rect 22428 53454 22430 53506
rect 22482 53454 22484 53506
rect 21364 53228 21588 53284
rect 21308 53218 21364 53228
rect 21420 53060 21476 53070
rect 21196 53058 21476 53060
rect 21196 53006 21422 53058
rect 21474 53006 21476 53058
rect 21196 53004 21476 53006
rect 21420 52994 21476 53004
rect 21532 52274 21588 53228
rect 21532 52222 21534 52274
rect 21586 52222 21588 52274
rect 21532 52210 21588 52222
rect 22428 51492 22484 53454
rect 22540 53618 22708 53620
rect 22540 53566 22654 53618
rect 22706 53566 22708 53618
rect 22540 53564 22708 53566
rect 22540 51938 22596 53564
rect 22652 53554 22708 53564
rect 23100 53620 23156 53630
rect 23100 53526 23156 53564
rect 23548 53620 23604 53630
rect 23212 53508 23268 53518
rect 23212 53414 23268 53452
rect 23100 52948 23156 52958
rect 23100 52276 23156 52892
rect 23548 52834 23604 53564
rect 23884 53508 23940 53518
rect 23884 53058 23940 53452
rect 23996 53170 24052 53676
rect 24556 53730 24836 53732
rect 24556 53678 24782 53730
rect 24834 53678 24836 53730
rect 24556 53676 24836 53678
rect 23996 53118 23998 53170
rect 24050 53118 24052 53170
rect 23996 53106 24052 53118
rect 24332 53620 24388 53630
rect 23884 53006 23886 53058
rect 23938 53006 23940 53058
rect 23884 52994 23940 53006
rect 24220 52948 24276 52958
rect 24220 52854 24276 52892
rect 23548 52782 23550 52834
rect 23602 52782 23604 52834
rect 23548 52770 23604 52782
rect 23100 52162 23156 52220
rect 23100 52110 23102 52162
rect 23154 52110 23156 52162
rect 23100 52098 23156 52110
rect 24332 52050 24388 53564
rect 24556 52274 24612 53676
rect 24780 53666 24836 53676
rect 25340 53730 25396 55580
rect 25340 53678 25342 53730
rect 25394 53678 25396 53730
rect 24668 53172 24724 53182
rect 24668 53078 24724 53116
rect 25340 53172 25396 53678
rect 25340 53078 25396 53116
rect 24556 52222 24558 52274
rect 24610 52222 24612 52274
rect 24556 52210 24612 52222
rect 24332 51998 24334 52050
rect 24386 51998 24388 52050
rect 24332 51986 24388 51998
rect 22540 51886 22542 51938
rect 22594 51886 22596 51938
rect 22540 51874 22596 51886
rect 22428 51426 22484 51436
rect 23772 51492 23828 51502
rect 21532 49924 21588 49934
rect 21532 49922 21700 49924
rect 21532 49870 21534 49922
rect 21586 49870 21700 49922
rect 21532 49868 21700 49870
rect 21532 49858 21588 49868
rect 21196 49810 21252 49822
rect 21196 49758 21198 49810
rect 21250 49758 21252 49810
rect 21196 49588 21252 49758
rect 21420 49812 21476 49822
rect 21420 49718 21476 49756
rect 21532 49588 21588 49598
rect 21196 49586 21588 49588
rect 21196 49534 21534 49586
rect 21586 49534 21588 49586
rect 21196 49532 21588 49534
rect 21532 49522 21588 49532
rect 21420 48916 21476 48926
rect 21420 48822 21476 48860
rect 21308 48804 21364 48814
rect 21308 48710 21364 48748
rect 21532 48804 21588 48814
rect 21644 48804 21700 49868
rect 23772 49812 23828 51436
rect 25452 50594 25508 50606
rect 25452 50542 25454 50594
rect 25506 50542 25508 50594
rect 25116 50484 25172 50494
rect 25452 50484 25508 50542
rect 25116 50482 25508 50484
rect 25116 50430 25118 50482
rect 25170 50430 25508 50482
rect 25116 50428 25508 50430
rect 23772 49810 24052 49812
rect 23772 49758 23774 49810
rect 23826 49758 24052 49810
rect 23772 49756 24052 49758
rect 23772 49746 23828 49756
rect 23660 49698 23716 49710
rect 23660 49646 23662 49698
rect 23714 49646 23716 49698
rect 23436 49588 23492 49598
rect 22092 49586 23492 49588
rect 22092 49534 23438 49586
rect 23490 49534 23492 49586
rect 22092 49532 23492 49534
rect 21532 48802 21700 48804
rect 21532 48750 21534 48802
rect 21586 48750 21700 48802
rect 21532 48748 21700 48750
rect 21980 49026 22036 49038
rect 21980 48974 21982 49026
rect 22034 48974 22036 49026
rect 21532 48692 21588 48748
rect 21532 47684 21588 48636
rect 21980 48468 22036 48974
rect 21980 48402 22036 48412
rect 22092 48466 22148 49532
rect 23436 49522 23492 49532
rect 23548 49140 23604 49150
rect 22540 49028 22596 49038
rect 22540 48934 22596 48972
rect 22988 49028 23044 49038
rect 22988 48934 23044 48972
rect 22092 48414 22094 48466
rect 22146 48414 22148 48466
rect 22092 48402 22148 48414
rect 23324 48468 23380 48478
rect 23380 48412 23492 48468
rect 23324 48402 23380 48412
rect 21532 47618 21588 47628
rect 22428 48242 22484 48254
rect 22428 48190 22430 48242
rect 22482 48190 22484 48242
rect 22428 47460 22484 48190
rect 22652 47684 22708 47694
rect 22652 47590 22708 47628
rect 23100 47572 23156 47582
rect 23100 47478 23156 47516
rect 22876 47460 22932 47470
rect 22428 47458 22932 47460
rect 22428 47406 22878 47458
rect 22930 47406 22932 47458
rect 22428 47404 22932 47406
rect 21084 47170 21140 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46900 20244 46910
rect 19404 46676 19460 46686
rect 19404 46582 19460 46620
rect 19740 46452 19796 46462
rect 19740 46358 19796 46396
rect 19068 43708 19124 45948
rect 20188 46002 20244 46844
rect 22876 46116 22932 47404
rect 22988 46116 23044 46126
rect 22876 46060 22988 46116
rect 22988 46050 23044 46060
rect 20188 45950 20190 46002
rect 20242 45950 20244 46002
rect 20188 45938 20244 45950
rect 20748 45668 20804 45678
rect 20748 45574 20804 45612
rect 21420 45668 21476 45678
rect 21420 45574 21476 45612
rect 23100 45666 23156 45678
rect 23100 45614 23102 45666
rect 23154 45614 23156 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 22316 45332 22372 45342
rect 22316 45238 22372 45276
rect 21644 45220 21700 45230
rect 21644 45106 21700 45164
rect 21644 45054 21646 45106
rect 21698 45054 21700 45106
rect 20972 44994 21028 45006
rect 20972 44942 20974 44994
rect 21026 44942 21028 44994
rect 19628 44434 19684 44446
rect 19628 44382 19630 44434
rect 19682 44382 19684 44434
rect 19628 43708 19684 44382
rect 20972 44324 21028 44942
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 18284 43650 18340 43662
rect 18284 43598 18286 43650
rect 18338 43598 18340 43650
rect 18284 42980 18340 43598
rect 19068 43652 19684 43708
rect 19068 43538 19124 43652
rect 19068 43486 19070 43538
rect 19122 43486 19124 43538
rect 19068 43474 19124 43486
rect 19628 43204 19684 43652
rect 20524 43652 20580 43662
rect 20580 43596 20692 43652
rect 20524 43586 20580 43596
rect 19740 43428 19796 43438
rect 19740 43334 19796 43372
rect 19628 43138 19684 43148
rect 18060 42924 18340 42980
rect 20188 42980 20244 42990
rect 18060 42644 18116 42924
rect 20188 42886 20244 42924
rect 18172 42756 18228 42766
rect 18172 42754 18564 42756
rect 18172 42702 18174 42754
rect 18226 42702 18564 42754
rect 18172 42700 18564 42702
rect 18172 42690 18228 42700
rect 18060 42578 18116 42588
rect 17948 42364 18228 42420
rect 17836 42130 17892 42140
rect 18060 41524 18116 41534
rect 18172 41524 18228 42364
rect 18396 42082 18452 42094
rect 18396 42030 18398 42082
rect 18450 42030 18452 42082
rect 18116 41468 18228 41524
rect 18284 41970 18340 41982
rect 18284 41918 18286 41970
rect 18338 41918 18340 41970
rect 18060 41458 18116 41468
rect 18284 41188 18340 41918
rect 17500 40402 17668 40404
rect 17500 40350 17502 40402
rect 17554 40350 17668 40402
rect 17500 40348 17668 40350
rect 17500 40338 17556 40348
rect 17388 39394 17444 40124
rect 17500 39620 17556 39630
rect 17500 39526 17556 39564
rect 17388 39342 17390 39394
rect 17442 39342 17444 39394
rect 17388 39330 17444 39342
rect 16828 38836 16884 38846
rect 16716 38780 16828 38836
rect 16828 38770 16884 38780
rect 16716 38276 16772 38286
rect 16716 38274 16884 38276
rect 16716 38222 16718 38274
rect 16770 38222 16884 38274
rect 16716 38220 16884 38222
rect 16716 38210 16772 38220
rect 16604 38164 16660 38174
rect 16604 38070 16660 38108
rect 16828 37380 16884 38220
rect 17612 38052 17668 40348
rect 17948 40514 18004 40526
rect 17948 40462 17950 40514
rect 18002 40462 18004 40514
rect 17724 39732 17780 39742
rect 17724 39638 17780 39676
rect 17612 37986 17668 37996
rect 17724 38724 17780 38734
rect 17052 37940 17108 37950
rect 17052 37846 17108 37884
rect 16828 37268 16884 37324
rect 17276 37268 17332 37278
rect 17388 37268 17444 37278
rect 16828 37212 16996 37268
rect 16380 37174 16436 37212
rect 16268 37044 16324 37100
rect 16716 37154 16772 37166
rect 16716 37102 16718 37154
rect 16770 37102 16772 37154
rect 16716 37044 16772 37102
rect 16268 36988 16772 37044
rect 16156 36654 16158 36706
rect 16210 36654 16212 36706
rect 16156 36642 16212 36654
rect 16940 36706 16996 37212
rect 17332 37266 17444 37268
rect 17332 37214 17390 37266
rect 17442 37214 17444 37266
rect 17332 37212 17444 37214
rect 16940 36654 16942 36706
rect 16994 36654 16996 36706
rect 16940 36642 16996 36654
rect 17164 36932 17220 36942
rect 15708 35196 15876 35252
rect 15932 36594 15988 36606
rect 15932 36542 15934 36594
rect 15986 36542 15988 36594
rect 15932 36484 15988 36542
rect 15932 35474 15988 36428
rect 16828 36594 16884 36606
rect 16828 36542 16830 36594
rect 16882 36542 16884 36594
rect 16828 36484 16884 36542
rect 16828 36418 16884 36428
rect 17164 36482 17220 36876
rect 17164 36430 17166 36482
rect 17218 36430 17220 36482
rect 17164 36418 17220 36430
rect 15932 35422 15934 35474
rect 15986 35422 15988 35474
rect 14476 33966 14478 34018
rect 14530 33966 14532 34018
rect 14476 33954 14532 33966
rect 14812 34242 14868 34254
rect 14812 34190 14814 34242
rect 14866 34190 14868 34242
rect 14812 33684 14868 34190
rect 14812 33618 14868 33628
rect 13916 33406 13918 33458
rect 13970 33406 13972 33458
rect 13916 33394 13972 33406
rect 15148 33346 15204 33358
rect 15148 33294 15150 33346
rect 15202 33294 15204 33346
rect 14812 33124 14868 33134
rect 15148 33124 15204 33294
rect 14812 33122 15204 33124
rect 14812 33070 14814 33122
rect 14866 33070 15204 33122
rect 14812 33068 15204 33070
rect 14812 33058 14868 33068
rect 13916 31892 13972 31902
rect 13916 31780 13972 31836
rect 14252 31890 14308 31902
rect 14252 31838 14254 31890
rect 14306 31838 14308 31890
rect 14028 31780 14084 31790
rect 13916 31778 14084 31780
rect 13916 31726 14030 31778
rect 14082 31726 14084 31778
rect 13916 31724 14084 31726
rect 12796 28082 13188 28084
rect 12796 28030 12798 28082
rect 12850 28030 13188 28082
rect 12796 28028 13188 28030
rect 13468 29932 13748 29988
rect 13804 30212 13860 30222
rect 13916 30212 13972 31724
rect 14028 31714 14084 31724
rect 13804 30210 13972 30212
rect 13804 30158 13806 30210
rect 13858 30158 13972 30210
rect 13804 30156 13972 30158
rect 14140 31666 14196 31678
rect 14140 31614 14142 31666
rect 14194 31614 14196 31666
rect 14140 30210 14196 31614
rect 14140 30158 14142 30210
rect 14194 30158 14196 30210
rect 12796 28018 12852 28028
rect 12684 27806 12686 27858
rect 12738 27806 12740 27858
rect 12684 27794 12740 27806
rect 12908 27858 12964 27870
rect 12908 27806 12910 27858
rect 12962 27806 12964 27858
rect 12460 27186 12572 27188
rect 12460 27134 12462 27186
rect 12514 27134 12572 27186
rect 12460 27132 12572 27134
rect 12460 27122 12516 27132
rect 12572 27094 12628 27132
rect 12236 27076 12292 27086
rect 11788 26852 11956 26908
rect 10220 26514 10724 26516
rect 10220 26462 10670 26514
rect 10722 26462 10724 26514
rect 10220 26460 10724 26462
rect 10220 26290 10276 26460
rect 10668 26450 10724 26460
rect 10220 26238 10222 26290
rect 10274 26238 10276 26290
rect 10220 26226 10276 26238
rect 11788 26292 11844 26302
rect 11900 26292 11956 26852
rect 11788 26290 11956 26292
rect 11788 26238 11790 26290
rect 11842 26238 11956 26290
rect 11788 26236 11956 26238
rect 9996 25284 10052 25452
rect 11004 26180 11060 26190
rect 9996 25228 10164 25284
rect 8988 24894 8990 24946
rect 9042 24894 9044 24946
rect 8988 24882 9044 24894
rect 10108 24722 10164 25228
rect 10108 24670 10110 24722
rect 10162 24670 10164 24722
rect 10108 24658 10164 24670
rect 10780 24612 10836 24622
rect 10780 24518 10836 24556
rect 11004 16324 11060 26124
rect 11788 25620 11844 26236
rect 12236 26178 12292 27020
rect 12236 26126 12238 26178
rect 12290 26126 12292 26178
rect 12236 26114 12292 26126
rect 12908 27074 12964 27806
rect 13468 27748 13524 29932
rect 13804 29764 13860 30156
rect 13468 27682 13524 27692
rect 13580 29708 13860 29764
rect 13916 29988 13972 29998
rect 12908 27022 12910 27074
rect 12962 27022 12964 27074
rect 11788 25554 11844 25564
rect 12236 25508 12292 25518
rect 12236 25414 12292 25452
rect 12796 25508 12852 25518
rect 12796 25414 12852 25452
rect 11564 25396 11620 25406
rect 11564 25302 11620 25340
rect 12908 24610 12964 27022
rect 13580 27076 13636 29708
rect 13916 29314 13972 29932
rect 13916 29262 13918 29314
rect 13970 29262 13972 29314
rect 13916 29250 13972 29262
rect 14140 28980 14196 30158
rect 14252 31668 14308 31838
rect 14252 29426 14308 31612
rect 15036 31890 15092 33068
rect 15036 31838 15038 31890
rect 15090 31838 15092 31890
rect 15036 31780 15092 31838
rect 15372 31780 15428 31790
rect 15036 31778 15428 31780
rect 15036 31726 15374 31778
rect 15426 31726 15428 31778
rect 15036 31724 15428 31726
rect 15036 31444 15092 31724
rect 15372 31714 15428 31724
rect 15036 31378 15092 31388
rect 14812 30212 14868 30222
rect 14812 30118 14868 30156
rect 15708 30212 15764 35196
rect 15820 35028 15876 35038
rect 15932 35028 15988 35422
rect 15820 35026 15988 35028
rect 15820 34974 15822 35026
rect 15874 34974 15988 35026
rect 15820 34972 15988 34974
rect 16156 35700 16212 35710
rect 15820 34962 15876 34972
rect 16156 34132 16212 35644
rect 17276 35138 17332 37212
rect 17388 37202 17444 37212
rect 17724 36708 17780 38668
rect 17948 38724 18004 40462
rect 18060 38836 18116 38846
rect 18060 38742 18116 38780
rect 18284 38668 18340 41132
rect 18396 40404 18452 42030
rect 18396 40338 18452 40348
rect 18508 39956 18564 42700
rect 19404 42754 19460 42766
rect 19404 42702 19406 42754
rect 19458 42702 19460 42754
rect 19404 41860 19460 42702
rect 20300 42644 20356 42654
rect 20300 42550 20356 42588
rect 20524 42530 20580 42542
rect 20524 42478 20526 42530
rect 20578 42478 20580 42530
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20524 42308 20580 42478
rect 19836 42298 20100 42308
rect 20300 42252 20580 42308
rect 19852 41972 19908 41982
rect 20300 41972 20356 42252
rect 20636 42196 20692 43596
rect 20972 43540 21028 44268
rect 21644 44324 21700 45054
rect 21644 44258 21700 44268
rect 21756 45218 21812 45230
rect 21756 45166 21758 45218
rect 21810 45166 21812 45218
rect 21756 45108 21812 45166
rect 22204 45220 22260 45230
rect 23100 45220 23156 45614
rect 23212 45332 23268 45342
rect 23268 45276 23380 45332
rect 23212 45266 23268 45276
rect 22204 45126 22260 45164
rect 22876 45164 23156 45220
rect 21756 44322 21812 45052
rect 21980 45106 22036 45118
rect 21980 45054 21982 45106
rect 22034 45054 22036 45106
rect 21980 44996 22036 45054
rect 22428 45108 22484 45118
rect 22428 45014 22484 45052
rect 22876 45106 22932 45164
rect 22876 45054 22878 45106
rect 22930 45054 22932 45106
rect 22316 44996 22372 45006
rect 21980 44940 22316 44996
rect 22316 44930 22372 44940
rect 21756 44270 21758 44322
rect 21810 44270 21812 44322
rect 21756 43708 21812 44270
rect 22092 44324 22148 44334
rect 22092 44230 22148 44268
rect 22316 44212 22372 44222
rect 22652 44212 22708 44222
rect 22204 44210 22708 44212
rect 22204 44158 22318 44210
rect 22370 44158 22654 44210
rect 22706 44158 22708 44210
rect 22204 44156 22708 44158
rect 21756 43652 21924 43708
rect 20972 43474 21028 43484
rect 21868 43426 21924 43652
rect 22204 43650 22260 44156
rect 22316 44146 22372 44156
rect 22652 44146 22708 44156
rect 22764 44098 22820 44110
rect 22764 44046 22766 44098
rect 22818 44046 22820 44098
rect 22204 43598 22206 43650
rect 22258 43598 22260 43650
rect 22204 43586 22260 43598
rect 22540 43988 22596 43998
rect 22540 43650 22596 43932
rect 22540 43598 22542 43650
rect 22594 43598 22596 43650
rect 22540 43586 22596 43598
rect 22764 43650 22820 44046
rect 22876 44098 22932 45054
rect 23324 45106 23380 45276
rect 23324 45054 23326 45106
rect 23378 45054 23380 45106
rect 23324 45042 23380 45054
rect 23100 44996 23156 45006
rect 23100 44902 23156 44940
rect 23436 44436 23492 48412
rect 23548 48354 23604 49084
rect 23660 49138 23716 49646
rect 23660 49086 23662 49138
rect 23714 49086 23716 49138
rect 23660 49074 23716 49086
rect 23548 48302 23550 48354
rect 23602 48302 23604 48354
rect 23548 48290 23604 48302
rect 23884 48132 23940 48142
rect 23884 48038 23940 48076
rect 23660 47460 23716 47470
rect 23660 47366 23716 47404
rect 23996 47346 24052 49756
rect 24444 49140 24500 49150
rect 24444 48468 24500 49084
rect 25116 49028 25172 50428
rect 25116 48962 25172 48972
rect 24444 48466 24836 48468
rect 24444 48414 24446 48466
rect 24498 48414 24836 48466
rect 24444 48412 24836 48414
rect 24444 48402 24500 48412
rect 24668 48132 24724 48142
rect 24668 48038 24724 48076
rect 24332 48018 24388 48030
rect 24332 47966 24334 48018
rect 24386 47966 24388 48018
rect 24332 47572 24388 47966
rect 24332 47506 24388 47516
rect 24556 47460 24612 47470
rect 24556 47366 24612 47404
rect 23996 47294 23998 47346
rect 24050 47294 24052 47346
rect 23996 47282 24052 47294
rect 24780 47346 24836 48412
rect 24780 47294 24782 47346
rect 24834 47294 24836 47346
rect 24780 47282 24836 47294
rect 24892 48132 24948 48142
rect 24892 47458 24948 48076
rect 24892 47406 24894 47458
rect 24946 47406 24948 47458
rect 24332 47236 24388 47246
rect 24332 47142 24388 47180
rect 24668 47236 24724 47246
rect 23660 47124 23716 47134
rect 23660 46786 23716 47068
rect 24556 46900 24612 46910
rect 24556 46806 24612 46844
rect 23660 46734 23662 46786
rect 23714 46734 23716 46786
rect 23660 46722 23716 46734
rect 23548 46676 23604 46686
rect 24444 46676 24500 46686
rect 23548 46582 23604 46620
rect 24108 46674 24500 46676
rect 24108 46622 24446 46674
rect 24498 46622 24500 46674
rect 24108 46620 24500 46622
rect 23660 46116 23716 46126
rect 23660 45330 23716 46060
rect 23660 45278 23662 45330
rect 23714 45278 23716 45330
rect 23660 45266 23716 45278
rect 24108 45330 24164 46620
rect 24444 46610 24500 46620
rect 24668 45668 24724 47180
rect 24892 47124 24948 47406
rect 24892 47058 24948 47068
rect 25452 47236 25508 47246
rect 25452 47012 25508 47180
rect 25452 46946 25508 46956
rect 24108 45278 24110 45330
rect 24162 45278 24164 45330
rect 24108 45266 24164 45278
rect 24332 45612 24724 45668
rect 25228 46676 25284 46686
rect 23324 44324 23380 44334
rect 23436 44324 23492 44380
rect 24108 44436 24164 44446
rect 24108 44342 24164 44380
rect 22876 44046 22878 44098
rect 22930 44046 22932 44098
rect 22876 43988 22932 44046
rect 22876 43922 22932 43932
rect 23100 44322 23492 44324
rect 23100 44270 23326 44322
rect 23378 44270 23492 44322
rect 23100 44268 23492 44270
rect 22764 43598 22766 43650
rect 22818 43598 22820 43650
rect 22764 43586 22820 43598
rect 21868 43374 21870 43426
rect 21922 43374 21924 43426
rect 21868 43362 21924 43374
rect 22316 43428 22372 43438
rect 22316 43334 22372 43372
rect 20860 43204 20916 43214
rect 20524 42140 20692 42196
rect 20748 42642 20804 42654
rect 20748 42590 20750 42642
rect 20802 42590 20804 42642
rect 20524 42084 20580 42140
rect 19852 41970 20244 41972
rect 19852 41918 19854 41970
rect 19906 41918 20244 41970
rect 19852 41916 20244 41918
rect 19852 41906 19908 41916
rect 19068 41186 19124 41198
rect 19068 41134 19070 41186
rect 19122 41134 19124 41186
rect 17948 38658 18004 38668
rect 18172 38612 18340 38668
rect 18396 39900 18564 39956
rect 18844 41074 18900 41086
rect 18844 41022 18846 41074
rect 18898 41022 18900 41074
rect 17948 38164 18004 38174
rect 17948 37266 18004 38108
rect 18172 37380 18228 38612
rect 18284 37380 18340 37390
rect 18172 37378 18340 37380
rect 18172 37326 18286 37378
rect 18338 37326 18340 37378
rect 18172 37324 18340 37326
rect 17948 37214 17950 37266
rect 18002 37214 18004 37266
rect 17948 37202 18004 37214
rect 17612 36652 17780 36708
rect 17500 36482 17556 36494
rect 17500 36430 17502 36482
rect 17554 36430 17556 36482
rect 17500 35476 17556 36430
rect 17500 35410 17556 35420
rect 17276 35086 17278 35138
rect 17330 35086 17332 35138
rect 17276 35074 17332 35086
rect 16268 34916 16324 34926
rect 16604 34916 16660 34926
rect 16268 34914 16604 34916
rect 16268 34862 16270 34914
rect 16322 34862 16604 34914
rect 16268 34860 16604 34862
rect 16268 34850 16324 34860
rect 16604 34822 16660 34860
rect 16828 34914 16884 34926
rect 16828 34862 16830 34914
rect 16882 34862 16884 34914
rect 16828 34132 16884 34862
rect 15708 30146 15764 30156
rect 15820 34076 16884 34132
rect 17612 34132 17668 36652
rect 17948 36484 18004 36494
rect 17948 35810 18004 36428
rect 17948 35758 17950 35810
rect 18002 35758 18004 35810
rect 17948 35746 18004 35758
rect 15596 29988 15652 29998
rect 15372 29652 15428 29662
rect 14812 29538 14868 29550
rect 14812 29486 14814 29538
rect 14866 29486 14868 29538
rect 14588 29428 14644 29438
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 14252 29362 14308 29374
rect 14364 29426 14644 29428
rect 14364 29374 14590 29426
rect 14642 29374 14644 29426
rect 14364 29372 14644 29374
rect 14140 28914 14196 28924
rect 14364 28756 14420 29372
rect 14588 29362 14644 29372
rect 14700 29316 14756 29326
rect 14700 29222 14756 29260
rect 14812 29092 14868 29486
rect 14812 29026 14868 29036
rect 15036 29426 15092 29438
rect 15036 29374 15038 29426
rect 15090 29374 15092 29426
rect 13916 28700 14420 28756
rect 13916 28644 13972 28700
rect 13580 27010 13636 27020
rect 13692 28642 13972 28644
rect 13692 28590 13918 28642
rect 13970 28590 13972 28642
rect 13692 28588 13972 28590
rect 13468 26964 13524 27002
rect 13468 26898 13524 26908
rect 13692 26404 13748 28588
rect 13916 28578 13972 28588
rect 14700 28644 14756 28654
rect 14700 28550 14756 28588
rect 14140 28532 14196 28542
rect 14140 28438 14196 28476
rect 14252 28530 14308 28542
rect 14252 28478 14254 28530
rect 14306 28478 14308 28530
rect 14028 28420 14084 28430
rect 14028 28326 14084 28364
rect 14140 28084 14196 28094
rect 14252 28084 14308 28478
rect 14140 28082 14308 28084
rect 14140 28030 14142 28082
rect 14194 28030 14308 28082
rect 14140 28028 14308 28030
rect 14924 28308 14980 28318
rect 14924 28082 14980 28252
rect 14924 28030 14926 28082
rect 14978 28030 14980 28082
rect 14140 28018 14196 28028
rect 14924 28018 14980 28030
rect 14364 27970 14420 27982
rect 14364 27918 14366 27970
rect 14418 27918 14420 27970
rect 14364 27748 14420 27918
rect 14364 27682 14420 27692
rect 14476 27860 14532 27870
rect 14812 27860 14868 27870
rect 14476 27858 14868 27860
rect 14476 27806 14478 27858
rect 14530 27806 14814 27858
rect 14866 27806 14868 27858
rect 14476 27804 14868 27806
rect 14476 27300 14532 27804
rect 14140 27244 14532 27300
rect 14140 27076 14196 27244
rect 14588 27188 14644 27198
rect 14644 27132 14756 27188
rect 14588 27122 14644 27132
rect 13804 27074 14196 27076
rect 13804 27022 14142 27074
rect 14194 27022 14196 27074
rect 13804 27020 14196 27022
rect 13804 26962 13860 27020
rect 14140 27010 14196 27020
rect 14252 27076 14308 27086
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13804 26898 13860 26910
rect 14252 26962 14308 27020
rect 14252 26910 14254 26962
rect 14306 26910 14308 26962
rect 14252 26898 14308 26910
rect 14700 26908 14756 27132
rect 14812 27076 14868 27804
rect 14924 27636 14980 27646
rect 15036 27636 15092 29374
rect 15372 29426 15428 29596
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15372 29362 15428 29374
rect 15596 29092 15652 29932
rect 15596 29026 15652 29036
rect 14924 27634 15092 27636
rect 14924 27582 14926 27634
rect 14978 27582 15092 27634
rect 14924 27580 15092 27582
rect 15148 28642 15204 28654
rect 15148 28590 15150 28642
rect 15202 28590 15204 28642
rect 15148 28532 15204 28590
rect 14924 27570 14980 27580
rect 15148 27524 15204 28476
rect 15148 27458 15204 27468
rect 14924 27076 14980 27086
rect 14812 27074 14980 27076
rect 14812 27022 14926 27074
rect 14978 27022 14980 27074
rect 14812 27020 14980 27022
rect 14924 27010 14980 27020
rect 14476 26852 14532 26862
rect 13244 26290 13300 26302
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 25620 13300 26238
rect 13244 25554 13300 25564
rect 13356 25508 13412 25518
rect 13356 24946 13412 25452
rect 13692 25284 13748 26348
rect 14364 26850 14532 26852
rect 14364 26798 14478 26850
rect 14530 26798 14532 26850
rect 14364 26796 14532 26798
rect 13916 26178 13972 26190
rect 13916 26126 13918 26178
rect 13970 26126 13972 26178
rect 13916 25508 13972 26126
rect 14364 26068 14420 26796
rect 14476 26786 14532 26796
rect 14588 26850 14644 26862
rect 14700 26852 14868 26908
rect 14588 26798 14590 26850
rect 14642 26798 14644 26850
rect 13916 25442 13972 25452
rect 14252 26012 14420 26068
rect 14476 26628 14532 26638
rect 14028 25396 14084 25406
rect 14028 25302 14084 25340
rect 14252 25394 14308 26012
rect 14252 25342 14254 25394
rect 14306 25342 14308 25394
rect 14252 25330 14308 25342
rect 14476 25394 14532 26572
rect 14476 25342 14478 25394
rect 14530 25342 14532 25394
rect 13916 25284 13972 25294
rect 13692 25282 13972 25284
rect 13692 25230 13918 25282
rect 13970 25230 13972 25282
rect 13692 25228 13972 25230
rect 13356 24894 13358 24946
rect 13410 24894 13412 24946
rect 13356 24882 13412 24894
rect 13916 24946 13972 25228
rect 14140 25282 14196 25294
rect 14140 25230 14142 25282
rect 14194 25230 14196 25282
rect 14140 25172 14196 25230
rect 14140 25106 14196 25116
rect 13916 24894 13918 24946
rect 13970 24894 13972 24946
rect 13916 24882 13972 24894
rect 14140 24836 14196 24846
rect 14140 24834 14308 24836
rect 14140 24782 14142 24834
rect 14194 24782 14308 24834
rect 14140 24780 14308 24782
rect 14140 24770 14196 24780
rect 12908 24558 12910 24610
rect 12962 24558 12964 24610
rect 12908 24546 12964 24558
rect 13916 24724 13972 24734
rect 13916 23042 13972 24668
rect 14028 24612 14084 24622
rect 14028 24518 14084 24556
rect 14252 24612 14308 24780
rect 14476 24834 14532 25342
rect 14476 24782 14478 24834
rect 14530 24782 14532 24834
rect 14476 24770 14532 24782
rect 14364 24722 14420 24734
rect 14364 24670 14366 24722
rect 14418 24670 14420 24722
rect 14364 24612 14420 24670
rect 14588 24612 14644 26798
rect 14812 26850 14868 26852
rect 14812 26798 14814 26850
rect 14866 26798 14868 26850
rect 14812 26786 14868 26798
rect 15596 26404 15652 26414
rect 15596 26310 15652 26348
rect 15484 25956 15540 25966
rect 15484 25620 15540 25900
rect 15484 25526 15540 25564
rect 14364 24556 14644 24612
rect 14700 25508 14756 25518
rect 14252 24546 14308 24556
rect 13916 22990 13918 23042
rect 13970 22990 13972 23042
rect 13916 22978 13972 22990
rect 14700 20916 14756 25452
rect 15148 25172 15204 25182
rect 15148 24946 15204 25116
rect 15148 24894 15150 24946
rect 15202 24894 15204 24946
rect 15148 24882 15204 24894
rect 15820 24724 15876 34076
rect 17612 34066 17668 34076
rect 17836 34916 17892 34926
rect 17836 34130 17892 34860
rect 17948 34804 18004 34814
rect 18004 34748 18116 34804
rect 17948 34710 18004 34748
rect 17836 34078 17838 34130
rect 17890 34078 17892 34130
rect 17836 34066 17892 34078
rect 18060 33458 18116 34748
rect 18284 34692 18340 37324
rect 18396 37154 18452 39900
rect 18844 39732 18900 41022
rect 18844 39638 18900 39676
rect 18956 41076 19012 41086
rect 18956 39618 19012 41020
rect 18956 39566 18958 39618
rect 19010 39566 19012 39618
rect 18956 39172 19012 39566
rect 18732 39116 19012 39172
rect 19068 39620 19124 41134
rect 19404 40626 19460 41804
rect 19964 41748 20020 41758
rect 19964 41654 20020 41692
rect 20076 41300 20132 41310
rect 20076 41206 20132 41244
rect 19852 41188 19908 41198
rect 19852 41094 19908 41132
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19404 40574 19406 40626
rect 19458 40574 19460 40626
rect 19404 40562 19460 40574
rect 20188 40628 20244 41916
rect 20300 41906 20356 41916
rect 20412 42082 20580 42084
rect 20412 42030 20526 42082
rect 20578 42030 20580 42082
rect 20412 42028 20580 42030
rect 20300 41074 20356 41086
rect 20300 41022 20302 41074
rect 20354 41022 20356 41074
rect 20300 40852 20356 41022
rect 20412 40852 20468 42028
rect 20524 42018 20580 42028
rect 20636 41970 20692 41982
rect 20636 41918 20638 41970
rect 20690 41918 20692 41970
rect 20524 41076 20580 41086
rect 20524 40982 20580 41020
rect 20412 40796 20580 40852
rect 20300 40786 20356 40796
rect 20412 40628 20468 40638
rect 20188 40626 20468 40628
rect 20188 40574 20414 40626
rect 20466 40574 20468 40626
rect 20188 40572 20468 40574
rect 18508 38834 18564 38846
rect 18508 38782 18510 38834
rect 18562 38782 18564 38834
rect 18508 38612 18564 38782
rect 18620 38724 18676 38734
rect 18732 38724 18788 39116
rect 18844 38948 18900 38958
rect 18844 38834 18900 38892
rect 18844 38782 18846 38834
rect 18898 38782 18900 38834
rect 18844 38770 18900 38782
rect 18676 38668 18788 38724
rect 18620 38630 18676 38668
rect 18508 38276 18564 38556
rect 18956 38276 19012 38286
rect 18508 38220 18676 38276
rect 18620 38164 18676 38220
rect 18844 38220 18956 38276
rect 18620 38162 18788 38164
rect 18620 38110 18622 38162
rect 18674 38110 18788 38162
rect 18620 38108 18788 38110
rect 18620 38098 18676 38108
rect 18396 37102 18398 37154
rect 18450 37102 18452 37154
rect 18396 37090 18452 37102
rect 18508 38052 18564 38062
rect 18508 37156 18564 37996
rect 18508 37090 18564 37100
rect 18620 37828 18676 37838
rect 18508 36596 18564 36606
rect 18620 36596 18676 37772
rect 18508 36594 18676 36596
rect 18508 36542 18510 36594
rect 18562 36542 18676 36594
rect 18508 36540 18676 36542
rect 18508 36530 18564 36540
rect 18508 34804 18564 34814
rect 18564 34748 18676 34804
rect 18508 34710 18564 34748
rect 18060 33406 18062 33458
rect 18114 33406 18116 33458
rect 18060 33394 18116 33406
rect 18172 34636 18340 34692
rect 15932 33236 15988 33246
rect 15932 33142 15988 33180
rect 17948 32004 18004 32014
rect 17500 31892 17556 31902
rect 16156 31668 16212 31678
rect 16156 31666 16436 31668
rect 16156 31614 16158 31666
rect 16210 31614 16436 31666
rect 16156 31612 16436 31614
rect 16156 31602 16212 31612
rect 16268 30212 16324 30222
rect 16044 29428 16100 29438
rect 16044 29334 16100 29372
rect 15932 28756 15988 28766
rect 16268 28756 16324 30156
rect 16380 29316 16436 31612
rect 16716 31444 16772 31454
rect 16604 29988 16660 29998
rect 16604 29650 16660 29932
rect 16604 29598 16606 29650
rect 16658 29598 16660 29650
rect 16604 29586 16660 29598
rect 16492 29540 16548 29550
rect 16492 29446 16548 29484
rect 16492 29316 16548 29326
rect 16380 29314 16548 29316
rect 16380 29262 16494 29314
rect 16546 29262 16548 29314
rect 16380 29260 16548 29262
rect 16492 29250 16548 29260
rect 15932 28754 16324 28756
rect 15932 28702 15934 28754
rect 15986 28702 16324 28754
rect 15932 28700 16324 28702
rect 15932 28690 15988 28700
rect 16156 28532 16212 28542
rect 16156 28438 16212 28476
rect 16268 28530 16324 28700
rect 16716 28644 16772 31388
rect 17500 29650 17556 31836
rect 17948 29764 18004 31948
rect 18172 31668 18228 34636
rect 18620 34354 18676 34748
rect 18620 34302 18622 34354
rect 18674 34302 18676 34354
rect 18620 34290 18676 34302
rect 18284 34132 18340 34142
rect 18284 34038 18340 34076
rect 18508 33234 18564 33246
rect 18508 33182 18510 33234
rect 18562 33182 18564 33234
rect 18508 33124 18564 33182
rect 18620 33236 18676 33246
rect 18620 33142 18676 33180
rect 18508 33058 18564 33068
rect 18732 32786 18788 38108
rect 18844 37156 18900 38220
rect 18956 38210 19012 38220
rect 19068 38274 19124 39564
rect 19180 40516 19236 40526
rect 19180 40290 19236 40460
rect 19180 40238 19182 40290
rect 19234 40238 19236 40290
rect 19180 38668 19236 40238
rect 19292 39618 19348 39630
rect 19292 39566 19294 39618
rect 19346 39566 19348 39618
rect 19292 38948 19348 39566
rect 20188 39620 20244 40572
rect 20412 40562 20468 40572
rect 20300 40404 20356 40414
rect 20524 40404 20580 40796
rect 20300 40310 20356 40348
rect 20412 40348 20580 40404
rect 20412 40178 20468 40348
rect 20412 40126 20414 40178
rect 20466 40126 20468 40178
rect 20412 40114 20468 40126
rect 20188 39554 20244 39564
rect 20188 39394 20244 39406
rect 20188 39342 20190 39394
rect 20242 39342 20244 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19292 38882 19348 38892
rect 19852 38946 19908 38958
rect 19852 38894 19854 38946
rect 19906 38894 19908 38946
rect 19180 38612 19348 38668
rect 19068 38222 19070 38274
rect 19122 38222 19124 38274
rect 19068 38210 19124 38222
rect 18956 37940 19012 37950
rect 18956 37378 19012 37884
rect 18956 37326 18958 37378
rect 19010 37326 19012 37378
rect 18956 37314 19012 37326
rect 19068 37268 19124 37278
rect 18844 37100 19012 37156
rect 18844 36482 18900 36494
rect 18844 36430 18846 36482
rect 18898 36430 18900 36482
rect 18844 36372 18900 36430
rect 18844 35698 18900 36316
rect 18956 35922 19012 37100
rect 18956 35870 18958 35922
rect 19010 35870 19012 35922
rect 18956 35858 19012 35870
rect 19068 36370 19124 37212
rect 19068 36318 19070 36370
rect 19122 36318 19124 36370
rect 18844 35646 18846 35698
rect 18898 35646 18900 35698
rect 18844 33572 18900 35646
rect 19068 35026 19124 36318
rect 19068 34974 19070 35026
rect 19122 34974 19124 35026
rect 19068 34962 19124 34974
rect 19180 35586 19236 35598
rect 19180 35534 19182 35586
rect 19234 35534 19236 35586
rect 19180 35476 19236 35534
rect 19180 34356 19236 35420
rect 19068 34300 19236 34356
rect 19068 33908 19124 34300
rect 19180 34132 19236 34142
rect 19180 34038 19236 34076
rect 19068 33852 19236 33908
rect 18844 33516 19012 33572
rect 18844 33348 18900 33358
rect 18844 33254 18900 33292
rect 18732 32734 18734 32786
rect 18786 32734 18788 32786
rect 18732 32722 18788 32734
rect 18620 32450 18676 32462
rect 18620 32398 18622 32450
rect 18674 32398 18676 32450
rect 18284 31892 18340 31902
rect 18620 31892 18676 32398
rect 18284 31890 18676 31892
rect 18284 31838 18286 31890
rect 18338 31838 18676 31890
rect 18284 31836 18676 31838
rect 18284 31826 18340 31836
rect 18620 31778 18676 31836
rect 18956 31892 19012 33516
rect 19068 33234 19124 33246
rect 19068 33182 19070 33234
rect 19122 33182 19124 33234
rect 19068 33012 19124 33182
rect 19068 32946 19124 32956
rect 19068 31892 19124 31902
rect 19012 31890 19124 31892
rect 19012 31838 19070 31890
rect 19122 31838 19124 31890
rect 19012 31836 19124 31838
rect 18956 31798 19012 31836
rect 19068 31826 19124 31836
rect 18620 31726 18622 31778
rect 18674 31726 18676 31778
rect 18620 31714 18676 31726
rect 19180 31668 19236 33852
rect 18172 31612 18340 31668
rect 17948 29698 18004 29708
rect 18060 29988 18116 29998
rect 17500 29598 17502 29650
rect 17554 29598 17556 29650
rect 17500 29586 17556 29598
rect 18060 29650 18116 29932
rect 18060 29598 18062 29650
rect 18114 29598 18116 29650
rect 18060 29586 18116 29598
rect 17276 29540 17332 29550
rect 17276 29446 17332 29484
rect 16828 29428 16884 29438
rect 16828 29426 17220 29428
rect 16828 29374 16830 29426
rect 16882 29374 17220 29426
rect 16828 29372 17220 29374
rect 16828 29362 16884 29372
rect 16828 28644 16884 28654
rect 16268 28478 16270 28530
rect 16322 28478 16324 28530
rect 16268 28466 16324 28478
rect 16380 28642 16884 28644
rect 16380 28590 16830 28642
rect 16882 28590 16884 28642
rect 16380 28588 16884 28590
rect 16380 28082 16436 28588
rect 16828 28578 16884 28588
rect 16492 28420 16548 28430
rect 16492 28326 16548 28364
rect 16380 28030 16382 28082
rect 16434 28030 16436 28082
rect 16380 26908 16436 28030
rect 17164 28084 17220 29372
rect 17612 29426 17668 29438
rect 17612 29374 17614 29426
rect 17666 29374 17668 29426
rect 17612 28644 17668 29374
rect 17612 28588 17892 28644
rect 17500 28530 17556 28542
rect 17500 28478 17502 28530
rect 17554 28478 17556 28530
rect 17388 28084 17444 28094
rect 17164 28082 17444 28084
rect 17164 28030 17390 28082
rect 17442 28030 17444 28082
rect 17164 28028 17444 28030
rect 17164 26908 17220 28028
rect 17388 28018 17444 28028
rect 17500 28082 17556 28478
rect 17612 28532 17668 28588
rect 17612 28466 17668 28476
rect 17500 28030 17502 28082
rect 17554 28030 17556 28082
rect 17500 28018 17556 28030
rect 17724 28420 17780 28430
rect 17612 27972 17668 27982
rect 17612 27878 17668 27916
rect 17724 27970 17780 28364
rect 17724 27918 17726 27970
rect 17778 27918 17780 27970
rect 17724 27906 17780 27918
rect 17836 27748 17892 28588
rect 17724 27692 17892 27748
rect 18172 27858 18228 27870
rect 18172 27806 18174 27858
rect 18226 27806 18228 27858
rect 17724 26908 17780 27692
rect 18172 27636 18228 27806
rect 15932 26852 15988 26862
rect 15932 26404 15988 26796
rect 15932 26310 15988 26348
rect 16044 26852 16436 26908
rect 16492 26852 17220 26908
rect 17388 26852 17780 26908
rect 17836 27524 17892 27534
rect 15932 25620 15988 25630
rect 16044 25620 16100 26852
rect 16492 26514 16548 26852
rect 16492 26462 16494 26514
rect 16546 26462 16548 26514
rect 16492 26450 16548 26462
rect 15988 25564 16100 25620
rect 15932 25526 15988 25564
rect 16268 25508 16324 25518
rect 16268 25414 16324 25452
rect 16380 25282 16436 25294
rect 16604 25284 16660 25294
rect 16380 25230 16382 25282
rect 16434 25230 16436 25282
rect 16044 24948 16100 24958
rect 16044 24854 16100 24892
rect 15820 24658 15876 24668
rect 16268 24834 16324 24846
rect 16268 24782 16270 24834
rect 16322 24782 16324 24834
rect 15596 24612 15652 24622
rect 15596 24518 15652 24556
rect 16156 24610 16212 24622
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 16044 23268 16100 23278
rect 16156 23268 16212 24558
rect 16268 24612 16324 24782
rect 16380 24724 16436 25230
rect 16380 24658 16436 24668
rect 16492 25282 16660 25284
rect 16492 25230 16606 25282
rect 16658 25230 16660 25282
rect 16492 25228 16660 25230
rect 16492 24722 16548 25228
rect 16604 25218 16660 25228
rect 16716 24948 16772 26852
rect 17388 26402 17444 26852
rect 17388 26350 17390 26402
rect 17442 26350 17444 26402
rect 16828 26290 16884 26302
rect 16828 26238 16830 26290
rect 16882 26238 16884 26290
rect 16828 26180 16884 26238
rect 16828 26114 16884 26124
rect 17388 26292 17444 26350
rect 16716 24882 16772 24892
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 16492 24658 16548 24670
rect 16716 24722 16772 24734
rect 16716 24670 16718 24722
rect 16770 24670 16772 24722
rect 16268 23828 16324 24556
rect 16716 24500 16772 24670
rect 16716 24434 16772 24444
rect 16268 23762 16324 23772
rect 16044 23266 16212 23268
rect 16044 23214 16046 23266
rect 16098 23214 16212 23266
rect 16044 23212 16212 23214
rect 16044 23202 16100 23212
rect 16828 23156 16884 25454
rect 17388 25508 17444 26236
rect 17388 25442 17444 25452
rect 17724 26290 17780 26302
rect 17724 26238 17726 26290
rect 17778 26238 17780 26290
rect 17724 26180 17780 26238
rect 17724 25508 17780 26124
rect 17724 25442 17780 25452
rect 17612 25396 17668 25406
rect 17500 25394 17668 25396
rect 17500 25342 17614 25394
rect 17666 25342 17668 25394
rect 17500 25340 17668 25342
rect 17388 24948 17444 24958
rect 17388 24854 17444 24892
rect 17500 24946 17556 25340
rect 17612 25330 17668 25340
rect 17836 25284 17892 27468
rect 18172 27186 18228 27580
rect 18172 27134 18174 27186
rect 18226 27134 18228 27186
rect 18172 27122 18228 27134
rect 18172 26404 18228 26414
rect 18284 26404 18340 31612
rect 19068 31612 19236 31668
rect 18844 29428 18900 29438
rect 18844 28082 18900 29372
rect 18844 28030 18846 28082
rect 18898 28030 18900 28082
rect 18844 28018 18900 28030
rect 18620 27972 18676 27982
rect 18620 27186 18676 27916
rect 18620 27134 18622 27186
rect 18674 27134 18676 27186
rect 18620 26908 18676 27134
rect 18956 27636 19012 27646
rect 18620 26852 18788 26908
rect 18620 26404 18676 26414
rect 18172 26402 18676 26404
rect 18172 26350 18174 26402
rect 18226 26350 18622 26402
rect 18674 26350 18676 26402
rect 18172 26348 18676 26350
rect 18172 26338 18228 26348
rect 18620 26338 18676 26348
rect 18060 26292 18116 26302
rect 18060 26198 18116 26236
rect 17500 24894 17502 24946
rect 17554 24894 17556 24946
rect 17500 24882 17556 24894
rect 17724 25228 17892 25284
rect 18172 26066 18228 26078
rect 18172 26014 18174 26066
rect 18226 26014 18228 26066
rect 17612 24836 17668 24846
rect 17724 24836 17780 25228
rect 17668 24780 17780 24836
rect 18060 24948 18116 24958
rect 17612 24742 17668 24780
rect 17836 24724 17892 24734
rect 17836 24630 17892 24668
rect 18060 24722 18116 24892
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 17836 24500 17892 24510
rect 18060 24500 18116 24670
rect 18172 24724 18228 26014
rect 18732 25172 18788 26852
rect 18620 24836 18676 24846
rect 18620 24742 18676 24780
rect 18172 24658 18228 24668
rect 17892 24444 18116 24500
rect 17836 24050 17892 24444
rect 17836 23998 17838 24050
rect 17890 23998 17892 24050
rect 17836 23986 17892 23998
rect 17276 23828 17332 23838
rect 17276 23734 17332 23772
rect 18732 23716 18788 25116
rect 18956 24948 19012 27580
rect 19068 26908 19124 31612
rect 19180 30324 19236 30334
rect 19292 30324 19348 38612
rect 19852 38612 19908 38894
rect 19852 38546 19908 38556
rect 20188 38388 20244 39342
rect 20412 38948 20468 38958
rect 20412 38668 20468 38892
rect 20188 38322 20244 38332
rect 20300 38612 20468 38668
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37492 19684 37502
rect 19404 37380 19460 37390
rect 19404 34356 19460 37324
rect 19628 37266 19684 37436
rect 19628 37214 19630 37266
rect 19682 37214 19684 37266
rect 19516 35028 19572 35038
rect 19628 35028 19684 37214
rect 20188 37492 20244 37502
rect 19740 37156 19796 37166
rect 19740 37062 19796 37100
rect 20188 36482 20244 37436
rect 20300 36932 20356 38612
rect 20636 38276 20692 41918
rect 20748 41748 20804 42590
rect 20748 41682 20804 41692
rect 20748 40292 20804 40302
rect 20748 39730 20804 40236
rect 20748 39678 20750 39730
rect 20802 39678 20804 39730
rect 20748 39666 20804 39678
rect 20636 38210 20692 38220
rect 20748 38834 20804 38846
rect 20748 38782 20750 38834
rect 20802 38782 20804 38834
rect 20748 38052 20804 38782
rect 20860 38668 20916 43148
rect 22092 43204 22148 43214
rect 22092 42866 22148 43148
rect 22092 42814 22094 42866
rect 22146 42814 22148 42866
rect 22092 42802 22148 42814
rect 21420 42532 21476 42542
rect 21476 42476 21588 42532
rect 21420 42438 21476 42476
rect 20972 42196 21028 42206
rect 20972 42102 21028 42140
rect 21084 41972 21140 41982
rect 20972 40628 21028 40638
rect 20972 40534 21028 40572
rect 20972 38948 21028 38958
rect 21084 38948 21140 41916
rect 21420 41970 21476 41982
rect 21420 41918 21422 41970
rect 21474 41918 21476 41970
rect 21196 41860 21252 41870
rect 21196 41766 21252 41804
rect 21420 41636 21476 41918
rect 21420 41570 21476 41580
rect 21308 41524 21364 41534
rect 21308 41298 21364 41468
rect 21308 41246 21310 41298
rect 21362 41246 21364 41298
rect 21308 41234 21364 41246
rect 21420 40628 21476 40638
rect 21532 40628 21588 42476
rect 22652 42084 22708 42094
rect 21868 40964 21924 40974
rect 22316 40964 22372 40974
rect 21868 40962 22316 40964
rect 21868 40910 21870 40962
rect 21922 40910 22316 40962
rect 21868 40908 22316 40910
rect 21868 40898 21924 40908
rect 21476 40572 21588 40628
rect 21420 40534 21476 40572
rect 22204 39732 22260 39742
rect 22204 39638 22260 39676
rect 22316 39172 22372 40908
rect 22652 40516 22708 42028
rect 22988 40852 23044 40862
rect 22876 40516 22932 40526
rect 22540 40514 22932 40516
rect 22540 40462 22878 40514
rect 22930 40462 22932 40514
rect 22540 40460 22932 40462
rect 22428 39172 22484 39182
rect 22316 39116 22428 39172
rect 22428 39106 22484 39116
rect 20972 38946 21140 38948
rect 20972 38894 20974 38946
rect 21026 38894 21140 38946
rect 20972 38892 21140 38894
rect 20972 38882 21028 38892
rect 20860 38612 21028 38668
rect 20412 38050 20804 38052
rect 20412 37998 20750 38050
rect 20802 37998 20804 38050
rect 20412 37996 20804 37998
rect 20412 37268 20468 37996
rect 20748 37986 20804 37996
rect 20412 37174 20468 37212
rect 20860 37266 20916 37278
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 20748 37156 20804 37166
rect 20748 37062 20804 37100
rect 20356 36876 20804 36932
rect 20300 36838 20356 36876
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 20188 36418 20244 36430
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20300 35700 20356 35710
rect 19516 35026 19684 35028
rect 19516 34974 19518 35026
rect 19570 34974 19684 35026
rect 19516 34972 19684 34974
rect 19964 35698 20356 35700
rect 19964 35646 20302 35698
rect 20354 35646 20356 35698
rect 19964 35644 20356 35646
rect 19516 34962 19572 34972
rect 19964 34916 20020 35644
rect 20300 35634 20356 35644
rect 20748 35586 20804 36876
rect 20748 35534 20750 35586
rect 20802 35534 20804 35586
rect 20748 35522 20804 35534
rect 20860 35476 20916 37214
rect 20860 35410 20916 35420
rect 20860 35028 20916 35038
rect 20972 35028 21028 38612
rect 21308 38388 21364 38398
rect 21308 37938 21364 38332
rect 21308 37886 21310 37938
rect 21362 37886 21364 37938
rect 21308 37874 21364 37886
rect 21644 37828 21700 37838
rect 22204 37828 22260 37838
rect 21644 37826 22260 37828
rect 21644 37774 21646 37826
rect 21698 37774 22206 37826
rect 22258 37774 22260 37826
rect 21644 37772 22260 37774
rect 21308 36258 21364 36270
rect 21308 36206 21310 36258
rect 21362 36206 21364 36258
rect 21308 35588 21364 36206
rect 21644 36258 21700 37772
rect 22204 37762 22260 37772
rect 22540 36596 22596 40460
rect 22876 40450 22932 40460
rect 22988 40290 23044 40796
rect 23100 40740 23156 44268
rect 23324 44258 23380 44268
rect 23660 44098 23716 44110
rect 23660 44046 23662 44098
rect 23714 44046 23716 44098
rect 23212 43988 23268 43998
rect 23212 43762 23268 43932
rect 23660 43988 23716 44046
rect 23660 43922 23716 43932
rect 23212 43710 23214 43762
rect 23266 43710 23268 43762
rect 23212 43698 23268 43710
rect 23884 42082 23940 42094
rect 23884 42030 23886 42082
rect 23938 42030 23940 42082
rect 23548 41972 23604 41982
rect 23436 41970 23604 41972
rect 23436 41918 23550 41970
rect 23602 41918 23604 41970
rect 23436 41916 23604 41918
rect 23100 40674 23156 40684
rect 23212 41298 23268 41310
rect 23212 41246 23214 41298
rect 23266 41246 23268 41298
rect 22988 40238 22990 40290
rect 23042 40238 23044 40290
rect 22988 40226 23044 40238
rect 22652 40178 22708 40190
rect 22652 40126 22654 40178
rect 22706 40126 22708 40178
rect 22652 39620 22708 40126
rect 23212 39732 23268 41246
rect 23324 41186 23380 41198
rect 23324 41134 23326 41186
rect 23378 41134 23380 41186
rect 23324 40628 23380 41134
rect 23324 40562 23380 40572
rect 23436 40852 23492 41916
rect 23548 41906 23604 41916
rect 23772 41300 23828 41310
rect 23772 41206 23828 41244
rect 23884 40852 23940 42030
rect 23436 40402 23492 40796
rect 23436 40350 23438 40402
rect 23490 40350 23492 40402
rect 23436 40338 23492 40350
rect 23548 40796 23884 40852
rect 23436 39732 23492 39742
rect 23212 39676 23436 39732
rect 22652 39618 23380 39620
rect 22652 39566 22654 39618
rect 22706 39566 23380 39618
rect 22652 39564 23380 39566
rect 22652 39554 22708 39564
rect 23212 39172 23268 39182
rect 22988 37940 23044 37950
rect 22876 37156 22932 37166
rect 22876 37062 22932 37100
rect 22988 36708 23044 37884
rect 23100 36708 23156 36718
rect 22988 36706 23156 36708
rect 22988 36654 23102 36706
rect 23154 36654 23156 36706
rect 22988 36652 23156 36654
rect 23100 36642 23156 36652
rect 22540 36594 22708 36596
rect 22540 36542 22542 36594
rect 22594 36542 22708 36594
rect 22540 36540 22708 36542
rect 22540 36530 22596 36540
rect 21644 36206 21646 36258
rect 21698 36206 21700 36258
rect 21364 35532 21476 35588
rect 21308 35494 21364 35532
rect 20860 35026 21364 35028
rect 20860 34974 20862 35026
rect 20914 34974 21364 35026
rect 20860 34972 21364 34974
rect 20860 34962 20916 34972
rect 19628 34914 20020 34916
rect 19628 34862 19966 34914
rect 20018 34862 20020 34914
rect 19628 34860 20020 34862
rect 19404 34300 19572 34356
rect 19516 34132 19572 34300
rect 19516 33348 19572 34076
rect 19628 33572 19684 34860
rect 19964 34850 20020 34860
rect 21308 34914 21364 34972
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34850 21364 34862
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 21420 34244 21476 35532
rect 21308 34188 21476 34244
rect 19628 33516 19796 33572
rect 19628 33348 19684 33358
rect 19572 33346 19684 33348
rect 19572 33294 19630 33346
rect 19682 33294 19684 33346
rect 19572 33292 19684 33294
rect 19516 33282 19572 33292
rect 19628 33282 19684 33292
rect 19404 33124 19460 33134
rect 19404 32452 19460 33068
rect 19516 33122 19572 33134
rect 19740 33124 19796 33516
rect 20076 33348 20132 33358
rect 20076 33346 20244 33348
rect 20076 33294 20078 33346
rect 20130 33294 20244 33346
rect 20076 33292 20244 33294
rect 20076 33282 20132 33292
rect 19516 33070 19518 33122
rect 19570 33070 19572 33122
rect 19516 33012 19572 33070
rect 19516 32946 19572 32956
rect 19628 33068 19796 33124
rect 19404 32358 19460 32396
rect 19180 30322 19348 30324
rect 19180 30270 19182 30322
rect 19234 30270 19348 30322
rect 19180 30268 19348 30270
rect 19180 30212 19236 30268
rect 19180 30146 19236 30156
rect 19628 30210 19684 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32450 20244 33292
rect 20524 33124 20580 33134
rect 20524 33122 20804 33124
rect 20524 33070 20526 33122
rect 20578 33070 20804 33122
rect 20524 33068 20804 33070
rect 20524 33058 20580 33068
rect 20188 32398 20190 32450
rect 20242 32398 20244 32450
rect 20188 32340 20244 32398
rect 20188 32004 20244 32284
rect 20188 31938 20244 31948
rect 20748 32452 20804 33068
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 30884 20356 30894
rect 19628 30158 19630 30210
rect 19682 30158 19684 30210
rect 19628 28754 19684 30158
rect 20188 30828 20300 30884
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19628 28702 19630 28754
rect 19682 28702 19684 28754
rect 19628 28690 19684 28702
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19180 28084 19236 28094
rect 19180 27990 19236 28028
rect 19516 28084 19572 28094
rect 19516 27186 19572 28028
rect 19516 27134 19518 27186
rect 19570 27134 19572 27186
rect 19516 27122 19572 27134
rect 19628 27860 19684 27870
rect 19068 26852 19236 26908
rect 19180 26290 19236 26852
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 19180 25732 19236 26238
rect 19628 25844 19684 27804
rect 20188 27524 20244 30828
rect 20300 30818 20356 30828
rect 20748 30660 20804 32396
rect 21196 30884 21252 30894
rect 21196 30790 21252 30828
rect 20636 30604 20804 30660
rect 20412 29316 20468 29326
rect 20300 29260 20412 29316
rect 20300 27970 20356 29260
rect 20412 29250 20468 29260
rect 20300 27918 20302 27970
rect 20354 27918 20356 27970
rect 20300 27906 20356 27918
rect 20636 27524 20692 30604
rect 21308 29764 21364 34188
rect 21644 33460 21700 36206
rect 22092 34804 22148 34814
rect 21644 33394 21700 33404
rect 21868 34802 22148 34804
rect 21868 34750 22094 34802
rect 22146 34750 22148 34802
rect 21868 34748 22148 34750
rect 21420 33346 21476 33358
rect 21420 33294 21422 33346
rect 21474 33294 21476 33346
rect 21420 33124 21476 33294
rect 21420 33058 21476 33068
rect 21532 30996 21588 31006
rect 21420 30994 21588 30996
rect 21420 30942 21534 30994
rect 21586 30942 21588 30994
rect 21420 30940 21588 30942
rect 21420 30100 21476 30940
rect 21532 30930 21588 30940
rect 21868 30436 21924 34748
rect 22092 34738 22148 34748
rect 22092 33346 22148 33358
rect 22092 33294 22094 33346
rect 22146 33294 22148 33346
rect 22092 33236 22148 33294
rect 22204 33236 22260 33246
rect 22092 33180 22204 33236
rect 22204 33170 22260 33180
rect 21980 31106 22036 31118
rect 21980 31054 21982 31106
rect 22034 31054 22036 31106
rect 21980 30996 22036 31054
rect 21980 30930 22036 30940
rect 22092 31106 22148 31118
rect 22092 31054 22094 31106
rect 22146 31054 22148 31106
rect 22092 30884 22148 31054
rect 22204 31108 22260 31118
rect 22204 31014 22260 31052
rect 22092 30818 22148 30828
rect 22316 30994 22372 31006
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 22204 30436 22260 30446
rect 21532 30380 21924 30436
rect 21980 30380 22204 30436
rect 21532 30322 21588 30380
rect 21532 30270 21534 30322
rect 21586 30270 21588 30322
rect 21532 30258 21588 30270
rect 21868 30212 21924 30222
rect 21756 30100 21812 30110
rect 21420 30098 21812 30100
rect 21420 30046 21758 30098
rect 21810 30046 21812 30098
rect 21420 30044 21812 30046
rect 21308 29698 21364 29708
rect 21084 29652 21140 29662
rect 21084 29426 21140 29596
rect 21756 29652 21812 30044
rect 21756 29586 21812 29596
rect 21868 29650 21924 30156
rect 21980 30098 22036 30380
rect 22204 30370 22260 30380
rect 22316 30212 22372 30942
rect 22540 30996 22596 31006
rect 22540 30902 22596 30940
rect 22316 30118 22372 30156
rect 21980 30046 21982 30098
rect 22034 30046 22036 30098
rect 21980 30034 22036 30046
rect 22092 30098 22148 30110
rect 22092 30046 22094 30098
rect 22146 30046 22148 30098
rect 22092 29988 22148 30046
rect 22204 29988 22260 29998
rect 22092 29932 22204 29988
rect 22204 29922 22260 29932
rect 22652 29764 22708 36540
rect 22764 36482 22820 36494
rect 22764 36430 22766 36482
rect 22818 36430 22820 36482
rect 22764 35924 22820 36430
rect 22764 35858 22820 35868
rect 22764 35700 22820 35710
rect 22764 35606 22820 35644
rect 22764 33572 22820 33582
rect 22764 31218 22820 33516
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 31154 22820 31166
rect 22876 30996 22932 31006
rect 23100 30996 23156 31006
rect 22876 30902 22932 30940
rect 22988 30994 23156 30996
rect 22988 30942 23102 30994
rect 23154 30942 23156 30994
rect 22988 30940 23156 30942
rect 22988 30436 23044 30940
rect 23100 30930 23156 30940
rect 23212 30772 23268 39116
rect 23324 37044 23380 39564
rect 23436 38834 23492 39676
rect 23436 38782 23438 38834
rect 23490 38782 23492 38834
rect 23436 38770 23492 38782
rect 23548 37604 23604 40796
rect 23884 40758 23940 40796
rect 24108 42082 24164 42094
rect 24108 42030 24110 42082
rect 24162 42030 24164 42082
rect 23772 40628 23828 40638
rect 24108 40628 24164 42030
rect 24220 41748 24276 41758
rect 24220 41654 24276 41692
rect 24332 40964 24388 45612
rect 25228 45218 25284 46620
rect 25228 45166 25230 45218
rect 25282 45166 25284 45218
rect 25228 45154 25284 45166
rect 25340 45106 25396 45118
rect 25340 45054 25342 45106
rect 25394 45054 25396 45106
rect 24668 44996 24724 45006
rect 24668 44902 24724 44940
rect 24444 44882 24500 44894
rect 24444 44830 24446 44882
rect 24498 44830 24500 44882
rect 24444 44324 24500 44830
rect 24444 44210 24500 44268
rect 24780 44324 24836 44334
rect 24780 44230 24836 44268
rect 25340 44324 25396 45054
rect 24444 44158 24446 44210
rect 24498 44158 24500 44210
rect 24444 44146 24500 44158
rect 25340 42866 25396 44268
rect 25564 44996 25620 45006
rect 25564 44436 25620 44940
rect 25564 44210 25620 44380
rect 25564 44158 25566 44210
rect 25618 44158 25620 44210
rect 25564 44146 25620 44158
rect 25340 42814 25342 42866
rect 25394 42814 25396 42866
rect 25340 42802 25396 42814
rect 25228 42754 25284 42766
rect 25228 42702 25230 42754
rect 25282 42702 25284 42754
rect 25116 42642 25172 42654
rect 25116 42590 25118 42642
rect 25170 42590 25172 42642
rect 25116 42196 25172 42590
rect 25228 42308 25284 42702
rect 25228 42252 25396 42308
rect 25116 42140 25284 42196
rect 24332 40898 24388 40908
rect 24444 42082 24500 42094
rect 24444 42030 24446 42082
rect 24498 42030 24500 42082
rect 23828 40572 24164 40628
rect 24444 40628 24500 42030
rect 24556 42084 24612 42094
rect 24556 41990 24612 42028
rect 24780 41972 24836 41982
rect 25116 41972 25172 41982
rect 24780 41970 25172 41972
rect 24780 41918 24782 41970
rect 24834 41918 25118 41970
rect 25170 41918 25172 41970
rect 24780 41916 25172 41918
rect 24780 41906 24836 41916
rect 25116 41906 25172 41916
rect 25228 41300 25284 42140
rect 25228 41186 25284 41244
rect 25228 41134 25230 41186
rect 25282 41134 25284 41186
rect 25228 41122 25284 41134
rect 25340 41188 25396 42252
rect 25676 41746 25732 56812
rect 26124 56802 26180 56812
rect 26684 56774 26740 56812
rect 26796 56756 26852 56766
rect 26796 56662 26852 56700
rect 26684 54628 26740 54638
rect 26684 54534 26740 54572
rect 26796 54402 26852 54414
rect 26796 54350 26798 54402
rect 26850 54350 26852 54402
rect 26796 53956 26852 54350
rect 26012 53900 26852 53956
rect 26012 53842 26068 53900
rect 26012 53790 26014 53842
rect 26066 53790 26068 53842
rect 26012 53778 26068 53790
rect 26236 50484 26292 50494
rect 26236 50390 26292 50428
rect 26908 50428 26964 57820
rect 27468 57764 27524 58382
rect 27132 57708 27524 57764
rect 27020 57652 27076 57662
rect 27132 57652 27188 57708
rect 27580 57652 27636 58494
rect 28140 58322 28196 61180
rect 28364 60786 28420 60798
rect 28364 60734 28366 60786
rect 28418 60734 28420 60786
rect 28364 60228 28420 60734
rect 28364 60134 28420 60172
rect 28140 58270 28142 58322
rect 28194 58270 28196 58322
rect 28140 58258 28196 58270
rect 28252 57764 28308 57774
rect 28252 57670 28308 57708
rect 27020 57650 27188 57652
rect 27020 57598 27022 57650
rect 27074 57598 27188 57650
rect 27020 57596 27188 57598
rect 27244 57650 27636 57652
rect 27244 57598 27582 57650
rect 27634 57598 27636 57650
rect 27244 57596 27636 57598
rect 27020 55860 27076 57596
rect 27244 57090 27300 57596
rect 27580 57586 27636 57596
rect 27244 57038 27246 57090
rect 27298 57038 27300 57090
rect 27244 57026 27300 57038
rect 27132 56756 27188 56766
rect 27132 56662 27188 56700
rect 27020 55794 27076 55804
rect 27692 56644 27748 56654
rect 27692 55300 27748 56588
rect 28476 56308 28532 62860
rect 28588 62850 28644 62860
rect 28924 62916 28980 62926
rect 28924 62466 28980 62860
rect 29036 62578 29092 63756
rect 29036 62526 29038 62578
rect 29090 62526 29092 62578
rect 29036 62514 29092 62526
rect 28924 62414 28926 62466
rect 28978 62414 28980 62466
rect 28924 62402 28980 62414
rect 29148 62354 29204 64652
rect 29484 64708 29540 64718
rect 29484 64614 29540 64652
rect 30380 64708 30436 64718
rect 30380 64614 30436 64652
rect 30940 64596 30996 64606
rect 32508 64596 32564 64764
rect 30940 64502 30996 64540
rect 32396 64594 32564 64596
rect 32396 64542 32510 64594
rect 32562 64542 32564 64594
rect 32396 64540 32564 64542
rect 29596 64482 29652 64494
rect 29596 64430 29598 64482
rect 29650 64430 29652 64482
rect 29596 63364 29652 64430
rect 29148 62302 29150 62354
rect 29202 62302 29204 62354
rect 29148 62290 29204 62302
rect 29372 63308 29652 63364
rect 29708 64482 29764 64494
rect 29708 64430 29710 64482
rect 29762 64430 29764 64482
rect 29372 62354 29428 63308
rect 29484 63026 29540 63038
rect 29484 62974 29486 63026
rect 29538 62974 29540 63026
rect 29484 62916 29540 62974
rect 29708 62916 29764 64430
rect 30828 64482 30884 64494
rect 30828 64430 30830 64482
rect 30882 64430 30884 64482
rect 30828 63812 30884 64430
rect 31052 64484 31108 64494
rect 31500 64484 31556 64494
rect 32284 64484 32340 64494
rect 31052 64482 31556 64484
rect 31052 64430 31054 64482
rect 31106 64430 31502 64482
rect 31554 64430 31556 64482
rect 31052 64428 31556 64430
rect 30940 63812 30996 63822
rect 30828 63810 30996 63812
rect 30828 63758 30942 63810
rect 30994 63758 30996 63810
rect 30828 63756 30996 63758
rect 30156 63140 30212 63150
rect 30156 63046 30212 63084
rect 30380 63138 30436 63150
rect 30380 63086 30382 63138
rect 30434 63086 30436 63138
rect 29540 62860 29764 62916
rect 29484 62822 29540 62860
rect 29372 62302 29374 62354
rect 29426 62302 29428 62354
rect 29372 62290 29428 62302
rect 29484 62244 29540 62254
rect 30380 62244 30436 63086
rect 30940 63140 30996 63756
rect 30940 63074 30996 63084
rect 31052 63028 31108 64428
rect 31500 64418 31556 64428
rect 32172 64482 32340 64484
rect 32172 64430 32286 64482
rect 32338 64430 32340 64482
rect 32172 64428 32340 64430
rect 31948 64034 32004 64046
rect 31948 63982 31950 64034
rect 32002 63982 32004 64034
rect 31276 63140 31332 63150
rect 31164 63028 31220 63038
rect 31052 63026 31220 63028
rect 31052 62974 31166 63026
rect 31218 62974 31220 63026
rect 31052 62972 31220 62974
rect 30828 62244 30884 62254
rect 31164 62244 31220 62972
rect 31276 63026 31332 63084
rect 31276 62974 31278 63026
rect 31330 62974 31332 63026
rect 31276 62962 31332 62974
rect 31500 62916 31556 62926
rect 31500 62822 31556 62860
rect 31948 62468 32004 63982
rect 32060 63922 32116 63934
rect 32060 63870 32062 63922
rect 32114 63870 32116 63922
rect 32060 63250 32116 63870
rect 32172 63924 32228 64428
rect 32284 64418 32340 64428
rect 32284 64148 32340 64158
rect 32396 64148 32452 64540
rect 32508 64530 32564 64540
rect 32620 64594 32676 64606
rect 32620 64542 32622 64594
rect 32674 64542 32676 64594
rect 32620 64372 32676 64542
rect 32956 64596 33012 64606
rect 32956 64502 33012 64540
rect 33068 64482 33124 64494
rect 33068 64430 33070 64482
rect 33122 64430 33124 64482
rect 33068 64372 33124 64430
rect 33292 64484 33348 64494
rect 33292 64390 33348 64428
rect 32284 64146 32452 64148
rect 32284 64094 32286 64146
rect 32338 64094 32452 64146
rect 32284 64092 32452 64094
rect 32508 64316 32676 64372
rect 32844 64316 33124 64372
rect 32284 64082 32340 64092
rect 32508 63924 32564 64316
rect 32172 63868 32340 63924
rect 32060 63198 32062 63250
rect 32114 63198 32116 63250
rect 32060 63186 32116 63198
rect 32284 63138 32340 63868
rect 32396 63812 32452 63822
rect 32396 63718 32452 63756
rect 32284 63086 32286 63138
rect 32338 63086 32340 63138
rect 32284 63074 32340 63086
rect 32060 62916 32116 62926
rect 32060 62822 32116 62860
rect 32508 62580 32564 63868
rect 32620 64036 32676 64046
rect 32620 63138 32676 63980
rect 32620 63086 32622 63138
rect 32674 63086 32676 63138
rect 32620 63074 32676 63086
rect 32844 62916 32900 64316
rect 33180 63924 33236 63934
rect 33180 63810 33236 63868
rect 33516 63922 33572 64764
rect 33516 63870 33518 63922
rect 33570 63870 33572 63922
rect 33516 63858 33572 63870
rect 33180 63758 33182 63810
rect 33234 63758 33236 63810
rect 33180 63746 33236 63758
rect 32844 62850 32900 62860
rect 32956 62914 33012 62926
rect 32956 62862 32958 62914
rect 33010 62862 33012 62914
rect 32284 62524 32564 62580
rect 32060 62468 32116 62478
rect 31948 62412 32060 62468
rect 32060 62402 32116 62412
rect 31276 62244 31332 62254
rect 30380 62242 31332 62244
rect 30380 62190 30830 62242
rect 30882 62190 31278 62242
rect 31330 62190 31332 62242
rect 30380 62188 31332 62190
rect 29484 62132 29764 62188
rect 29596 61124 29652 61134
rect 29596 60898 29652 61068
rect 29596 60846 29598 60898
rect 29650 60846 29652 60898
rect 29596 60834 29652 60846
rect 28924 60788 28980 60798
rect 28980 60732 29092 60788
rect 28924 60694 28980 60732
rect 28700 60676 28756 60686
rect 28700 60582 28756 60620
rect 29036 60002 29092 60732
rect 29036 59950 29038 60002
rect 29090 59950 29092 60002
rect 29036 59938 29092 59950
rect 29260 60228 29316 60238
rect 29260 59890 29316 60172
rect 29372 60004 29428 60014
rect 29372 59910 29428 59948
rect 29260 59838 29262 59890
rect 29314 59838 29316 59890
rect 29260 59826 29316 59838
rect 29708 58100 29764 62132
rect 30492 62132 30884 62188
rect 31276 62178 31332 62188
rect 30044 60676 30100 60686
rect 30492 60676 30548 62132
rect 32284 61010 32340 62524
rect 32956 62468 33012 62862
rect 32732 61460 32788 61470
rect 32732 61458 32900 61460
rect 32732 61406 32734 61458
rect 32786 61406 32900 61458
rect 32732 61404 32900 61406
rect 32732 61394 32788 61404
rect 32284 60958 32286 61010
rect 32338 60958 32340 61010
rect 31948 60786 32004 60798
rect 31948 60734 31950 60786
rect 32002 60734 32004 60786
rect 30044 60674 30548 60676
rect 30044 60622 30046 60674
rect 30098 60622 30494 60674
rect 30546 60622 30548 60674
rect 30044 60620 30548 60622
rect 30044 60610 30100 60620
rect 29932 60564 29988 60574
rect 29932 60470 29988 60508
rect 30380 60004 30436 60014
rect 30380 59778 30436 59948
rect 30380 59726 30382 59778
rect 30434 59726 30436 59778
rect 29820 58324 29876 58334
rect 29820 58230 29876 58268
rect 29932 58210 29988 58222
rect 29932 58158 29934 58210
rect 29986 58158 29988 58210
rect 29708 58044 29876 58100
rect 29820 57090 29876 58044
rect 29820 57038 29822 57090
rect 29874 57038 29876 57090
rect 29820 57026 29876 57038
rect 29932 56978 29988 58158
rect 30044 58210 30100 58222
rect 30044 58158 30046 58210
rect 30098 58158 30100 58210
rect 30044 57762 30100 58158
rect 30380 58100 30436 59726
rect 30492 58828 30548 60620
rect 31612 60676 31668 60686
rect 31948 60676 32004 60734
rect 31612 60674 32004 60676
rect 31612 60622 31614 60674
rect 31666 60622 32004 60674
rect 31612 60620 32004 60622
rect 31164 60002 31220 60014
rect 31164 59950 31166 60002
rect 31218 59950 31220 60002
rect 30716 59778 30772 59790
rect 30716 59726 30718 59778
rect 30770 59726 30772 59778
rect 30716 59108 30772 59726
rect 31164 59780 31220 59950
rect 30940 59108 30996 59118
rect 31164 59108 31220 59724
rect 30716 59106 31220 59108
rect 30716 59054 30942 59106
rect 30994 59054 31220 59106
rect 30716 59052 31220 59054
rect 31612 60002 31668 60620
rect 32060 60564 32116 60574
rect 32060 60114 32116 60508
rect 32060 60062 32062 60114
rect 32114 60062 32116 60114
rect 32060 60050 32116 60062
rect 31612 59950 31614 60002
rect 31666 59950 31668 60002
rect 31612 59108 31668 59950
rect 32284 59668 32340 60958
rect 32396 61346 32452 61358
rect 32620 61348 32676 61358
rect 32396 61294 32398 61346
rect 32450 61294 32452 61346
rect 32396 60788 32452 61294
rect 32396 60722 32452 60732
rect 32508 61346 32676 61348
rect 32508 61294 32622 61346
rect 32674 61294 32676 61346
rect 32508 61292 32676 61294
rect 32508 60226 32564 61292
rect 32620 61282 32676 61292
rect 32508 60174 32510 60226
rect 32562 60174 32564 60226
rect 32508 60162 32564 60174
rect 32396 60004 32452 60014
rect 32396 59910 32452 59948
rect 32844 60002 32900 61404
rect 32844 59950 32846 60002
rect 32898 59950 32900 60002
rect 32844 59938 32900 59950
rect 32508 59778 32564 59790
rect 32508 59726 32510 59778
rect 32562 59726 32564 59778
rect 32508 59668 32564 59726
rect 32284 59612 32564 59668
rect 30940 59042 30996 59052
rect 30492 58772 30772 58828
rect 30380 58034 30436 58044
rect 30492 58324 30548 58334
rect 30044 57710 30046 57762
rect 30098 57710 30100 57762
rect 30044 57316 30100 57710
rect 30044 57250 30100 57260
rect 30156 57652 30212 57662
rect 29932 56926 29934 56978
rect 29986 56926 29988 56978
rect 29932 56914 29988 56926
rect 28364 56306 28532 56308
rect 28364 56254 28478 56306
rect 28530 56254 28532 56306
rect 28364 56252 28532 56254
rect 28364 55300 28420 56252
rect 28476 56242 28532 56252
rect 30156 56866 30212 57596
rect 30268 57652 30324 57662
rect 30492 57652 30548 58268
rect 30268 57650 30548 57652
rect 30268 57598 30270 57650
rect 30322 57598 30548 57650
rect 30268 57596 30548 57598
rect 30604 58210 30660 58222
rect 30604 58158 30606 58210
rect 30658 58158 30660 58210
rect 30268 57586 30324 57596
rect 30156 56814 30158 56866
rect 30210 56814 30212 56866
rect 30156 55524 30212 56814
rect 30156 55468 30324 55524
rect 27692 55244 28084 55300
rect 27020 55076 27076 55086
rect 27692 55076 27748 55086
rect 27020 54626 27076 55020
rect 27020 54574 27022 54626
rect 27074 54574 27076 54626
rect 27020 54562 27076 54574
rect 27580 55074 27748 55076
rect 27580 55022 27694 55074
rect 27746 55022 27748 55074
rect 27580 55020 27748 55022
rect 27244 54514 27300 54526
rect 27244 54462 27246 54514
rect 27298 54462 27300 54514
rect 27244 54292 27300 54462
rect 27580 54516 27636 55020
rect 27692 55010 27748 55020
rect 27804 55074 27860 55086
rect 27804 55022 27806 55074
rect 27858 55022 27860 55074
rect 27580 54422 27636 54460
rect 27804 54292 27860 55022
rect 27916 55076 27972 55086
rect 27916 54982 27972 55020
rect 27244 54236 27860 54292
rect 28028 50428 28084 55244
rect 28252 55298 28420 55300
rect 28252 55246 28366 55298
rect 28418 55246 28420 55298
rect 28252 55244 28420 55246
rect 28140 54514 28196 54526
rect 28140 54462 28142 54514
rect 28194 54462 28196 54514
rect 28140 53844 28196 54462
rect 28140 53750 28196 53788
rect 28252 50428 28308 55244
rect 28364 55234 28420 55244
rect 29260 55298 29316 55310
rect 30156 55300 30212 55310
rect 29260 55246 29262 55298
rect 29314 55246 29316 55298
rect 28476 54404 28532 54414
rect 28476 54310 28532 54348
rect 28924 54402 28980 54414
rect 28924 54350 28926 54402
rect 28978 54350 28980 54402
rect 28924 53844 28980 54350
rect 29148 54404 29204 54414
rect 29260 54404 29316 55246
rect 29484 55298 30212 55300
rect 29484 55246 30158 55298
rect 30210 55246 30212 55298
rect 29484 55244 30212 55246
rect 29372 55186 29428 55198
rect 29372 55134 29374 55186
rect 29426 55134 29428 55186
rect 29372 55076 29428 55134
rect 29372 54516 29428 55020
rect 29484 54738 29540 55244
rect 30156 55234 30212 55244
rect 30156 55076 30212 55086
rect 30268 55076 30324 55468
rect 30380 55188 30436 57596
rect 30604 57316 30660 58158
rect 30604 57250 30660 57260
rect 30716 56644 30772 58772
rect 30828 58210 30884 58222
rect 30828 58158 30830 58210
rect 30882 58158 30884 58210
rect 30828 56866 30884 58158
rect 30940 57652 30996 57662
rect 30940 57558 30996 57596
rect 30828 56814 30830 56866
rect 30882 56814 30884 56866
rect 30828 56802 30884 56814
rect 30716 56588 30884 56644
rect 30716 55188 30772 55198
rect 30380 55132 30716 55188
rect 30716 55094 30772 55132
rect 30156 55074 30324 55076
rect 30156 55022 30158 55074
rect 30210 55022 30324 55074
rect 30156 55020 30324 55022
rect 30156 55010 30212 55020
rect 29484 54686 29486 54738
rect 29538 54686 29540 54738
rect 29484 54674 29540 54686
rect 29372 54460 29876 54516
rect 29260 54348 29764 54404
rect 29148 54068 29204 54348
rect 29148 54012 29428 54068
rect 29372 53956 29428 54012
rect 29372 53862 29428 53900
rect 29708 53954 29764 54348
rect 29708 53902 29710 53954
rect 29762 53902 29764 53954
rect 29708 53890 29764 53902
rect 29148 53844 29204 53854
rect 28980 53842 29204 53844
rect 28980 53790 29150 53842
rect 29202 53790 29204 53842
rect 28980 53788 29204 53790
rect 28924 53750 28980 53788
rect 29148 53778 29204 53788
rect 28924 53508 28980 53518
rect 28364 51378 28420 51390
rect 28364 51326 28366 51378
rect 28418 51326 28420 51378
rect 28364 50762 28420 51326
rect 28476 51380 28532 51390
rect 28532 51324 28756 51380
rect 28476 51286 28532 51324
rect 28364 50710 28366 50762
rect 28418 50710 28420 50762
rect 28364 50698 28420 50710
rect 26908 50372 27188 50428
rect 25788 49140 25844 49150
rect 25788 49046 25844 49084
rect 26124 48244 26180 48254
rect 25900 47570 25956 47582
rect 25900 47518 25902 47570
rect 25954 47518 25956 47570
rect 25900 46676 25956 47518
rect 26124 47346 26180 48188
rect 26908 47796 26964 47806
rect 26908 47348 26964 47740
rect 26124 47294 26126 47346
rect 26178 47294 26180 47346
rect 26124 47282 26180 47294
rect 26796 47292 26964 47348
rect 26012 46676 26068 46686
rect 25900 46674 26068 46676
rect 25900 46622 26014 46674
rect 26066 46622 26068 46674
rect 25900 46620 26068 46622
rect 26012 46564 26068 46620
rect 26012 46498 26068 46508
rect 26236 46564 26292 46574
rect 26236 45780 26292 46508
rect 26796 46562 26852 47292
rect 26796 46510 26798 46562
rect 26850 46510 26852 46562
rect 26796 46498 26852 46510
rect 26236 45714 26292 45724
rect 27020 45892 27076 45902
rect 25788 45106 25844 45118
rect 25788 45054 25790 45106
rect 25842 45054 25844 45106
rect 25788 44322 25844 45054
rect 25788 44270 25790 44322
rect 25842 44270 25844 44322
rect 25788 43708 25844 44270
rect 25788 43652 26404 43708
rect 26012 42756 26068 42766
rect 26012 42662 26068 42700
rect 26236 42754 26292 42766
rect 26236 42702 26238 42754
rect 26290 42702 26292 42754
rect 25900 41972 25956 41982
rect 26236 41972 26292 42702
rect 25900 41970 26292 41972
rect 25900 41918 25902 41970
rect 25954 41918 26292 41970
rect 25900 41916 26292 41918
rect 25676 41694 25678 41746
rect 25730 41694 25732 41746
rect 25676 41682 25732 41694
rect 25788 41858 25844 41870
rect 25788 41806 25790 41858
rect 25842 41806 25844 41858
rect 25564 41298 25620 41310
rect 25564 41246 25566 41298
rect 25618 41246 25620 41298
rect 25452 41188 25508 41198
rect 25340 41186 25508 41188
rect 25340 41134 25454 41186
rect 25506 41134 25508 41186
rect 25340 41132 25508 41134
rect 25452 40964 25508 41132
rect 25564 41188 25620 41246
rect 25564 41122 25620 41132
rect 25564 40964 25620 40974
rect 25452 40908 25564 40964
rect 25564 40898 25620 40908
rect 23660 39620 23716 39630
rect 23660 38834 23716 39564
rect 23660 38782 23662 38834
rect 23714 38782 23716 38834
rect 23660 38770 23716 38782
rect 23772 39618 23828 40572
rect 24444 40516 24500 40572
rect 24108 40460 24500 40516
rect 23884 40404 23940 40414
rect 23884 40310 23940 40348
rect 23772 39566 23774 39618
rect 23826 39566 23828 39618
rect 23548 37538 23604 37548
rect 23660 37378 23716 37390
rect 23660 37326 23662 37378
rect 23714 37326 23716 37378
rect 23660 37044 23716 37326
rect 23324 36988 23716 37044
rect 23660 36370 23716 36988
rect 23660 36318 23662 36370
rect 23714 36318 23716 36370
rect 23324 35924 23380 35934
rect 23324 35830 23380 35868
rect 23660 35700 23716 36318
rect 23660 35634 23716 35644
rect 23324 35364 23380 35374
rect 23324 31218 23380 35308
rect 23772 34580 23828 39566
rect 24108 39394 24164 40460
rect 25004 39732 25060 39742
rect 24668 39620 24724 39630
rect 24724 39564 24836 39620
rect 24668 39554 24724 39564
rect 24108 39342 24110 39394
rect 24162 39342 24164 39394
rect 24108 39330 24164 39342
rect 24220 39396 24276 39406
rect 23884 38836 23940 38846
rect 23884 38742 23940 38780
rect 24108 38834 24164 38846
rect 24108 38782 24110 38834
rect 24162 38782 24164 38834
rect 24108 38668 24164 38782
rect 23884 38612 24164 38668
rect 23884 37492 23940 38612
rect 24220 38610 24276 39340
rect 24220 38558 24222 38610
rect 24274 38558 24276 38610
rect 24220 38500 24276 38558
rect 23996 38444 24276 38500
rect 24332 38948 24388 38958
rect 23996 37940 24052 38444
rect 23996 37846 24052 37884
rect 24220 38052 24276 38062
rect 24332 38052 24388 38892
rect 24556 38724 24612 38734
rect 24556 38274 24612 38668
rect 24556 38222 24558 38274
rect 24610 38222 24612 38274
rect 24556 38210 24612 38222
rect 24220 38050 24388 38052
rect 24220 37998 24222 38050
rect 24274 37998 24388 38050
rect 24220 37996 24388 37998
rect 24668 38164 24724 38174
rect 23996 37604 24052 37614
rect 24052 37548 24164 37604
rect 23996 37538 24052 37548
rect 23884 37426 23940 37436
rect 23996 36932 24052 36942
rect 23548 34524 23828 34580
rect 23884 36876 23996 36932
rect 23548 34018 23604 34524
rect 23884 34132 23940 36876
rect 23996 36866 24052 36876
rect 24108 36594 24164 37548
rect 24220 37492 24276 37996
rect 24556 37492 24612 37502
rect 24220 37490 24612 37492
rect 24220 37438 24558 37490
rect 24610 37438 24612 37490
rect 24220 37436 24612 37438
rect 24556 37426 24612 37436
rect 24668 37268 24724 38108
rect 24556 37266 24724 37268
rect 24556 37214 24670 37266
rect 24722 37214 24724 37266
rect 24556 37212 24724 37214
rect 24556 36706 24612 37212
rect 24668 37202 24724 37212
rect 24556 36654 24558 36706
rect 24610 36654 24612 36706
rect 24556 36642 24612 36654
rect 24108 36542 24110 36594
rect 24162 36542 24164 36594
rect 24108 36530 24164 36542
rect 23996 36482 24052 36494
rect 23996 36430 23998 36482
rect 24050 36430 24052 36482
rect 23996 35698 24052 36430
rect 24332 36484 24388 36494
rect 24668 36484 24724 36494
rect 24780 36484 24836 39564
rect 25004 39506 25060 39676
rect 25004 39454 25006 39506
rect 25058 39454 25060 39506
rect 25004 39442 25060 39454
rect 25564 39618 25620 39630
rect 25788 39620 25844 41806
rect 25900 41186 25956 41916
rect 25900 41134 25902 41186
rect 25954 41134 25956 41186
rect 25900 41122 25956 41134
rect 26012 41188 26068 41198
rect 26012 39842 26068 41132
rect 26348 40180 26404 43652
rect 26908 41970 26964 41982
rect 26908 41918 26910 41970
rect 26962 41918 26964 41970
rect 26572 41748 26628 41758
rect 26572 41186 26628 41692
rect 26572 41134 26574 41186
rect 26626 41134 26628 41186
rect 26572 41122 26628 41134
rect 26908 41188 26964 41918
rect 27020 41412 27076 45836
rect 27132 43988 27188 50372
rect 27804 50372 28084 50428
rect 28140 50372 28308 50428
rect 28364 50596 28420 50606
rect 27356 49476 27412 49486
rect 27356 48466 27412 49420
rect 27356 48414 27358 48466
rect 27410 48414 27412 48466
rect 27356 48402 27412 48414
rect 27244 48242 27300 48254
rect 27244 48190 27246 48242
rect 27298 48190 27300 48242
rect 27244 47796 27300 48190
rect 27244 47730 27300 47740
rect 27468 48244 27524 48254
rect 27356 47458 27412 47470
rect 27356 47406 27358 47458
rect 27410 47406 27412 47458
rect 27244 47348 27300 47358
rect 27244 46898 27300 47292
rect 27244 46846 27246 46898
rect 27298 46846 27300 46898
rect 27244 46834 27300 46846
rect 27356 46564 27412 47406
rect 27468 47012 27524 48188
rect 27468 46956 27636 47012
rect 27356 46498 27412 46508
rect 27468 46674 27524 46686
rect 27468 46622 27470 46674
rect 27522 46622 27524 46674
rect 27468 46004 27524 46622
rect 27580 46114 27636 46956
rect 27580 46062 27582 46114
rect 27634 46062 27636 46114
rect 27580 46050 27636 46062
rect 27468 45938 27524 45948
rect 27244 45892 27300 45902
rect 27244 45798 27300 45836
rect 27132 43932 27412 43988
rect 27132 42756 27188 42766
rect 27132 42662 27188 42700
rect 27244 42084 27300 42094
rect 27244 41990 27300 42028
rect 27132 41412 27188 41422
rect 27020 41410 27188 41412
rect 27020 41358 27134 41410
rect 27186 41358 27188 41410
rect 27020 41356 27188 41358
rect 27132 41346 27188 41356
rect 27356 41410 27412 43932
rect 27356 41358 27358 41410
rect 27410 41358 27412 41410
rect 27356 41346 27412 41358
rect 27468 42754 27524 42766
rect 27468 42702 27470 42754
rect 27522 42702 27524 42754
rect 27468 41300 27524 42702
rect 27692 42754 27748 42766
rect 27692 42702 27694 42754
rect 27746 42702 27748 42754
rect 27692 42644 27748 42702
rect 27468 41234 27524 41244
rect 27580 42588 27692 42644
rect 26908 41122 26964 41132
rect 26460 41076 26516 41086
rect 26460 40982 26516 41020
rect 26684 41074 26740 41086
rect 26684 41022 26686 41074
rect 26738 41022 26740 41074
rect 26348 40114 26404 40124
rect 26012 39790 26014 39842
rect 26066 39790 26068 39842
rect 26012 39778 26068 39790
rect 26124 39732 26180 39742
rect 26124 39638 26180 39676
rect 25564 39566 25566 39618
rect 25618 39566 25620 39618
rect 25564 39508 25620 39566
rect 25564 38722 25620 39452
rect 25564 38670 25566 38722
rect 25618 38670 25620 38722
rect 25340 37492 25396 37502
rect 25340 37398 25396 37436
rect 25228 37156 25284 37166
rect 25228 37062 25284 37100
rect 24220 36036 24276 36046
rect 24220 35922 24276 35980
rect 24220 35870 24222 35922
rect 24274 35870 24276 35922
rect 24220 35858 24276 35870
rect 23996 35646 23998 35698
rect 24050 35646 24052 35698
rect 23996 35028 24052 35646
rect 24220 35028 24276 35038
rect 23996 35026 24276 35028
rect 23996 34974 24222 35026
rect 24274 34974 24276 35026
rect 23996 34972 24276 34974
rect 24220 34962 24276 34972
rect 23884 34130 24276 34132
rect 23884 34078 23886 34130
rect 23938 34078 24276 34130
rect 23884 34076 24276 34078
rect 23884 34066 23940 34076
rect 23548 33966 23550 34018
rect 23602 33966 23604 34018
rect 23548 33572 23604 33966
rect 23548 33506 23604 33516
rect 24220 33458 24276 34076
rect 24220 33406 24222 33458
rect 24274 33406 24276 33458
rect 24220 33394 24276 33406
rect 24332 33236 24388 36428
rect 24108 33180 24388 33236
rect 24444 36482 24836 36484
rect 24444 36430 24670 36482
rect 24722 36430 24836 36482
rect 24444 36428 24836 36430
rect 25228 36932 25284 36942
rect 23324 31166 23326 31218
rect 23378 31166 23380 31218
rect 23324 31154 23380 31166
rect 23884 33124 23940 33134
rect 23884 31778 23940 33068
rect 24108 32786 24164 33180
rect 24444 32788 24500 36428
rect 24668 36418 24724 36428
rect 25228 36036 25284 36876
rect 25228 35922 25284 35980
rect 25228 35870 25230 35922
rect 25282 35870 25284 35922
rect 25228 35858 25284 35870
rect 25452 35588 25508 35598
rect 25564 35588 25620 38670
rect 25676 39564 25844 39620
rect 26236 39620 26292 39630
rect 25676 38834 25732 39564
rect 26236 39526 26292 39564
rect 26572 39618 26628 39630
rect 26572 39566 26574 39618
rect 26626 39566 26628 39618
rect 26572 39508 26628 39566
rect 26572 39442 26628 39452
rect 26684 39060 26740 41022
rect 27356 41076 27412 41086
rect 26684 38994 26740 39004
rect 27132 40402 27188 40414
rect 27132 40350 27134 40402
rect 27186 40350 27188 40402
rect 27132 38948 27188 40350
rect 25676 38782 25678 38834
rect 25730 38782 25732 38834
rect 25676 38724 25732 38782
rect 26348 38836 26404 38846
rect 26348 38742 26404 38780
rect 27020 38836 27076 38846
rect 27132 38836 27188 38892
rect 27020 38834 27188 38836
rect 27020 38782 27022 38834
rect 27074 38782 27188 38834
rect 27020 38780 27188 38782
rect 27244 40404 27300 40414
rect 27244 38834 27300 40348
rect 27244 38782 27246 38834
rect 27298 38782 27300 38834
rect 27020 38770 27076 38780
rect 25676 38658 25732 38668
rect 26012 38724 26068 38734
rect 26012 38274 26068 38668
rect 26796 38610 26852 38622
rect 26796 38558 26798 38610
rect 26850 38558 26852 38610
rect 26012 38222 26014 38274
rect 26066 38222 26068 38274
rect 26012 38210 26068 38222
rect 26124 38500 26180 38510
rect 26124 38050 26180 38444
rect 26796 38388 26852 38558
rect 26796 38322 26852 38332
rect 26908 38500 26964 38510
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 26124 37986 26180 37998
rect 26572 38052 26628 38062
rect 26012 37828 26068 37838
rect 26012 37378 26068 37772
rect 26012 37326 26014 37378
rect 26066 37326 26068 37378
rect 26012 36932 26068 37326
rect 26124 37380 26180 37390
rect 26124 37286 26180 37324
rect 26572 37266 26628 37996
rect 26572 37214 26574 37266
rect 26626 37214 26628 37266
rect 26572 37202 26628 37214
rect 26796 37378 26852 37390
rect 26796 37326 26798 37378
rect 26850 37326 26852 37378
rect 26796 37268 26852 37326
rect 26796 37202 26852 37212
rect 26012 36866 26068 36876
rect 26908 36708 26964 38444
rect 27020 38164 27076 38174
rect 27020 38070 27076 38108
rect 27132 38050 27188 38062
rect 27132 37998 27134 38050
rect 27186 37998 27188 38050
rect 27132 37380 27188 37998
rect 27132 37266 27188 37324
rect 27132 37214 27134 37266
rect 27186 37214 27188 37266
rect 27132 37202 27188 37214
rect 27244 37042 27300 38782
rect 27356 38274 27412 41020
rect 27468 40964 27524 40974
rect 27468 40870 27524 40908
rect 27580 40628 27636 42588
rect 27692 42578 27748 42588
rect 27804 42420 27860 50372
rect 28140 48356 28196 50372
rect 28364 49922 28420 50540
rect 28700 50428 28756 51324
rect 28476 50372 28756 50428
rect 28924 50428 28980 53452
rect 29148 51380 29204 51390
rect 29204 51324 29540 51380
rect 29148 51286 29204 51324
rect 29036 51266 29092 51278
rect 29036 51214 29038 51266
rect 29090 51214 29092 51266
rect 29036 50820 29092 51214
rect 29036 50596 29092 50764
rect 29372 50708 29428 50718
rect 29260 50596 29316 50606
rect 29036 50540 29260 50596
rect 29260 50502 29316 50540
rect 28924 50372 29204 50428
rect 28476 50034 28532 50372
rect 28476 49982 28478 50034
rect 28530 49982 28532 50034
rect 28476 49970 28532 49982
rect 28700 50036 28756 50046
rect 28700 49942 28756 49980
rect 28364 49870 28366 49922
rect 28418 49870 28420 49922
rect 28364 49858 28420 49870
rect 29036 49922 29092 49934
rect 29036 49870 29038 49922
rect 29090 49870 29092 49922
rect 29036 49812 29092 49870
rect 29036 49746 29092 49756
rect 28140 48300 28532 48356
rect 27916 48242 27972 48254
rect 27916 48190 27918 48242
rect 27970 48190 27972 48242
rect 27916 47684 27972 48190
rect 28364 47684 28420 47694
rect 27916 47682 28420 47684
rect 27916 47630 28366 47682
rect 28418 47630 28420 47682
rect 27916 47628 28420 47630
rect 28364 47618 28420 47628
rect 27916 47460 27972 47470
rect 27916 47366 27972 47404
rect 28252 47348 28308 47358
rect 28252 47254 28308 47292
rect 28364 47234 28420 47246
rect 28364 47182 28366 47234
rect 28418 47182 28420 47234
rect 28364 47124 28420 47182
rect 28364 47058 28420 47068
rect 28476 46900 28532 48300
rect 29148 47684 29204 50372
rect 29372 50034 29428 50652
rect 29484 50594 29540 51324
rect 29820 51266 29876 54460
rect 30604 54402 30660 54414
rect 30604 54350 30606 54402
rect 30658 54350 30660 54402
rect 30380 53844 30436 53854
rect 30380 53618 30436 53788
rect 30380 53566 30382 53618
rect 30434 53566 30436 53618
rect 30380 53554 30436 53566
rect 30044 53508 30100 53518
rect 30044 53414 30100 53452
rect 30604 53508 30660 54350
rect 30604 53442 30660 53452
rect 30716 53732 30772 53742
rect 30716 52836 30772 53676
rect 30828 52948 30884 56588
rect 31052 55300 31108 59052
rect 31612 59042 31668 59052
rect 32284 59108 32340 59118
rect 32284 59014 32340 59052
rect 32284 57762 32340 57774
rect 32284 57710 32286 57762
rect 32338 57710 32340 57762
rect 31612 57540 31668 57550
rect 32060 57540 32116 57550
rect 31612 57538 32116 57540
rect 31612 57486 31614 57538
rect 31666 57486 32062 57538
rect 32114 57486 32116 57538
rect 31612 57484 32116 57486
rect 31612 57474 31668 57484
rect 32060 57474 32116 57484
rect 32284 57540 32340 57710
rect 32284 57474 32340 57484
rect 32844 57540 32900 57550
rect 32396 57426 32452 57438
rect 32396 57374 32398 57426
rect 32450 57374 32452 57426
rect 31612 57316 31668 57326
rect 31612 56978 31668 57260
rect 31612 56926 31614 56978
rect 31666 56926 31668 56978
rect 31612 56914 31668 56926
rect 32396 56980 32452 57374
rect 32396 56914 32452 56924
rect 31836 56196 31892 56206
rect 31724 56194 31892 56196
rect 31724 56142 31838 56194
rect 31890 56142 31892 56194
rect 31724 56140 31892 56142
rect 31388 55970 31444 55982
rect 31388 55918 31390 55970
rect 31442 55918 31444 55970
rect 31388 55524 31444 55918
rect 30940 55244 31108 55300
rect 31164 55468 31444 55524
rect 30940 54180 30996 55244
rect 31052 55076 31108 55086
rect 31164 55076 31220 55468
rect 31612 55300 31668 55310
rect 31052 55074 31220 55076
rect 31052 55022 31054 55074
rect 31106 55022 31220 55074
rect 31052 55020 31220 55022
rect 31388 55186 31444 55198
rect 31388 55134 31390 55186
rect 31442 55134 31444 55186
rect 31052 54514 31108 55020
rect 31052 54462 31054 54514
rect 31106 54462 31108 54514
rect 31052 54404 31108 54462
rect 31052 54338 31108 54348
rect 30940 54124 31220 54180
rect 30828 52882 30884 52892
rect 30716 52050 30772 52780
rect 30716 51998 30718 52050
rect 30770 51998 30772 52050
rect 30716 51986 30772 51998
rect 30940 52164 30996 52174
rect 30940 51604 30996 52108
rect 30716 51548 30996 51604
rect 30156 51380 30212 51390
rect 29820 51214 29822 51266
rect 29874 51214 29876 51266
rect 29820 51202 29876 51214
rect 30044 51378 30212 51380
rect 30044 51326 30158 51378
rect 30210 51326 30212 51378
rect 30044 51324 30212 51326
rect 29484 50542 29486 50594
rect 29538 50542 29540 50594
rect 29484 50530 29540 50542
rect 29596 50596 29652 50606
rect 29372 49982 29374 50034
rect 29426 49982 29428 50034
rect 29372 49970 29428 49982
rect 29484 50036 29540 50046
rect 29596 50036 29652 50540
rect 30044 50428 30100 51324
rect 30156 51314 30212 51324
rect 30156 50596 30212 50634
rect 30380 50596 30436 50606
rect 30212 50594 30436 50596
rect 30212 50542 30382 50594
rect 30434 50542 30436 50594
rect 30212 50540 30436 50542
rect 30156 50530 30212 50540
rect 30380 50530 30436 50540
rect 30604 50484 30660 50522
rect 29932 50372 29988 50382
rect 30044 50372 30212 50428
rect 30604 50418 30660 50428
rect 29484 50034 29652 50036
rect 29484 49982 29486 50034
rect 29538 49982 29652 50034
rect 29484 49980 29652 49982
rect 29820 50036 29876 50046
rect 29484 49970 29540 49980
rect 29820 49922 29876 49980
rect 29820 49870 29822 49922
rect 29874 49870 29876 49922
rect 29820 49858 29876 49870
rect 29932 49922 29988 50316
rect 30156 50034 30212 50372
rect 30156 49982 30158 50034
rect 30210 49982 30212 50034
rect 30156 49970 30212 49982
rect 29932 49870 29934 49922
rect 29986 49870 29988 49922
rect 29036 47628 29204 47684
rect 29260 49810 29316 49822
rect 29260 49758 29262 49810
rect 29314 49758 29316 49810
rect 29260 49700 29316 49758
rect 29932 49700 29988 49870
rect 29260 49644 29988 49700
rect 30492 49812 30548 49822
rect 30492 49698 30548 49756
rect 30492 49646 30494 49698
rect 30546 49646 30548 49698
rect 29036 47460 29092 47628
rect 29036 47404 29204 47460
rect 28252 46844 28532 46900
rect 28588 47124 28644 47134
rect 27916 45890 27972 45902
rect 27916 45838 27918 45890
rect 27970 45838 27972 45890
rect 27916 45108 27972 45838
rect 27916 45042 27972 45052
rect 28028 42420 28084 42430
rect 27804 42364 28028 42420
rect 28028 42354 28084 42364
rect 28028 42194 28084 42206
rect 28028 42142 28030 42194
rect 28082 42142 28084 42194
rect 27916 42084 27972 42094
rect 27916 41970 27972 42028
rect 27916 41918 27918 41970
rect 27970 41918 27972 41970
rect 27916 41906 27972 41918
rect 28028 41972 28084 42142
rect 28028 41906 28084 41916
rect 28140 41970 28196 41982
rect 28140 41918 28142 41970
rect 28194 41918 28196 41970
rect 28140 41860 28196 41918
rect 27692 41746 27748 41758
rect 27692 41694 27694 41746
rect 27746 41694 27748 41746
rect 27692 41188 27748 41694
rect 28140 41300 28196 41804
rect 27692 41122 27748 41132
rect 27804 41244 28196 41300
rect 27692 40964 27748 40974
rect 27804 40964 27860 41244
rect 27692 40962 27860 40964
rect 27692 40910 27694 40962
rect 27746 40910 27860 40962
rect 27692 40908 27860 40910
rect 27692 40898 27748 40908
rect 27580 40572 27748 40628
rect 27580 40404 27636 40414
rect 27580 40290 27636 40348
rect 27580 40238 27582 40290
rect 27634 40238 27636 40290
rect 27580 40226 27636 40238
rect 27692 39732 27748 40572
rect 27804 40516 27860 40908
rect 27804 40402 27860 40460
rect 27804 40350 27806 40402
rect 27858 40350 27860 40402
rect 27804 40338 27860 40350
rect 27916 41076 27972 41086
rect 27916 40068 27972 41020
rect 28028 40964 28084 40974
rect 28028 40290 28084 40908
rect 28028 40238 28030 40290
rect 28082 40238 28084 40290
rect 28028 40226 28084 40238
rect 27916 40012 28196 40068
rect 27916 39732 27972 39742
rect 27692 39730 27972 39732
rect 27692 39678 27918 39730
rect 27970 39678 27972 39730
rect 27692 39676 27972 39678
rect 27916 39666 27972 39676
rect 27468 39396 27524 39406
rect 27524 39340 27972 39396
rect 27468 39302 27524 39340
rect 27692 39060 27748 39070
rect 27692 38966 27748 39004
rect 27916 39058 27972 39340
rect 27916 39006 27918 39058
rect 27970 39006 27972 39058
rect 27916 38994 27972 39006
rect 28028 38836 28084 38846
rect 28028 38742 28084 38780
rect 27356 38222 27358 38274
rect 27410 38222 27412 38274
rect 27356 38210 27412 38222
rect 28140 38162 28196 40012
rect 28252 38276 28308 46844
rect 28588 46786 28644 47068
rect 28588 46734 28590 46786
rect 28642 46734 28644 46786
rect 28588 46564 28644 46734
rect 28700 46788 28756 46798
rect 28700 46694 28756 46732
rect 28924 46676 28980 46686
rect 28924 46674 29092 46676
rect 28924 46622 28926 46674
rect 28978 46622 29092 46674
rect 28924 46620 29092 46622
rect 28924 46610 28980 46620
rect 28588 46508 28756 46564
rect 28588 45668 28644 45678
rect 28476 45666 28644 45668
rect 28476 45614 28590 45666
rect 28642 45614 28644 45666
rect 28476 45612 28644 45614
rect 28476 45108 28532 45612
rect 28588 45602 28644 45612
rect 28700 45330 28756 46508
rect 29036 45890 29092 46620
rect 29036 45838 29038 45890
rect 29090 45838 29092 45890
rect 29036 45826 29092 45838
rect 29148 45892 29204 47404
rect 29260 46114 29316 49644
rect 30492 48804 30548 49646
rect 30492 48738 30548 48748
rect 29708 47570 29764 47582
rect 29708 47518 29710 47570
rect 29762 47518 29764 47570
rect 29372 47346 29428 47358
rect 29372 47294 29374 47346
rect 29426 47294 29428 47346
rect 29372 47124 29428 47294
rect 29708 47348 29764 47518
rect 29708 47292 30100 47348
rect 29372 46562 29428 47068
rect 29596 47234 29652 47246
rect 29596 47182 29598 47234
rect 29650 47182 29652 47234
rect 29596 46900 29652 47182
rect 29596 46844 29876 46900
rect 29372 46510 29374 46562
rect 29426 46510 29428 46562
rect 29372 46498 29428 46510
rect 29820 46788 29876 46844
rect 29260 46062 29262 46114
rect 29314 46062 29316 46114
rect 29260 46050 29316 46062
rect 29820 46004 29876 46732
rect 29820 45938 29876 45948
rect 30044 46002 30100 47292
rect 30716 46900 30772 51548
rect 30940 50708 30996 50718
rect 30940 50594 30996 50652
rect 30940 50542 30942 50594
rect 30994 50542 30996 50594
rect 30940 50530 30996 50542
rect 30828 50484 30884 50522
rect 30828 50418 30884 50428
rect 31052 49700 31108 49710
rect 31052 49606 31108 49644
rect 30380 46844 30772 46900
rect 30940 49028 30996 49038
rect 30044 45950 30046 46002
rect 30098 45950 30100 46002
rect 30044 45938 30100 45950
rect 30156 46228 30212 46238
rect 29148 45836 29540 45892
rect 28700 45278 28702 45330
rect 28754 45278 28756 45330
rect 28700 45266 28756 45278
rect 28476 45014 28532 45052
rect 29148 45108 29204 45118
rect 29148 44996 29204 45052
rect 29148 44994 29428 44996
rect 29148 44942 29150 44994
rect 29202 44942 29428 44994
rect 29148 44940 29428 44942
rect 29148 44930 29204 44940
rect 28364 42868 28420 42878
rect 28364 42756 28420 42812
rect 29148 42756 29204 42766
rect 28364 42754 28644 42756
rect 28364 42702 28366 42754
rect 28418 42702 28644 42754
rect 28364 42700 28644 42702
rect 28364 42690 28420 42700
rect 28476 42532 28532 42542
rect 28476 42438 28532 42476
rect 28364 42420 28420 42430
rect 28364 38612 28420 42364
rect 28588 42308 28644 42700
rect 29148 42662 29204 42700
rect 28700 42532 28756 42542
rect 29260 42532 29316 42542
rect 28700 42530 29316 42532
rect 28700 42478 28702 42530
rect 28754 42478 29262 42530
rect 29314 42478 29316 42530
rect 28700 42476 29316 42478
rect 28700 42466 28756 42476
rect 29260 42466 29316 42476
rect 28476 42252 28644 42308
rect 28924 42308 28980 42318
rect 29372 42308 29428 44940
rect 29484 42530 29540 45836
rect 30156 45890 30212 46172
rect 30156 45838 30158 45890
rect 30210 45838 30212 45890
rect 30156 45826 30212 45838
rect 29820 43652 29876 43662
rect 29820 43558 29876 43596
rect 29708 43538 29764 43550
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29708 42644 29764 43486
rect 29932 43538 29988 43550
rect 29932 43486 29934 43538
rect 29986 43486 29988 43538
rect 29932 42868 29988 43486
rect 29932 42802 29988 42812
rect 30268 43538 30324 43550
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 29708 42578 29764 42588
rect 30044 42754 30100 42766
rect 30044 42702 30046 42754
rect 30098 42702 30100 42754
rect 29484 42478 29486 42530
rect 29538 42478 29540 42530
rect 29484 42466 29540 42478
rect 29372 42252 29652 42308
rect 28476 42194 28532 42252
rect 28812 42196 28868 42206
rect 28476 42142 28478 42194
rect 28530 42142 28532 42194
rect 28476 42084 28532 42142
rect 28476 42018 28532 42028
rect 28588 42140 28812 42196
rect 28588 41970 28644 42140
rect 28812 42130 28868 42140
rect 28588 41918 28590 41970
rect 28642 41918 28644 41970
rect 28588 41906 28644 41918
rect 28700 41972 28756 41982
rect 28924 41972 28980 42252
rect 28700 41970 28980 41972
rect 28700 41918 28702 41970
rect 28754 41918 28980 41970
rect 28700 41916 28980 41918
rect 29036 41970 29092 41982
rect 29036 41918 29038 41970
rect 29090 41918 29092 41970
rect 28700 40964 28756 41916
rect 29036 41186 29092 41918
rect 29484 41972 29540 41982
rect 29484 41878 29540 41916
rect 29036 41134 29038 41186
rect 29090 41134 29092 41186
rect 29036 41122 29092 41134
rect 29372 41074 29428 41086
rect 29372 41022 29374 41074
rect 29426 41022 29428 41074
rect 29260 40964 29316 40974
rect 28700 40962 29316 40964
rect 28700 40910 29262 40962
rect 29314 40910 29316 40962
rect 28700 40908 29316 40910
rect 28924 40628 28980 40638
rect 28924 40402 28980 40572
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 40338 28980 40350
rect 28588 40180 28644 40190
rect 28588 38668 28644 40124
rect 28588 38612 28756 38668
rect 28364 38546 28420 38556
rect 28252 38220 28532 38276
rect 28140 38110 28142 38162
rect 28194 38110 28196 38162
rect 28140 38098 28196 38110
rect 27468 38052 27524 38062
rect 27468 37958 27524 37996
rect 28252 38052 28308 38062
rect 27580 37940 27636 37950
rect 27580 37492 27636 37884
rect 28140 37940 28196 37950
rect 28140 37846 28196 37884
rect 27580 37266 27636 37436
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 37202 27636 37214
rect 27244 36990 27246 37042
rect 27298 36990 27300 37042
rect 27244 36978 27300 36990
rect 27356 36708 27412 36718
rect 26908 36706 27412 36708
rect 26908 36654 27358 36706
rect 27410 36654 27412 36706
rect 26908 36652 27412 36654
rect 27356 36642 27412 36652
rect 28252 36594 28308 37996
rect 28364 37828 28420 37838
rect 28364 37734 28420 37772
rect 28252 36542 28254 36594
rect 28306 36542 28308 36594
rect 28252 36530 28308 36542
rect 26908 36484 26964 36494
rect 26908 36390 26964 36428
rect 27244 36482 27300 36494
rect 27244 36430 27246 36482
rect 27298 36430 27300 36482
rect 27244 35924 27300 36430
rect 27804 36260 27860 36270
rect 27244 35830 27300 35868
rect 27580 36258 27860 36260
rect 27580 36206 27806 36258
rect 27858 36206 27860 36258
rect 27580 36204 27860 36206
rect 27356 35812 27412 35822
rect 27580 35812 27636 36204
rect 27804 36194 27860 36204
rect 28364 35924 28420 35934
rect 28476 35924 28532 38220
rect 28588 38052 28644 38062
rect 28588 37958 28644 37996
rect 28700 37828 28756 38612
rect 29148 38276 29204 40908
rect 29260 40898 29316 40908
rect 29372 40516 29428 41022
rect 29260 40460 29428 40516
rect 29260 40402 29316 40460
rect 29260 40350 29262 40402
rect 29314 40350 29316 40402
rect 29260 38500 29316 40350
rect 29484 40404 29540 40414
rect 29484 40290 29540 40348
rect 29484 40238 29486 40290
rect 29538 40238 29540 40290
rect 29484 40226 29540 40238
rect 29596 38668 29652 42252
rect 30044 42196 30100 42702
rect 30044 42130 30100 42140
rect 29708 41970 29764 41982
rect 29708 41918 29710 41970
rect 29762 41918 29764 41970
rect 29708 40628 29764 41918
rect 29708 40562 29764 40572
rect 30156 41524 30212 41534
rect 30156 39284 30212 41468
rect 30268 40516 30324 43486
rect 30380 41970 30436 46844
rect 30940 43652 30996 48972
rect 31052 46786 31108 46798
rect 31052 46734 31054 46786
rect 31106 46734 31108 46786
rect 31052 46228 31108 46734
rect 31052 46162 31108 46172
rect 31052 46004 31108 46014
rect 31052 45910 31108 45948
rect 31164 45780 31220 54124
rect 31276 53956 31332 53966
rect 31276 53172 31332 53900
rect 31388 53844 31444 55134
rect 31500 55188 31556 55198
rect 31500 55094 31556 55132
rect 31500 54628 31556 54638
rect 31612 54628 31668 55244
rect 31724 55298 31780 56140
rect 31836 56130 31892 56140
rect 32508 56196 32564 56206
rect 32508 56102 32564 56140
rect 32284 56082 32340 56094
rect 32284 56030 32286 56082
rect 32338 56030 32340 56082
rect 32284 55522 32340 56030
rect 32284 55470 32286 55522
rect 32338 55470 32340 55522
rect 32284 55458 32340 55470
rect 31724 55246 31726 55298
rect 31778 55246 31780 55298
rect 31724 55234 31780 55246
rect 32284 55300 32340 55310
rect 32284 55186 32340 55244
rect 32284 55134 32286 55186
rect 32338 55134 32340 55186
rect 32284 55122 32340 55134
rect 32396 55186 32452 55198
rect 32396 55134 32398 55186
rect 32450 55134 32452 55186
rect 31500 54626 31668 54628
rect 31500 54574 31502 54626
rect 31554 54574 31668 54626
rect 31500 54572 31668 54574
rect 31500 54562 31556 54572
rect 31948 54404 32004 54414
rect 32396 54404 32452 55134
rect 32508 54404 32564 54414
rect 32396 54402 32564 54404
rect 32396 54350 32510 54402
rect 32562 54350 32564 54402
rect 32396 54348 32564 54350
rect 31948 54068 32004 54348
rect 32508 54292 32564 54348
rect 32508 54226 32564 54236
rect 31388 53778 31444 53788
rect 31724 54012 32004 54068
rect 31276 53078 31332 53116
rect 30940 43586 30996 43596
rect 31052 45724 31220 45780
rect 31276 52948 31332 52958
rect 31052 42866 31108 45724
rect 31164 44324 31220 44334
rect 31164 44230 31220 44268
rect 31276 42868 31332 52892
rect 31500 52946 31556 52958
rect 31500 52894 31502 52946
rect 31554 52894 31556 52946
rect 31500 52162 31556 52894
rect 31500 52110 31502 52162
rect 31554 52110 31556 52162
rect 31500 46788 31556 52110
rect 31724 50428 31780 54012
rect 32172 53172 32228 53182
rect 32172 52946 32228 53116
rect 32172 52894 32174 52946
rect 32226 52894 32228 52946
rect 32172 52882 32228 52894
rect 31948 52836 32004 52846
rect 31948 52742 32004 52780
rect 32508 52724 32564 52734
rect 32508 52722 32788 52724
rect 32508 52670 32510 52722
rect 32562 52670 32788 52722
rect 32508 52668 32788 52670
rect 32508 52658 32564 52668
rect 32508 52388 32564 52398
rect 32396 52276 32452 52286
rect 32396 52182 32452 52220
rect 31836 52164 31892 52174
rect 31836 52070 31892 52108
rect 32508 51602 32564 52332
rect 32732 52162 32788 52668
rect 32732 52110 32734 52162
rect 32786 52110 32788 52162
rect 32732 52098 32788 52110
rect 32508 51550 32510 51602
rect 32562 51550 32564 51602
rect 32508 51538 32564 51550
rect 32284 50820 32340 50830
rect 32284 50594 32340 50764
rect 32284 50542 32286 50594
rect 32338 50542 32340 50594
rect 32284 50428 32340 50542
rect 32508 50594 32564 50606
rect 32508 50542 32510 50594
rect 32562 50542 32564 50594
rect 31724 50372 31892 50428
rect 32284 50372 32452 50428
rect 31612 49812 31668 49822
rect 31612 49810 31780 49812
rect 31612 49758 31614 49810
rect 31666 49758 31780 49810
rect 31612 49756 31780 49758
rect 31612 49746 31668 49756
rect 31724 49028 31780 49756
rect 31724 48934 31780 48972
rect 31500 46722 31556 46732
rect 31388 46564 31444 46574
rect 31388 46470 31444 46508
rect 31724 46564 31780 46574
rect 31724 46470 31780 46508
rect 31500 45220 31556 45230
rect 31500 45126 31556 45164
rect 31724 45106 31780 45118
rect 31724 45054 31726 45106
rect 31778 45054 31780 45106
rect 31724 44546 31780 45054
rect 31724 44494 31726 44546
rect 31778 44494 31780 44546
rect 31724 44482 31780 44494
rect 31388 44436 31444 44446
rect 31388 44342 31444 44380
rect 31836 44324 31892 50372
rect 32060 49810 32116 49822
rect 32060 49758 32062 49810
rect 32114 49758 32116 49810
rect 32060 49028 32116 49758
rect 32396 49698 32452 50372
rect 32396 49646 32398 49698
rect 32450 49646 32452 49698
rect 32396 49634 32452 49646
rect 32508 49700 32564 50542
rect 32508 49634 32564 49644
rect 32732 49812 32788 49822
rect 32284 49252 32340 49262
rect 32172 49028 32228 49038
rect 32060 49026 32228 49028
rect 32060 48974 32174 49026
rect 32226 48974 32228 49026
rect 32060 48972 32228 48974
rect 31948 46786 32004 46798
rect 31948 46734 31950 46786
rect 32002 46734 32004 46786
rect 31948 46564 32004 46734
rect 31948 46498 32004 46508
rect 32060 46450 32116 46462
rect 32060 46398 32062 46450
rect 32114 46398 32116 46450
rect 31948 46228 32004 46238
rect 31948 44994 32004 46172
rect 32060 45780 32116 46398
rect 32060 45714 32116 45724
rect 31948 44942 31950 44994
rect 32002 44942 32004 44994
rect 31948 44930 32004 44942
rect 32060 44436 32116 44446
rect 31052 42814 31054 42866
rect 31106 42814 31108 42866
rect 31052 42802 31108 42814
rect 31164 42812 31332 42868
rect 31612 44268 31892 44324
rect 31948 44324 32004 44334
rect 30940 42754 30996 42766
rect 30940 42702 30942 42754
rect 30994 42702 30996 42754
rect 30380 41918 30382 41970
rect 30434 41918 30436 41970
rect 30380 41906 30436 41918
rect 30492 42642 30548 42654
rect 30492 42590 30494 42642
rect 30546 42590 30548 42642
rect 30492 41860 30548 42590
rect 30940 42532 30996 42702
rect 30940 42466 30996 42476
rect 31164 42308 31220 42812
rect 30492 41794 30548 41804
rect 30716 42252 31220 42308
rect 31276 42644 31332 42654
rect 30268 40450 30324 40460
rect 30156 39218 30212 39228
rect 30380 39060 30436 39070
rect 30380 38946 30436 39004
rect 30380 38894 30382 38946
rect 30434 38894 30436 38946
rect 30380 38882 30436 38894
rect 30044 38836 30100 38846
rect 29260 38434 29316 38444
rect 29484 38612 29652 38668
rect 29932 38724 29988 38762
rect 30044 38742 30100 38780
rect 30604 38834 30660 38846
rect 30604 38782 30606 38834
rect 30658 38782 30660 38834
rect 29932 38658 29988 38668
rect 29260 38276 29316 38286
rect 29148 38274 29316 38276
rect 29148 38222 29262 38274
rect 29314 38222 29316 38274
rect 29148 38220 29316 38222
rect 29260 38210 29316 38220
rect 28700 37762 28756 37772
rect 29148 38052 29204 38062
rect 29148 37266 29204 37996
rect 29260 37940 29316 37950
rect 29260 37846 29316 37884
rect 29372 37938 29428 37950
rect 29372 37886 29374 37938
rect 29426 37886 29428 37938
rect 29148 37214 29150 37266
rect 29202 37214 29204 37266
rect 29148 37202 29204 37214
rect 29372 37268 29428 37886
rect 27356 35810 27636 35812
rect 27356 35758 27358 35810
rect 27410 35758 27636 35810
rect 27356 35756 27636 35758
rect 27916 35922 28532 35924
rect 27916 35870 28366 35922
rect 28418 35870 28532 35922
rect 27916 35868 28532 35870
rect 25676 35588 25732 35598
rect 25564 35586 25732 35588
rect 25564 35534 25678 35586
rect 25730 35534 25732 35586
rect 25564 35532 25732 35534
rect 25452 34018 25508 35532
rect 25676 35364 25732 35532
rect 27356 35588 27412 35756
rect 27356 35522 27412 35532
rect 25676 35298 25732 35308
rect 27916 35028 27972 35868
rect 28364 35858 28420 35868
rect 29372 35140 29428 37212
rect 29260 35084 29428 35140
rect 27916 34934 27972 34972
rect 29148 35028 29204 35038
rect 28364 34690 28420 34702
rect 28364 34638 28366 34690
rect 28418 34638 28420 34690
rect 28364 34468 28420 34638
rect 28252 34412 28364 34468
rect 25452 33966 25454 34018
rect 25506 33966 25508 34018
rect 25452 33954 25508 33966
rect 27580 34020 27636 34030
rect 27580 34018 27972 34020
rect 27580 33966 27582 34018
rect 27634 33966 27972 34018
rect 27580 33964 27972 33966
rect 27580 33954 27636 33964
rect 25116 33460 25172 33470
rect 24668 33124 24724 33134
rect 24668 33030 24724 33068
rect 25116 33124 25172 33404
rect 27916 33458 27972 33964
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33394 27972 33406
rect 28140 33348 28196 33358
rect 28140 33254 28196 33292
rect 25788 33236 25844 33246
rect 25788 33142 25844 33180
rect 27804 33234 27860 33246
rect 27804 33182 27806 33234
rect 27858 33182 27860 33234
rect 25452 33124 25508 33134
rect 25116 33122 25508 33124
rect 25116 33070 25118 33122
rect 25170 33070 25454 33122
rect 25506 33070 25508 33122
rect 25116 33068 25508 33070
rect 24108 32734 24110 32786
rect 24162 32734 24164 32786
rect 24108 31892 24164 32734
rect 24108 31826 24164 31836
rect 24220 32786 24500 32788
rect 24220 32734 24446 32786
rect 24498 32734 24500 32786
rect 24220 32732 24500 32734
rect 23884 31726 23886 31778
rect 23938 31726 23940 31778
rect 22988 30370 23044 30380
rect 23100 30716 23268 30772
rect 23436 30996 23492 31006
rect 21868 29598 21870 29650
rect 21922 29598 21924 29650
rect 21868 29586 21924 29598
rect 22316 29708 22708 29764
rect 22764 29988 22820 29998
rect 22876 29988 22932 29998
rect 22820 29986 22932 29988
rect 22820 29934 22878 29986
rect 22930 29934 22932 29986
rect 22820 29932 22932 29934
rect 22316 29650 22372 29708
rect 22316 29598 22318 29650
rect 22370 29598 22372 29650
rect 21532 29540 21588 29550
rect 21532 29446 21588 29484
rect 21644 29538 21700 29550
rect 21644 29486 21646 29538
rect 21698 29486 21700 29538
rect 21084 29374 21086 29426
rect 21138 29374 21140 29426
rect 21084 29362 21140 29374
rect 20188 27468 20356 27524
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 25788 19908 25844
rect 19180 25676 19796 25732
rect 19740 25618 19796 25676
rect 19740 25566 19742 25618
rect 19794 25566 19796 25618
rect 19740 25554 19796 25566
rect 19852 25396 19908 25788
rect 19628 25340 19908 25396
rect 19068 24948 19124 24958
rect 19012 24946 19124 24948
rect 19012 24894 19070 24946
rect 19122 24894 19124 24946
rect 19012 24892 19124 24894
rect 18956 24854 19012 24892
rect 19068 24882 19124 24892
rect 19404 24948 19460 24958
rect 19404 24050 19460 24892
rect 19628 24724 19684 25340
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19740 24724 19796 24734
rect 19628 24722 19796 24724
rect 19628 24670 19742 24722
rect 19794 24670 19796 24722
rect 19628 24668 19796 24670
rect 19740 24658 19796 24668
rect 19404 23998 19406 24050
rect 19458 23998 19460 24050
rect 18732 23650 18788 23660
rect 18956 23938 19012 23950
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23828 19012 23886
rect 17500 23156 17556 23166
rect 16828 23154 17556 23156
rect 16828 23102 16830 23154
rect 16882 23102 17502 23154
rect 17554 23102 17556 23154
rect 16828 23100 17556 23102
rect 16828 21812 16884 23100
rect 17500 23090 17556 23100
rect 18956 22596 19012 23772
rect 18956 22530 19012 22540
rect 16716 21756 16884 21812
rect 18620 21812 18676 21822
rect 14700 20914 15092 20916
rect 14700 20862 14702 20914
rect 14754 20862 15092 20914
rect 14700 20860 15092 20862
rect 14700 20850 14756 20860
rect 15036 20802 15092 20860
rect 15036 20750 15038 20802
rect 15090 20750 15092 20802
rect 15036 20188 15092 20750
rect 15820 20692 15876 20702
rect 15820 20598 15876 20636
rect 14476 20132 15092 20188
rect 14476 19234 14532 20132
rect 15036 20066 15092 20076
rect 16716 20132 16772 21756
rect 18620 21718 18676 21756
rect 19292 21812 19348 21822
rect 19292 21718 19348 21756
rect 18284 21698 18340 21710
rect 18284 21646 18286 21698
rect 18338 21646 18340 21698
rect 17948 20916 18004 20926
rect 16716 20066 16772 20076
rect 17724 20914 18004 20916
rect 17724 20862 17950 20914
rect 18002 20862 18004 20914
rect 17724 20860 18004 20862
rect 17724 20020 17780 20860
rect 17948 20850 18004 20860
rect 18284 20804 18340 21646
rect 18956 21700 19012 21710
rect 19012 21644 19236 21700
rect 18956 21606 19012 21644
rect 18172 20802 18340 20804
rect 18172 20750 18286 20802
rect 18338 20750 18340 20802
rect 18172 20748 18340 20750
rect 18060 20132 18116 20142
rect 17724 19954 17780 19964
rect 17836 20076 18060 20132
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19170 14532 19182
rect 17276 19346 17332 19358
rect 17276 19294 17278 19346
rect 17330 19294 17332 19346
rect 15148 19122 15204 19134
rect 15148 19070 15150 19122
rect 15202 19070 15204 19122
rect 15148 18452 15204 19070
rect 15148 18386 15204 18396
rect 17276 19012 17332 19294
rect 17836 19346 17892 20076
rect 18060 20038 18116 20076
rect 17836 19294 17838 19346
rect 17890 19294 17892 19346
rect 17836 19282 17892 19294
rect 18172 19012 18228 20748
rect 18284 20738 18340 20748
rect 18620 20916 18676 20926
rect 18620 20802 18676 20860
rect 18620 20750 18622 20802
rect 18674 20750 18676 20802
rect 18620 20738 18676 20750
rect 18732 20802 18788 20814
rect 18732 20750 18734 20802
rect 18786 20750 18788 20802
rect 18396 20692 18452 20702
rect 18396 20598 18452 20636
rect 18508 20580 18564 20590
rect 18508 20468 18564 20524
rect 18396 20412 18564 20468
rect 18396 20132 18452 20412
rect 18732 20356 18788 20750
rect 18508 20300 18788 20356
rect 18508 20242 18564 20300
rect 18508 20190 18510 20242
rect 18562 20190 18564 20242
rect 18508 20178 18564 20190
rect 18284 20130 18452 20132
rect 18284 20078 18398 20130
rect 18450 20078 18452 20130
rect 18284 20076 18452 20078
rect 18284 19234 18340 20076
rect 18396 20066 18452 20076
rect 18620 20020 18676 20030
rect 18676 19964 18788 20020
rect 18620 19926 18676 19964
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 18284 19170 18340 19182
rect 14700 17444 14756 17454
rect 14700 16994 14756 17388
rect 16828 17108 16884 17118
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 16604 16996 16660 17006
rect 11004 16258 11060 16268
rect 14028 16882 14084 16894
rect 14028 16830 14030 16882
rect 14082 16830 14084 16882
rect 5852 11666 5908 11676
rect 14028 16100 14084 16830
rect 14028 13746 14084 16044
rect 15820 16772 15876 16782
rect 15820 16100 15876 16716
rect 16604 16210 16660 16940
rect 16828 16770 16884 17052
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 16604 16158 16606 16210
rect 16658 16158 16660 16210
rect 16604 16146 16660 16158
rect 15820 16006 15876 16044
rect 17276 14644 17332 18956
rect 17948 18956 18228 19012
rect 18396 19010 18452 19022
rect 18396 18958 18398 19010
rect 18450 18958 18452 19010
rect 17948 18452 18004 18956
rect 18396 18788 18452 18958
rect 18508 19012 18564 19022
rect 18508 18918 18564 18956
rect 18396 18732 18564 18788
rect 18508 18562 18564 18732
rect 18508 18510 18510 18562
rect 18562 18510 18564 18562
rect 18508 18498 18564 18510
rect 17388 18450 18004 18452
rect 17388 18398 17950 18450
rect 18002 18398 18004 18450
rect 17388 18396 18004 18398
rect 17388 17666 17444 18396
rect 17948 18386 18004 18396
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 18284 18452 18340 18462
rect 18284 18358 18340 18396
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 17388 17332 17444 17614
rect 17948 17668 18004 17678
rect 18396 17668 18452 17678
rect 17948 17666 18452 17668
rect 17948 17614 17950 17666
rect 18002 17614 18398 17666
rect 18450 17614 18452 17666
rect 17948 17612 18452 17614
rect 17948 17602 18004 17612
rect 18396 17602 18452 17612
rect 17724 17554 17780 17566
rect 17724 17502 17726 17554
rect 17778 17502 17780 17554
rect 17500 17444 17556 17454
rect 17500 17350 17556 17388
rect 17388 17266 17444 17276
rect 17724 17220 17780 17502
rect 18284 17444 18340 17482
rect 18284 17378 18340 17388
rect 18508 17442 18564 17454
rect 18508 17390 18510 17442
rect 18562 17390 18564 17442
rect 18396 17332 18452 17342
rect 17724 17154 17780 17164
rect 18284 17220 18340 17230
rect 18060 17108 18116 17118
rect 17612 16884 17668 16894
rect 17612 16790 17668 16828
rect 17276 14578 17332 14588
rect 14700 13972 14756 13982
rect 14700 13858 14756 13916
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 16828 13860 16884 13870
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13636 14084 13694
rect 14028 11396 14084 13580
rect 16828 13634 16884 13804
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 16828 13570 16884 13582
rect 17500 13636 17556 13646
rect 17500 13542 17556 13580
rect 17836 13188 17892 13198
rect 17836 13094 17892 13132
rect 17948 12852 18004 12862
rect 17948 12758 18004 12796
rect 17836 12740 17892 12750
rect 17612 12684 17836 12740
rect 17276 11508 17332 11518
rect 17276 11414 17332 11452
rect 14364 11396 14420 11406
rect 14028 11394 14420 11396
rect 14028 11342 14366 11394
rect 14418 11342 14420 11394
rect 14028 11340 14420 11342
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 14364 10164 14420 11340
rect 15148 11284 15204 11294
rect 15148 11282 15876 11284
rect 15148 11230 15150 11282
rect 15202 11230 15876 11282
rect 15148 11228 15876 11230
rect 15148 11218 15204 11228
rect 15820 10834 15876 11228
rect 15820 10782 15822 10834
rect 15874 10782 15876 10834
rect 15820 10770 15876 10782
rect 15932 11172 15988 11182
rect 15932 10722 15988 11116
rect 15932 10670 15934 10722
rect 15986 10670 15988 10722
rect 15932 10658 15988 10670
rect 14028 9044 14084 9054
rect 14364 9044 14420 10108
rect 17500 10164 17556 10174
rect 15932 9940 15988 9950
rect 15932 9846 15988 9884
rect 16828 9716 16884 9726
rect 14700 9604 14756 9614
rect 14700 9154 14756 9548
rect 15820 9604 15876 9614
rect 15820 9510 15876 9548
rect 14700 9102 14702 9154
rect 14754 9102 14756 9154
rect 14700 9090 14756 9102
rect 14028 9042 14420 9044
rect 14028 8990 14030 9042
rect 14082 8990 14420 9042
rect 14028 8988 14420 8990
rect 14028 8978 14084 8988
rect 16828 8930 16884 9660
rect 16828 8878 16830 8930
rect 16882 8878 16884 8930
rect 16828 8866 16884 8878
rect 17500 9266 17556 10108
rect 17612 9938 17668 12684
rect 17836 12646 17892 12684
rect 17724 11396 17780 11406
rect 17724 11170 17780 11340
rect 17724 11118 17726 11170
rect 17778 11118 17780 11170
rect 17724 10164 17780 11118
rect 18060 10722 18116 17052
rect 18284 17106 18340 17164
rect 18284 17054 18286 17106
rect 18338 17054 18340 17106
rect 18284 17042 18340 17054
rect 18396 16882 18452 17276
rect 18508 17108 18564 17390
rect 18508 17042 18564 17052
rect 18620 16996 18676 17006
rect 18620 16902 18676 16940
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18396 16818 18452 16830
rect 18732 16772 18788 19964
rect 18956 20018 19012 20030
rect 18956 19966 18958 20018
rect 19010 19966 19012 20018
rect 18956 19234 19012 19966
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 17666 19012 19182
rect 19068 18676 19124 18686
rect 19068 18452 19124 18620
rect 19068 18358 19124 18396
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18956 17556 19012 17614
rect 18956 17490 19012 17500
rect 19180 17666 19236 21644
rect 19292 20916 19348 20926
rect 19292 20822 19348 20860
rect 19404 20356 19460 23998
rect 19852 23938 19908 23950
rect 19852 23886 19854 23938
rect 19906 23886 19908 23938
rect 19852 23716 19908 23886
rect 19852 23650 19908 23660
rect 20300 23938 20356 27468
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19740 23042 19796 23054
rect 19740 22990 19742 23042
rect 19794 22990 19796 23042
rect 19740 22596 19796 22990
rect 19740 22530 19796 22540
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19964 21812 20020 21822
rect 19964 21718 20020 21756
rect 19628 21698 19684 21710
rect 19628 21646 19630 21698
rect 19682 21646 19684 21698
rect 19628 20580 19684 21646
rect 20076 21700 20132 21710
rect 20076 20802 20132 21644
rect 20300 20916 20356 23886
rect 20300 20850 20356 20860
rect 20412 27468 20692 27524
rect 20748 29314 20804 29326
rect 20748 29262 20750 29314
rect 20802 29262 20804 29314
rect 20748 29204 20804 29262
rect 21532 29316 21588 29326
rect 21532 29222 21588 29260
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 20076 20738 20132 20750
rect 19628 20514 19684 20524
rect 20300 20578 20356 20590
rect 20300 20526 20302 20578
rect 20354 20526 20356 20578
rect 19292 20300 19460 20356
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 19348 19348 20300
rect 19404 20132 19460 20142
rect 19404 20018 19460 20076
rect 20188 20132 20244 20142
rect 20300 20132 20356 20526
rect 20188 20130 20356 20132
rect 20188 20078 20190 20130
rect 20242 20078 20356 20130
rect 20188 20076 20356 20078
rect 20188 20066 20244 20076
rect 19404 19966 19406 20018
rect 19458 19966 19460 20018
rect 19404 19954 19460 19966
rect 19292 18676 19348 19292
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19292 18610 19348 18620
rect 19180 17614 19182 17666
rect 19234 17614 19236 17666
rect 19180 17444 19236 17614
rect 19852 17668 19908 17678
rect 19852 17574 19908 17612
rect 19180 17378 19236 17388
rect 19292 17442 19348 17454
rect 19292 17390 19294 17442
rect 19346 17390 19348 17442
rect 18844 16996 18900 17006
rect 19068 16996 19124 17006
rect 19292 16996 19348 17390
rect 18844 16994 19012 16996
rect 18844 16942 18846 16994
rect 18898 16942 19012 16994
rect 18844 16940 19012 16942
rect 18844 16930 18900 16940
rect 18620 16716 18788 16772
rect 18956 16772 19012 16940
rect 19068 16994 19348 16996
rect 19068 16942 19070 16994
rect 19122 16942 19348 16994
rect 19068 16940 19348 16942
rect 19404 17442 19460 17454
rect 19404 17390 19406 17442
rect 19458 17390 19460 17442
rect 19068 16930 19124 16940
rect 18956 16716 19124 16772
rect 18284 14644 18340 14654
rect 18284 14550 18340 14588
rect 18508 14532 18564 14542
rect 18508 14438 18564 14476
rect 18508 13860 18564 13870
rect 18284 13746 18340 13758
rect 18284 13694 18286 13746
rect 18338 13694 18340 13746
rect 18284 13188 18340 13694
rect 18284 13122 18340 13132
rect 18396 12962 18452 12974
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18284 12178 18340 12190
rect 18284 12126 18286 12178
rect 18338 12126 18340 12178
rect 18284 11956 18340 12126
rect 18284 11890 18340 11900
rect 18284 11508 18340 11518
rect 18396 11508 18452 12910
rect 18340 11452 18452 11508
rect 18284 11442 18340 11452
rect 18060 10670 18062 10722
rect 18114 10670 18116 10722
rect 18060 10658 18116 10670
rect 18172 10834 18228 10846
rect 18172 10782 18174 10834
rect 18226 10782 18228 10834
rect 17724 10098 17780 10108
rect 17836 10610 17892 10622
rect 17836 10558 17838 10610
rect 17890 10558 17892 10610
rect 17612 9886 17614 9938
rect 17666 9886 17668 9938
rect 17612 9828 17668 9886
rect 17612 9762 17668 9772
rect 17836 9716 17892 10558
rect 17948 10052 18004 10062
rect 18172 10052 18228 10782
rect 18508 10836 18564 13804
rect 18620 12962 18676 16716
rect 18732 16212 18788 16222
rect 18732 15148 18788 16156
rect 19068 15988 19124 16716
rect 19404 16212 19460 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16884 19684 16894
rect 19852 16884 19908 16894
rect 19684 16882 19908 16884
rect 19684 16830 19854 16882
rect 19906 16830 19908 16882
rect 19684 16828 19908 16830
rect 19628 16790 19684 16828
rect 19404 16146 19460 16156
rect 19740 16210 19796 16828
rect 19852 16818 19908 16828
rect 19740 16158 19742 16210
rect 19794 16158 19796 16210
rect 19740 16146 19796 16158
rect 20412 16212 20468 27468
rect 20748 25172 20804 29148
rect 21644 29204 21700 29486
rect 22092 29540 22148 29550
rect 22092 29446 22148 29484
rect 21644 29138 21700 29148
rect 22316 27748 22372 29598
rect 22428 29540 22484 29550
rect 22428 29446 22484 29484
rect 22428 27748 22484 27758
rect 22316 27746 22484 27748
rect 22316 27694 22430 27746
rect 22482 27694 22484 27746
rect 22316 27692 22484 27694
rect 22428 27682 22484 27692
rect 22316 26516 22372 26526
rect 22652 26516 22708 26526
rect 22372 26514 22708 26516
rect 22372 26462 22654 26514
rect 22706 26462 22708 26514
rect 22372 26460 22708 26462
rect 22316 26422 22372 26460
rect 22652 26450 22708 26460
rect 21420 25508 21476 25518
rect 21420 25506 21700 25508
rect 21420 25454 21422 25506
rect 21474 25454 21700 25506
rect 21420 25452 21700 25454
rect 21420 25442 21476 25452
rect 20748 25106 20804 25116
rect 21532 25282 21588 25294
rect 21532 25230 21534 25282
rect 21586 25230 21588 25282
rect 21532 24948 21588 25230
rect 20524 24892 21588 24948
rect 20524 24834 20580 24892
rect 20524 24782 20526 24834
rect 20578 24782 20580 24834
rect 20524 24770 20580 24782
rect 21644 23940 21700 25452
rect 21756 25394 21812 25406
rect 21756 25342 21758 25394
rect 21810 25342 21812 25394
rect 21756 25284 21812 25342
rect 21980 25396 22036 25406
rect 21980 25394 22372 25396
rect 21980 25342 21982 25394
rect 22034 25342 22372 25394
rect 21980 25340 22372 25342
rect 21980 25330 22036 25340
rect 21756 25218 21812 25228
rect 22316 24050 22372 25340
rect 22316 23998 22318 24050
rect 22370 23998 22372 24050
rect 22316 23986 22372 23998
rect 22540 25284 22596 25294
rect 21644 23874 21700 23884
rect 22204 23940 22260 23950
rect 20748 23716 20804 23726
rect 20748 22708 20804 23660
rect 21980 23714 22036 23726
rect 21980 23662 21982 23714
rect 22034 23662 22036 23714
rect 21980 23492 22036 23662
rect 21980 23426 22036 23436
rect 22204 23156 22260 23884
rect 22428 23714 22484 23726
rect 22428 23662 22430 23714
rect 22482 23662 22484 23714
rect 22428 23604 22484 23662
rect 22428 23538 22484 23548
rect 22540 23268 22596 25228
rect 22764 24836 22820 29932
rect 22876 29922 22932 29932
rect 22876 29652 22932 29662
rect 22876 29558 22932 29596
rect 22876 27860 22932 27870
rect 22876 26964 22932 27804
rect 22876 26898 22932 26908
rect 22764 24770 22820 24780
rect 22652 24724 22708 24734
rect 22652 24610 22708 24668
rect 22988 24612 23044 24622
rect 22652 24558 22654 24610
rect 22706 24558 22708 24610
rect 22652 24546 22708 24558
rect 22764 24610 23044 24612
rect 22764 24558 22990 24610
rect 23042 24558 23044 24610
rect 22764 24556 23044 24558
rect 22428 23212 22596 23268
rect 22652 23714 22708 23726
rect 22652 23662 22654 23714
rect 22706 23662 22708 23714
rect 22652 23492 22708 23662
rect 22764 23604 22820 24556
rect 22988 24546 23044 24556
rect 22764 23538 22820 23548
rect 22316 23156 22372 23166
rect 22204 23154 22372 23156
rect 22204 23102 22318 23154
rect 22370 23102 22372 23154
rect 22204 23100 22372 23102
rect 22316 23090 22372 23100
rect 22428 22932 22484 23212
rect 20748 22642 20804 22652
rect 22316 22876 22484 22932
rect 22540 23042 22596 23054
rect 22540 22990 22542 23042
rect 22594 22990 22596 23042
rect 20524 21700 20580 21710
rect 20524 20802 20580 21644
rect 21756 21588 21812 21598
rect 21756 21494 21812 21532
rect 20524 20750 20526 20802
rect 20578 20750 20580 20802
rect 20524 20738 20580 20750
rect 20748 20692 20804 20702
rect 20748 20598 20804 20636
rect 21980 20692 22036 20702
rect 21980 20598 22036 20636
rect 21868 20580 21924 20590
rect 21868 20188 21924 20524
rect 21756 20132 21924 20188
rect 22092 20578 22148 20590
rect 22092 20526 22094 20578
rect 22146 20526 22148 20578
rect 21756 18674 21812 20132
rect 22092 19908 22148 20526
rect 22316 20580 22372 22876
rect 22428 21700 22484 21710
rect 22540 21700 22596 22990
rect 22428 21698 22596 21700
rect 22428 21646 22430 21698
rect 22482 21646 22596 21698
rect 22428 21644 22596 21646
rect 22428 21634 22484 21644
rect 22540 20804 22596 20814
rect 22652 20804 22708 23436
rect 22764 23268 22820 23278
rect 22764 21700 22820 23212
rect 22988 23156 23044 23166
rect 22988 23062 23044 23100
rect 22764 21634 22820 21644
rect 22876 20804 22932 20814
rect 22540 20802 22932 20804
rect 22540 20750 22542 20802
rect 22594 20750 22878 20802
rect 22930 20750 22932 20802
rect 22540 20748 22932 20750
rect 22540 20738 22596 20748
rect 22876 20738 22932 20748
rect 23100 20580 23156 30716
rect 23212 29652 23268 29662
rect 23212 29558 23268 29596
rect 23436 29540 23492 30940
rect 23884 30212 23940 31726
rect 24108 31220 24164 31230
rect 24220 31220 24276 32732
rect 24444 32722 24500 32732
rect 24668 31668 24724 31678
rect 24668 31666 25060 31668
rect 24668 31614 24670 31666
rect 24722 31614 25060 31666
rect 24668 31612 25060 31614
rect 24668 31602 24724 31612
rect 24108 31218 24276 31220
rect 24108 31166 24110 31218
rect 24162 31166 24276 31218
rect 24108 31164 24276 31166
rect 24108 31154 24164 31164
rect 23996 30996 24052 31006
rect 23996 30902 24052 30940
rect 24332 30996 24388 31006
rect 24332 30994 24612 30996
rect 24332 30942 24334 30994
rect 24386 30942 24612 30994
rect 24332 30940 24612 30942
rect 24332 30930 24388 30940
rect 23996 30212 24052 30222
rect 23884 30156 23996 30212
rect 23996 30146 24052 30156
rect 24220 30100 24276 30110
rect 24276 30044 24388 30100
rect 24220 30006 24276 30044
rect 24332 29650 24388 30044
rect 24556 30098 24612 30940
rect 25004 30322 25060 31612
rect 25004 30270 25006 30322
rect 25058 30270 25060 30322
rect 25004 30258 25060 30270
rect 24556 30046 24558 30098
rect 24610 30046 24612 30098
rect 24556 30034 24612 30046
rect 24780 30098 24836 30110
rect 24780 30046 24782 30098
rect 24834 30046 24836 30098
rect 24444 29988 24500 29998
rect 24444 29894 24500 29932
rect 24332 29598 24334 29650
rect 24386 29598 24388 29650
rect 24332 29586 24388 29598
rect 23660 29540 23716 29550
rect 23436 29484 23660 29540
rect 23660 29446 23716 29484
rect 23996 29426 24052 29438
rect 23996 29374 23998 29426
rect 24050 29374 24052 29426
rect 23996 29316 24052 29374
rect 24556 29426 24612 29438
rect 24556 29374 24558 29426
rect 24610 29374 24612 29426
rect 24556 29316 24612 29374
rect 24780 29428 24836 30046
rect 24780 29362 24836 29372
rect 23996 29260 24612 29316
rect 23436 27748 23492 27758
rect 23324 26516 23380 26526
rect 23212 26178 23268 26190
rect 23212 26126 23214 26178
rect 23266 26126 23268 26178
rect 23212 25396 23268 26126
rect 23324 25618 23380 26460
rect 23436 25956 23492 27692
rect 24556 27298 24612 29260
rect 24556 27246 24558 27298
rect 24610 27246 24612 27298
rect 24556 27234 24612 27246
rect 23996 26964 24052 26974
rect 23772 26516 23828 26526
rect 23772 26290 23828 26460
rect 23772 26238 23774 26290
rect 23826 26238 23828 26290
rect 23772 26226 23828 26238
rect 23436 25890 23492 25900
rect 23324 25566 23326 25618
rect 23378 25566 23380 25618
rect 23324 25554 23380 25566
rect 23884 25508 23940 25518
rect 23884 25414 23940 25452
rect 23212 25330 23268 25340
rect 23436 25284 23492 25294
rect 23324 25228 23436 25284
rect 22316 20524 22596 20580
rect 22316 19908 22372 19918
rect 22092 19906 22484 19908
rect 22092 19854 22318 19906
rect 22370 19854 22484 19906
rect 22092 19852 22484 19854
rect 22316 19842 22372 19852
rect 21756 18622 21758 18674
rect 21810 18622 21812 18674
rect 21756 18610 21812 18622
rect 21980 18452 22036 18462
rect 21980 18450 22260 18452
rect 21980 18398 21982 18450
rect 22034 18398 22260 18450
rect 21980 18396 22260 18398
rect 21980 18386 22036 18396
rect 21868 18338 21924 18350
rect 21868 18286 21870 18338
rect 21922 18286 21924 18338
rect 21644 17780 21700 17790
rect 21196 17666 21252 17678
rect 21196 17614 21198 17666
rect 21250 17614 21252 17666
rect 21196 17444 21252 17614
rect 21644 17666 21700 17724
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 17602 21700 17614
rect 21868 17666 21924 18286
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17602 21924 17614
rect 21196 17378 21252 17388
rect 21420 17442 21476 17454
rect 21420 17390 21422 17442
rect 21474 17390 21476 17442
rect 21420 17108 21476 17390
rect 20636 17052 21476 17108
rect 20636 16994 20692 17052
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 22204 16884 22260 18396
rect 22316 18450 22372 18462
rect 22316 18398 22318 18450
rect 22370 18398 22372 18450
rect 22316 18338 22372 18398
rect 22316 18286 22318 18338
rect 22370 18286 22372 18338
rect 22316 18274 22372 18286
rect 22428 18116 22484 19852
rect 22540 18340 22596 20524
rect 22876 20524 23156 20580
rect 23212 24836 23268 24846
rect 22540 18274 22596 18284
rect 22764 18338 22820 18350
rect 22764 18286 22766 18338
rect 22818 18286 22820 18338
rect 22428 18060 22708 18116
rect 22316 17780 22372 17790
rect 22316 17686 22372 17724
rect 22652 17220 22708 18060
rect 22764 17556 22820 18286
rect 22876 18228 22932 20524
rect 23212 19460 23268 24780
rect 23324 23492 23380 25228
rect 23436 25218 23492 25228
rect 23436 24724 23492 24734
rect 23436 24630 23492 24668
rect 23324 23380 23380 23436
rect 23996 24610 24052 26908
rect 24668 26962 24724 26974
rect 24668 26910 24670 26962
rect 24722 26910 24724 26962
rect 24556 26852 24612 26862
rect 24220 26290 24276 26302
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 24220 26180 24276 26238
rect 24220 26114 24276 26124
rect 24332 26180 24388 26190
rect 24332 26178 24500 26180
rect 24332 26126 24334 26178
rect 24386 26126 24500 26178
rect 24332 26124 24500 26126
rect 24332 26114 24388 26124
rect 24444 25956 24500 26124
rect 24108 25732 24164 25742
rect 24108 25394 24164 25676
rect 24220 25508 24276 25518
rect 24220 25414 24276 25452
rect 24108 25342 24110 25394
rect 24162 25342 24164 25394
rect 24108 25330 24164 25342
rect 23996 24558 23998 24610
rect 24050 24558 24052 24610
rect 23436 23380 23492 23390
rect 23996 23380 24052 24558
rect 24332 23826 24388 23838
rect 24332 23774 24334 23826
rect 24386 23774 24388 23826
rect 24332 23492 24388 23774
rect 24332 23426 24388 23436
rect 23324 23378 23716 23380
rect 23324 23326 23438 23378
rect 23490 23326 23716 23378
rect 23324 23324 23716 23326
rect 23436 23314 23492 23324
rect 23660 23154 23716 23324
rect 23660 23102 23662 23154
rect 23714 23102 23716 23154
rect 23660 23090 23716 23102
rect 23884 22260 23940 22270
rect 23884 22166 23940 22204
rect 23996 21588 24052 23324
rect 24332 23268 24388 23278
rect 24444 23268 24500 25900
rect 24556 25732 24612 26796
rect 24668 26068 24724 26910
rect 25116 26908 25172 33068
rect 25452 33058 25508 33068
rect 27580 33124 27636 33134
rect 27804 33124 27860 33182
rect 28252 33236 28308 34412
rect 28364 34402 28420 34412
rect 29148 34354 29204 34972
rect 29148 34302 29150 34354
rect 29202 34302 29204 34354
rect 29148 34290 29204 34302
rect 28364 34132 28420 34142
rect 28364 34130 28532 34132
rect 28364 34078 28366 34130
rect 28418 34078 28532 34130
rect 28364 34076 28532 34078
rect 28364 34066 28420 34076
rect 28364 33684 28420 33694
rect 28364 33346 28420 33628
rect 28364 33294 28366 33346
rect 28418 33294 28420 33346
rect 28364 33282 28420 33294
rect 28252 33170 28308 33180
rect 27580 33122 27804 33124
rect 27580 33070 27582 33122
rect 27634 33070 27804 33122
rect 27580 33068 27804 33070
rect 27580 33058 27636 33068
rect 27804 33058 27860 33068
rect 28476 32452 28532 34076
rect 28700 34130 28756 34142
rect 28700 34078 28702 34130
rect 28754 34078 28756 34130
rect 28700 33124 28756 34078
rect 28924 34132 28980 34142
rect 29260 34132 29316 35084
rect 29372 34692 29428 34702
rect 29372 34598 29428 34636
rect 28924 34130 29316 34132
rect 28924 34078 28926 34130
rect 28978 34078 29316 34130
rect 28924 34076 29316 34078
rect 28812 34018 28868 34030
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33684 28868 33966
rect 28812 33618 28868 33628
rect 28924 33348 28980 34076
rect 29484 33460 29540 38612
rect 30268 38610 30324 38622
rect 30268 38558 30270 38610
rect 30322 38558 30324 38610
rect 30156 37826 30212 37838
rect 30156 37774 30158 37826
rect 30210 37774 30212 37826
rect 30156 37156 30212 37774
rect 30268 37380 30324 38558
rect 30492 38276 30548 38286
rect 30604 38276 30660 38782
rect 30492 38274 30660 38276
rect 30492 38222 30494 38274
rect 30546 38222 30660 38274
rect 30492 38220 30660 38222
rect 30492 38210 30548 38220
rect 30604 37940 30660 37950
rect 30604 37846 30660 37884
rect 30268 37314 30324 37324
rect 30492 37826 30548 37838
rect 30492 37774 30494 37826
rect 30546 37774 30548 37826
rect 30492 37156 30548 37774
rect 30716 37490 30772 42252
rect 31164 40516 31220 40526
rect 31164 40290 31220 40460
rect 31276 40404 31332 42588
rect 31388 40404 31444 40414
rect 31276 40402 31444 40404
rect 31276 40350 31390 40402
rect 31442 40350 31444 40402
rect 31276 40348 31444 40350
rect 31388 40338 31444 40348
rect 31164 40238 31166 40290
rect 31218 40238 31220 40290
rect 31164 40226 31220 40238
rect 31276 39618 31332 39630
rect 31276 39566 31278 39618
rect 31330 39566 31332 39618
rect 30940 39396 30996 39406
rect 30940 38836 30996 39340
rect 31276 39060 31332 39566
rect 31276 38994 31332 39004
rect 31500 39618 31556 39630
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 30828 38612 30884 38622
rect 30828 38518 30884 38556
rect 30828 37828 30884 37838
rect 30828 37734 30884 37772
rect 30716 37438 30718 37490
rect 30770 37438 30772 37490
rect 30716 37426 30772 37438
rect 30156 37100 30548 37156
rect 29708 35700 29764 35710
rect 29708 35026 29764 35644
rect 30156 35140 30212 37100
rect 30716 36596 30772 36606
rect 30940 36596 30996 38780
rect 31276 38050 31332 38062
rect 31276 37998 31278 38050
rect 31330 37998 31332 38050
rect 31276 37492 31332 37998
rect 31276 37266 31332 37436
rect 31500 37940 31556 39566
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 37202 31332 37214
rect 31388 37380 31444 37390
rect 30716 36594 30996 36596
rect 30716 36542 30718 36594
rect 30770 36542 30996 36594
rect 30716 36540 30996 36542
rect 31052 37042 31108 37054
rect 31052 36990 31054 37042
rect 31106 36990 31108 37042
rect 30492 35700 30548 35710
rect 30492 35606 30548 35644
rect 30156 35084 30324 35140
rect 29708 34974 29710 35026
rect 29762 34974 29764 35026
rect 29708 34962 29764 34974
rect 29820 34916 29876 34926
rect 30156 34916 30212 34926
rect 29820 34822 29876 34860
rect 29932 34914 30212 34916
rect 29932 34862 30158 34914
rect 30210 34862 30212 34914
rect 29932 34860 30212 34862
rect 29596 34690 29652 34702
rect 29596 34638 29598 34690
rect 29650 34638 29652 34690
rect 29596 34244 29652 34638
rect 29596 34178 29652 34188
rect 29820 34356 29876 34366
rect 29932 34356 29988 34860
rect 30156 34850 30212 34860
rect 29820 34354 29988 34356
rect 29820 34302 29822 34354
rect 29874 34302 29988 34354
rect 29820 34300 29988 34302
rect 30044 34692 30100 34702
rect 30268 34692 30324 35084
rect 30044 34354 30100 34636
rect 30044 34302 30046 34354
rect 30098 34302 30100 34354
rect 29820 34020 29876 34300
rect 30044 34290 30100 34302
rect 30156 34636 30324 34692
rect 30716 34916 30772 36540
rect 30940 35810 30996 35822
rect 30940 35758 30942 35810
rect 30994 35758 30996 35810
rect 30940 35028 30996 35758
rect 30940 34962 30996 34972
rect 29820 33954 29876 33964
rect 29484 33394 29540 33404
rect 28924 33282 28980 33292
rect 28700 33058 28756 33068
rect 29372 33124 29428 33134
rect 29484 33124 29540 33134
rect 29428 33122 29540 33124
rect 29428 33070 29486 33122
rect 29538 33070 29540 33122
rect 29428 33068 29540 33070
rect 28588 32452 28644 32462
rect 28476 32450 28644 32452
rect 28476 32398 28590 32450
rect 28642 32398 28644 32450
rect 28476 32396 28644 32398
rect 26796 31892 26852 31902
rect 26796 31798 26852 31836
rect 27244 31554 27300 31566
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 29988 25508 30830
rect 27244 30884 27300 31502
rect 28140 30996 28196 31006
rect 28588 30996 28644 32396
rect 28140 30994 28644 30996
rect 28140 30942 28142 30994
rect 28194 30942 28644 30994
rect 28140 30940 28644 30942
rect 27692 30884 27748 30894
rect 28140 30884 28196 30940
rect 27244 30882 28196 30884
rect 27244 30830 27694 30882
rect 27746 30830 28196 30882
rect 27244 30828 28196 30830
rect 27692 30818 27748 30828
rect 25788 30212 25844 30222
rect 25900 30212 25956 30222
rect 25788 30210 25900 30212
rect 25788 30158 25790 30210
rect 25842 30158 25900 30210
rect 25788 30156 25900 30158
rect 25788 30146 25844 30156
rect 25228 29538 25284 29550
rect 25228 29486 25230 29538
rect 25282 29486 25284 29538
rect 25228 29428 25284 29486
rect 25228 29362 25284 29372
rect 25452 29092 25508 29932
rect 25452 29026 25508 29036
rect 25564 29652 25620 29662
rect 25564 28868 25620 29596
rect 25564 28802 25620 28812
rect 25788 27858 25844 27870
rect 25788 27806 25790 27858
rect 25842 27806 25844 27858
rect 25788 27748 25844 27806
rect 25900 27748 25956 30156
rect 28140 30212 28196 30828
rect 28812 30884 28868 30894
rect 28812 30882 29204 30884
rect 28812 30830 28814 30882
rect 28866 30830 29204 30882
rect 28812 30828 29204 30830
rect 28812 30818 28868 30828
rect 26460 30098 26516 30110
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 26460 29316 26516 30046
rect 26460 29250 26516 29260
rect 26908 29652 26964 29662
rect 26908 29204 26964 29596
rect 27804 29652 27860 29662
rect 27804 29558 27860 29596
rect 27580 29538 27636 29550
rect 27580 29486 27582 29538
rect 27634 29486 27636 29538
rect 27580 29428 27636 29486
rect 27692 29540 27748 29550
rect 27692 29446 27748 29484
rect 27580 29362 27636 29372
rect 28028 29426 28084 29438
rect 28028 29374 28030 29426
rect 28082 29374 28084 29426
rect 27692 29316 27748 29326
rect 27692 29222 27748 29260
rect 26908 29138 26964 29148
rect 28028 28868 28084 29374
rect 28140 29316 28196 30156
rect 28588 30772 28644 30782
rect 28588 30322 28644 30716
rect 28588 30270 28590 30322
rect 28642 30270 28644 30322
rect 28588 29652 28644 30270
rect 29148 30322 29204 30828
rect 29148 30270 29150 30322
rect 29202 30270 29204 30322
rect 29148 30258 29204 30270
rect 29372 29988 29428 33068
rect 29484 33058 29540 33068
rect 29932 31108 29988 31118
rect 29820 31052 29932 31108
rect 29708 30884 29764 30894
rect 29596 30324 29652 30334
rect 29148 29932 29428 29988
rect 29484 30098 29540 30110
rect 29484 30046 29486 30098
rect 29538 30046 29540 30098
rect 28700 29652 28756 29662
rect 28588 29650 29092 29652
rect 28588 29598 28702 29650
rect 28754 29598 29092 29650
rect 28588 29596 29092 29598
rect 28700 29586 28756 29596
rect 28476 29540 28532 29550
rect 28476 29446 28532 29484
rect 28140 29250 28196 29260
rect 28812 29426 28868 29438
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28700 29204 28756 29214
rect 28476 28868 28532 28878
rect 28028 28812 28476 28868
rect 28140 28642 28196 28654
rect 28140 28590 28142 28642
rect 28194 28590 28196 28642
rect 28140 27858 28196 28590
rect 28364 28644 28420 28654
rect 28364 28530 28420 28588
rect 28364 28478 28366 28530
rect 28418 28478 28420 28530
rect 28364 28466 28420 28478
rect 28476 28082 28532 28812
rect 28476 28030 28478 28082
rect 28530 28030 28532 28082
rect 28476 28018 28532 28030
rect 28700 28084 28756 29148
rect 28812 28644 28868 29374
rect 29036 28866 29092 29596
rect 29036 28814 29038 28866
rect 29090 28814 29092 28866
rect 29036 28802 29092 28814
rect 28812 28578 28868 28588
rect 28700 28018 28756 28028
rect 28924 28084 28980 28094
rect 28924 27990 28980 28028
rect 28140 27806 28142 27858
rect 28194 27806 28196 27858
rect 26348 27748 26404 27758
rect 25900 27746 26404 27748
rect 25900 27694 26350 27746
rect 26402 27694 26404 27746
rect 25900 27692 26404 27694
rect 25788 27682 25844 27692
rect 26012 27074 26068 27086
rect 26012 27022 26014 27074
rect 26066 27022 26068 27074
rect 24668 26002 24724 26012
rect 25004 26852 25172 26908
rect 25788 26962 25844 26974
rect 25788 26910 25790 26962
rect 25842 26910 25844 26962
rect 25788 26908 25844 26910
rect 25340 26852 25396 26862
rect 24668 25732 24724 25742
rect 24612 25730 24724 25732
rect 24612 25678 24670 25730
rect 24722 25678 24724 25730
rect 24612 25676 24724 25678
rect 24556 25638 24612 25676
rect 24668 25666 24724 25676
rect 24556 25396 24612 25406
rect 24556 25302 24612 25340
rect 24892 23938 24948 23950
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24892 23604 24948 23886
rect 24892 23538 24948 23548
rect 24332 23266 24500 23268
rect 24332 23214 24334 23266
rect 24386 23214 24500 23266
rect 24332 23212 24500 23214
rect 24332 23202 24388 23212
rect 24108 23154 24164 23166
rect 24108 23102 24110 23154
rect 24162 23102 24164 23154
rect 24108 22260 24164 23102
rect 24220 23156 24276 23166
rect 24220 23062 24276 23100
rect 24444 22372 24500 22382
rect 24500 22316 24612 22372
rect 24444 22278 24500 22316
rect 24108 22194 24164 22204
rect 23996 21522 24052 21532
rect 24556 21474 24612 22316
rect 24556 21422 24558 21474
rect 24610 21422 24612 21474
rect 24556 21410 24612 21422
rect 24892 21588 24948 21598
rect 24892 20914 24948 21532
rect 24892 20862 24894 20914
rect 24946 20862 24948 20914
rect 24892 20850 24948 20862
rect 23212 19394 23268 19404
rect 23212 19236 23268 19246
rect 23212 18676 23268 19180
rect 23660 19236 23716 19246
rect 23660 19142 23716 19180
rect 24332 19236 24388 19246
rect 24332 19142 24388 19180
rect 25004 19236 25060 26852
rect 25340 26514 25396 26796
rect 25564 26850 25620 26862
rect 25564 26798 25566 26850
rect 25618 26798 25620 26850
rect 25564 26628 25620 26798
rect 25564 26562 25620 26572
rect 25676 26850 25732 26862
rect 25788 26852 25956 26908
rect 25676 26798 25678 26850
rect 25730 26798 25732 26850
rect 25340 26462 25342 26514
rect 25394 26462 25396 26514
rect 25340 26450 25396 26462
rect 25116 26404 25172 26414
rect 25116 26310 25172 26348
rect 25452 26404 25508 26414
rect 25676 26404 25732 26798
rect 25900 26740 25956 26852
rect 25900 26674 25956 26684
rect 25452 26402 25732 26404
rect 25452 26350 25454 26402
rect 25506 26350 25732 26402
rect 25452 26348 25732 26350
rect 26012 26404 26068 27022
rect 25452 26338 25508 26348
rect 26012 26338 26068 26348
rect 26236 27074 26292 27086
rect 26236 27022 26238 27074
rect 26290 27022 26292 27074
rect 26236 26292 26292 27022
rect 26348 26964 26404 27692
rect 26684 27300 26740 27310
rect 26684 27206 26740 27244
rect 28140 27300 28196 27806
rect 28140 27234 28196 27244
rect 26572 26962 26628 26974
rect 26572 26910 26574 26962
rect 26626 26910 26628 26962
rect 26572 26908 26628 26910
rect 29148 26908 29204 29932
rect 29484 29540 29540 30046
rect 29596 30098 29652 30268
rect 29596 30046 29598 30098
rect 29650 30046 29652 30098
rect 29596 30034 29652 30046
rect 29708 29986 29764 30828
rect 29708 29934 29710 29986
rect 29762 29934 29764 29986
rect 29708 29540 29764 29934
rect 29484 29474 29540 29484
rect 29596 29484 29764 29540
rect 29260 29316 29316 29326
rect 29596 29316 29652 29484
rect 29260 29314 29652 29316
rect 29260 29262 29262 29314
rect 29314 29262 29652 29314
rect 29260 29260 29652 29262
rect 29708 29316 29764 29326
rect 29260 29250 29316 29260
rect 29372 28866 29428 28878
rect 29372 28814 29374 28866
rect 29426 28814 29428 28866
rect 29372 28754 29428 28814
rect 29372 28702 29374 28754
rect 29426 28702 29428 28754
rect 29372 28690 29428 28702
rect 29708 28644 29764 29260
rect 29708 28578 29764 28588
rect 29820 28308 29876 31052
rect 29932 31042 29988 31052
rect 30156 30772 30212 34636
rect 30268 34244 30324 34254
rect 30268 34150 30324 34188
rect 30380 34130 30436 34142
rect 30380 34078 30382 34130
rect 30434 34078 30436 34130
rect 30380 33124 30436 34078
rect 30716 34130 30772 34860
rect 31052 34804 31108 36990
rect 31388 36484 31444 37324
rect 31500 37156 31556 37884
rect 31500 37090 31556 37100
rect 31500 36484 31556 36494
rect 31388 36482 31556 36484
rect 31388 36430 31502 36482
rect 31554 36430 31556 36482
rect 31388 36428 31556 36430
rect 31500 36418 31556 36428
rect 31164 36260 31220 36270
rect 31164 36166 31220 36204
rect 31500 35924 31556 35934
rect 31612 35924 31668 44268
rect 31948 44212 32004 44268
rect 31836 44156 32004 44212
rect 31836 43538 31892 44156
rect 31836 43486 31838 43538
rect 31890 43486 31892 43538
rect 31836 43474 31892 43486
rect 32060 43538 32116 44380
rect 32060 43486 32062 43538
rect 32114 43486 32116 43538
rect 32060 43474 32116 43486
rect 32172 41410 32228 48972
rect 32284 48468 32340 49196
rect 32732 49140 32788 49756
rect 32396 49138 32788 49140
rect 32396 49086 32734 49138
rect 32786 49086 32788 49138
rect 32396 49084 32788 49086
rect 32396 49026 32452 49084
rect 32732 49074 32788 49084
rect 32396 48974 32398 49026
rect 32450 48974 32452 49026
rect 32396 48962 32452 48974
rect 32508 48468 32564 48478
rect 32284 48466 32564 48468
rect 32284 48414 32510 48466
rect 32562 48414 32564 48466
rect 32284 48412 32564 48414
rect 32508 48402 32564 48412
rect 32508 46564 32564 46574
rect 32508 46470 32564 46508
rect 32844 46564 32900 57484
rect 32956 56308 33012 62412
rect 33068 60844 33348 60900
rect 33068 60564 33124 60844
rect 33292 60788 33348 60844
rect 33404 60788 33460 60798
rect 33292 60786 33460 60788
rect 33292 60734 33406 60786
rect 33458 60734 33460 60786
rect 33292 60732 33460 60734
rect 33404 60722 33460 60732
rect 33068 59890 33124 60508
rect 33180 60674 33236 60686
rect 33180 60622 33182 60674
rect 33234 60622 33236 60674
rect 33180 60340 33236 60622
rect 33180 60002 33236 60284
rect 33180 59950 33182 60002
rect 33234 59950 33236 60002
rect 33180 59938 33236 59950
rect 33068 59838 33070 59890
rect 33122 59838 33124 59890
rect 33068 59826 33124 59838
rect 33628 59780 33684 59790
rect 33628 59686 33684 59724
rect 33404 59108 33460 59118
rect 33180 57540 33236 57550
rect 33180 57446 33236 57484
rect 32956 56252 33124 56308
rect 32956 55300 33012 55310
rect 32956 55206 33012 55244
rect 32956 49252 33012 49262
rect 32956 49158 33012 49196
rect 32844 46498 32900 46508
rect 33068 46340 33124 56252
rect 33180 55410 33236 55422
rect 33180 55358 33182 55410
rect 33234 55358 33236 55410
rect 33180 54402 33236 55358
rect 33180 54350 33182 54402
rect 33234 54350 33236 54402
rect 33180 54292 33236 54350
rect 33180 54226 33236 54236
rect 33180 53506 33236 53518
rect 33180 53454 33182 53506
rect 33234 53454 33236 53506
rect 33180 52836 33236 53454
rect 33292 52836 33348 52846
rect 33180 52780 33292 52836
rect 33292 52388 33348 52780
rect 33404 52500 33460 59052
rect 33740 57540 33796 65436
rect 34860 65492 34916 65550
rect 34860 65426 34916 65436
rect 35532 65492 35588 65502
rect 35532 65398 35588 65436
rect 36652 65490 36708 65502
rect 36652 65438 36654 65490
rect 36706 65438 36708 65490
rect 34972 65380 35028 65390
rect 34972 65286 35028 65324
rect 35644 65380 35700 65390
rect 35084 65266 35140 65278
rect 35084 65214 35086 65266
rect 35138 65214 35140 65266
rect 34636 64484 34692 64494
rect 34636 63922 34692 64428
rect 35084 64036 35140 65214
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35644 64818 35700 65324
rect 35644 64766 35646 64818
rect 35698 64766 35700 64818
rect 35644 64754 35700 64766
rect 36428 64708 36484 64718
rect 36652 64708 36708 65438
rect 37436 65378 37492 65390
rect 37436 65326 37438 65378
rect 37490 65326 37492 65378
rect 37436 65268 37492 65326
rect 37436 65202 37492 65212
rect 38556 65380 38612 65390
rect 36428 64706 36652 64708
rect 36428 64654 36430 64706
rect 36482 64654 36652 64706
rect 36428 64652 36652 64654
rect 36428 64642 36484 64652
rect 36652 64642 36708 64652
rect 37100 64708 37156 64718
rect 37100 64614 37156 64652
rect 38556 64708 38612 65324
rect 38556 64614 38612 64652
rect 39228 64594 39284 64606
rect 39228 64542 39230 64594
rect 39282 64542 39284 64594
rect 39228 64148 39284 64542
rect 39228 64082 39284 64092
rect 35196 64036 35252 64046
rect 35084 64034 35252 64036
rect 35084 63982 35198 64034
rect 35250 63982 35252 64034
rect 35084 63980 35252 63982
rect 35196 63970 35252 63980
rect 34636 63870 34638 63922
rect 34690 63870 34692 63922
rect 34636 63858 34692 63870
rect 39340 63924 39396 66220
rect 39564 66274 39844 66276
rect 39564 66222 39790 66274
rect 39842 66222 39844 66274
rect 39564 66220 39844 66222
rect 39564 65378 39620 66220
rect 39788 66210 39844 66220
rect 41020 65492 41076 69200
rect 43036 67172 43092 69200
rect 43036 67116 43876 67172
rect 43820 66498 43876 67116
rect 43820 66446 43822 66498
rect 43874 66446 43876 66498
rect 43820 66434 43876 66446
rect 45052 66500 45108 69200
rect 47068 67228 47124 69200
rect 47068 67172 47572 67228
rect 45052 66434 45108 66444
rect 46172 66274 46228 66286
rect 46172 66222 46174 66274
rect 46226 66222 46228 66274
rect 43036 66164 43092 66174
rect 43036 66070 43092 66108
rect 46172 66164 46228 66222
rect 41020 65426 41076 65436
rect 42700 65492 42756 65502
rect 39564 65326 39566 65378
rect 39618 65326 39620 65378
rect 39564 65314 39620 65326
rect 40124 65378 40180 65390
rect 40124 65326 40126 65378
rect 40178 65326 40180 65378
rect 40124 65268 40180 65326
rect 41132 65380 41188 65390
rect 41132 65286 41188 65324
rect 41580 65380 41636 65390
rect 42028 65380 42084 65390
rect 41580 65378 41860 65380
rect 41580 65326 41582 65378
rect 41634 65326 41860 65378
rect 41580 65324 41860 65326
rect 41580 65314 41636 65324
rect 39452 63924 39508 63934
rect 39340 63922 39508 63924
rect 39340 63870 39454 63922
rect 39506 63870 39508 63922
rect 39340 63868 39508 63870
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 37884 62468 37940 62478
rect 37884 62374 37940 62412
rect 36316 62356 36372 62366
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35532 61684 35588 61694
rect 35532 61682 35812 61684
rect 35532 61630 35534 61682
rect 35586 61630 35812 61682
rect 35532 61628 35812 61630
rect 35532 61618 35588 61628
rect 34636 61458 34692 61470
rect 34636 61406 34638 61458
rect 34690 61406 34692 61458
rect 34636 61124 34692 61406
rect 35196 61458 35252 61470
rect 35196 61406 35198 61458
rect 35250 61406 35252 61458
rect 34748 61346 34804 61358
rect 34748 61294 34750 61346
rect 34802 61294 34804 61346
rect 34748 61236 34804 61294
rect 34972 61348 35028 61358
rect 34972 61346 35140 61348
rect 34972 61294 34974 61346
rect 35026 61294 35140 61346
rect 34972 61292 35140 61294
rect 34972 61282 35028 61292
rect 34748 61170 34804 61180
rect 34636 61058 34692 61068
rect 33852 60900 33908 60910
rect 34748 60900 34804 60910
rect 33908 60844 34020 60900
rect 33852 60834 33908 60844
rect 33964 60452 34020 60844
rect 34748 60786 34804 60844
rect 34748 60734 34750 60786
rect 34802 60734 34804 60786
rect 34748 60722 34804 60734
rect 34076 60676 34132 60686
rect 34524 60676 34580 60686
rect 34076 60674 34580 60676
rect 34076 60622 34078 60674
rect 34130 60622 34526 60674
rect 34578 60622 34580 60674
rect 34076 60620 34580 60622
rect 34076 60610 34132 60620
rect 33964 60396 34244 60452
rect 34188 60114 34244 60396
rect 34412 60226 34468 60620
rect 34524 60610 34580 60620
rect 34412 60174 34414 60226
rect 34466 60174 34468 60226
rect 34412 60162 34468 60174
rect 34748 60564 34804 60574
rect 34748 60226 34804 60508
rect 34748 60174 34750 60226
rect 34802 60174 34804 60226
rect 34748 60162 34804 60174
rect 35084 60228 35140 61292
rect 35196 61124 35252 61406
rect 35644 61460 35700 61470
rect 35420 61346 35476 61358
rect 35420 61294 35422 61346
rect 35474 61294 35476 61346
rect 35420 61236 35476 61294
rect 35420 61170 35476 61180
rect 35196 61058 35252 61068
rect 35420 60900 35476 60910
rect 35420 60806 35476 60844
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35084 60172 35476 60228
rect 34188 60062 34190 60114
rect 34242 60062 34244 60114
rect 34188 60050 34244 60062
rect 35420 59218 35476 60172
rect 35420 59166 35422 59218
rect 35474 59166 35476 59218
rect 35420 59154 35476 59166
rect 35644 58994 35700 61404
rect 35756 59220 35812 61628
rect 36316 61682 36372 62300
rect 37212 62354 37268 62366
rect 38780 62356 38836 62366
rect 37212 62302 37214 62354
rect 37266 62302 37268 62354
rect 36316 61630 36318 61682
rect 36370 61630 36372 61682
rect 36316 61618 36372 61630
rect 36764 62244 36820 62254
rect 36428 61458 36484 61470
rect 36428 61406 36430 61458
rect 36482 61406 36484 61458
rect 36204 61346 36260 61358
rect 36204 61294 36206 61346
rect 36258 61294 36260 61346
rect 36092 61236 36148 61246
rect 35868 61124 35924 61134
rect 35868 60786 35924 61068
rect 35868 60734 35870 60786
rect 35922 60734 35924 60786
rect 35868 60722 35924 60734
rect 36092 60786 36148 61180
rect 36092 60734 36094 60786
rect 36146 60734 36148 60786
rect 36092 60722 36148 60734
rect 36204 59332 36260 61294
rect 35980 59220 36036 59230
rect 35756 59218 36036 59220
rect 35756 59166 35982 59218
rect 36034 59166 36036 59218
rect 35756 59164 36036 59166
rect 35980 59154 36036 59164
rect 35644 58942 35646 58994
rect 35698 58942 35700 58994
rect 35644 58930 35700 58942
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 36204 58546 36260 59276
rect 36428 59108 36484 61406
rect 36764 60898 36820 62188
rect 36764 60846 36766 60898
rect 36818 60846 36820 60898
rect 36764 60834 36820 60846
rect 36988 61458 37044 61470
rect 36988 61406 36990 61458
rect 37042 61406 37044 61458
rect 36988 60564 37044 61406
rect 37212 61460 37268 62302
rect 38668 62354 38836 62356
rect 38668 62302 38782 62354
rect 38834 62302 38836 62354
rect 38668 62300 38836 62302
rect 37436 62244 37492 62254
rect 38556 62244 38612 62254
rect 37324 62242 37492 62244
rect 37324 62190 37438 62242
rect 37490 62190 37492 62242
rect 37324 62188 37492 62190
rect 37324 61460 37380 62188
rect 37436 62178 37492 62188
rect 38220 62242 38612 62244
rect 38220 62190 38558 62242
rect 38610 62190 38612 62242
rect 38220 62188 38612 62190
rect 37436 61684 37492 61694
rect 38220 61684 38276 62188
rect 38556 62178 38612 62188
rect 38668 62020 38724 62300
rect 38780 62290 38836 62300
rect 37436 61682 38276 61684
rect 37436 61630 37438 61682
rect 37490 61630 38222 61682
rect 38274 61630 38276 61682
rect 37436 61628 38276 61630
rect 37436 61618 37492 61628
rect 38220 61618 38276 61628
rect 38556 61964 38724 62020
rect 38556 61570 38612 61964
rect 38556 61518 38558 61570
rect 38610 61518 38612 61570
rect 37548 61460 37604 61470
rect 37324 61458 37604 61460
rect 37324 61406 37550 61458
rect 37602 61406 37604 61458
rect 37324 61404 37604 61406
rect 37212 61366 37268 61404
rect 37548 60900 37604 61404
rect 38332 61346 38388 61358
rect 38332 61294 38334 61346
rect 38386 61294 38388 61346
rect 38332 61012 38388 61294
rect 38332 60946 38388 60956
rect 37548 60834 37604 60844
rect 37772 60788 37828 60798
rect 37772 60694 37828 60732
rect 36988 60498 37044 60508
rect 37324 60676 37380 60686
rect 37212 59332 37268 59342
rect 37212 59238 37268 59276
rect 36876 59108 36932 59118
rect 36428 59106 36932 59108
rect 36428 59054 36878 59106
rect 36930 59054 36932 59106
rect 36428 59052 36932 59054
rect 36876 58772 36932 59052
rect 37324 58996 37380 60620
rect 37996 60676 38052 60686
rect 37996 60582 38052 60620
rect 38556 60674 38612 61518
rect 39116 60900 39172 60938
rect 39116 60834 39172 60844
rect 39004 60786 39060 60798
rect 39004 60734 39006 60786
rect 39058 60734 39060 60786
rect 38556 60622 38558 60674
rect 38610 60622 38612 60674
rect 38556 60610 38612 60622
rect 38668 60676 38724 60686
rect 38668 60114 38724 60620
rect 39004 60676 39060 60734
rect 39004 60610 39060 60620
rect 38668 60062 38670 60114
rect 38722 60062 38724 60114
rect 38668 60050 38724 60062
rect 37324 58930 37380 58940
rect 38108 59780 38164 59790
rect 36876 58716 37044 58772
rect 36204 58494 36206 58546
rect 36258 58494 36260 58546
rect 36204 58482 36260 58494
rect 35980 58322 36036 58334
rect 35980 58270 35982 58322
rect 36034 58270 36036 58322
rect 35980 57764 36036 58270
rect 33740 57474 33796 57484
rect 35868 57708 35980 57764
rect 34972 57428 35028 57438
rect 33740 56980 33796 56990
rect 34972 56980 35028 57372
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 33740 56886 33796 56924
rect 34524 56978 35028 56980
rect 34524 56926 34974 56978
rect 35026 56926 35028 56978
rect 34524 56924 35028 56926
rect 34524 56866 34580 56924
rect 34972 56914 35028 56924
rect 34524 56814 34526 56866
rect 34578 56814 34580 56866
rect 34524 56802 34580 56814
rect 35196 56756 35252 56766
rect 35196 56194 35252 56700
rect 35196 56142 35198 56194
rect 35250 56142 35252 56194
rect 35196 56130 35252 56142
rect 35644 56196 35700 56206
rect 35644 56102 35700 56140
rect 33628 56084 33684 56094
rect 33628 56082 33796 56084
rect 33628 56030 33630 56082
rect 33682 56030 33796 56082
rect 33628 56028 33796 56030
rect 33628 56018 33684 56028
rect 33740 55412 33796 56028
rect 33740 54404 33796 55356
rect 34188 56082 34244 56094
rect 34188 56030 34190 56082
rect 34242 56030 34244 56082
rect 33852 55300 33908 55310
rect 34188 55300 34244 56030
rect 35868 56082 35924 57708
rect 35980 57698 36036 57708
rect 36204 58210 36260 58222
rect 36204 58158 36206 58210
rect 36258 58158 36260 58210
rect 36204 57538 36260 58158
rect 36428 57764 36484 57774
rect 36204 57486 36206 57538
rect 36258 57486 36260 57538
rect 35868 56030 35870 56082
rect 35922 56030 35924 56082
rect 35868 56018 35924 56030
rect 35980 56866 36036 56878
rect 35980 56814 35982 56866
rect 36034 56814 36036 56866
rect 35980 56084 36036 56814
rect 36092 56756 36148 56766
rect 36092 56662 36148 56700
rect 36204 56196 36260 57486
rect 36316 57762 36484 57764
rect 36316 57710 36430 57762
rect 36482 57710 36484 57762
rect 36316 57708 36484 57710
rect 36316 56978 36372 57708
rect 36428 57698 36484 57708
rect 36316 56926 36318 56978
rect 36370 56926 36372 56978
rect 36316 56914 36372 56926
rect 36428 56868 36484 56878
rect 36428 56756 36484 56812
rect 36204 56130 36260 56140
rect 36316 56754 36484 56756
rect 36316 56702 36430 56754
rect 36482 56702 36484 56754
rect 36316 56700 36484 56702
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 55524 35252 55534
rect 35196 55430 35252 55468
rect 35980 55524 36036 56028
rect 35980 55458 36036 55468
rect 36316 55972 36372 56700
rect 36428 56690 36484 56700
rect 36988 56532 37044 58716
rect 37772 58548 37828 58558
rect 37660 57764 37716 57774
rect 37660 57650 37716 57708
rect 37660 57598 37662 57650
rect 37714 57598 37716 57650
rect 37660 57586 37716 57598
rect 37772 57428 37828 58492
rect 37772 57204 37828 57372
rect 37660 57148 37828 57204
rect 37100 56868 37156 56878
rect 37100 56774 37156 56812
rect 37324 56866 37380 56878
rect 37324 56814 37326 56866
rect 37378 56814 37380 56866
rect 37324 56756 37380 56814
rect 37324 56690 37380 56700
rect 36988 56476 37380 56532
rect 37324 56194 37380 56476
rect 37324 56142 37326 56194
rect 37378 56142 37380 56194
rect 37324 56130 37380 56142
rect 37212 56084 37268 56094
rect 37212 55990 37268 56028
rect 34860 55412 34916 55422
rect 34860 55318 34916 55356
rect 34748 55300 34804 55310
rect 33852 55298 34804 55300
rect 33852 55246 33854 55298
rect 33906 55246 34750 55298
rect 34802 55246 34804 55298
rect 33852 55244 34804 55246
rect 33852 55234 33908 55244
rect 34748 55234 34804 55244
rect 33628 54348 33796 54404
rect 33516 52836 33572 52846
rect 33516 52742 33572 52780
rect 33404 52444 33572 52500
rect 33292 52162 33348 52332
rect 33292 52110 33294 52162
rect 33346 52110 33348 52162
rect 33292 52098 33348 52110
rect 33404 52164 33460 52174
rect 33404 50818 33460 52108
rect 33404 50766 33406 50818
rect 33458 50766 33460 50818
rect 33404 50754 33460 50766
rect 33292 50594 33348 50606
rect 33292 50542 33294 50594
rect 33346 50542 33348 50594
rect 33180 49698 33236 49710
rect 33180 49646 33182 49698
rect 33234 49646 33236 49698
rect 33180 49252 33236 49646
rect 33180 49186 33236 49196
rect 33292 49250 33348 50542
rect 33404 49812 33460 49822
rect 33404 49718 33460 49756
rect 33292 49198 33294 49250
rect 33346 49198 33348 49250
rect 33292 49186 33348 49198
rect 33068 46284 33460 46340
rect 33180 45780 33236 45790
rect 33180 45686 33236 45724
rect 32508 45106 32564 45118
rect 32508 45054 32510 45106
rect 32562 45054 32564 45106
rect 32396 44996 32452 45006
rect 32284 44436 32340 44446
rect 32284 44342 32340 44380
rect 32396 44324 32452 44940
rect 32396 44230 32452 44268
rect 32396 43764 32452 43774
rect 32508 43764 32564 45054
rect 33292 44996 33348 45006
rect 33292 44902 33348 44940
rect 33068 44324 33124 44334
rect 33068 44230 33124 44268
rect 32396 43762 32564 43764
rect 32396 43710 32398 43762
rect 32450 43710 32564 43762
rect 32396 43708 32564 43710
rect 32396 43698 32452 43708
rect 33180 43092 33236 43102
rect 33180 42978 33236 43036
rect 33180 42926 33182 42978
rect 33234 42926 33236 42978
rect 33180 42866 33236 42926
rect 33180 42814 33182 42866
rect 33234 42814 33236 42866
rect 33180 42802 33236 42814
rect 33404 41972 33460 46284
rect 33292 41916 33460 41972
rect 32508 41858 32564 41870
rect 32508 41806 32510 41858
rect 32562 41806 32564 41858
rect 32508 41524 32564 41806
rect 32508 41458 32564 41468
rect 32172 41358 32174 41410
rect 32226 41358 32228 41410
rect 32172 41346 32228 41358
rect 32508 41298 32564 41310
rect 32508 41246 32510 41298
rect 32562 41246 32564 41298
rect 32060 41186 32116 41198
rect 32060 41134 32062 41186
rect 32114 41134 32116 41186
rect 32060 39396 32116 41134
rect 32508 41188 32564 41246
rect 32172 39732 32228 39742
rect 32508 39732 32564 41132
rect 33180 41186 33236 41198
rect 33180 41134 33182 41186
rect 33234 41134 33236 41186
rect 33180 41076 33236 41134
rect 33180 41010 33236 41020
rect 32172 39638 32228 39676
rect 32284 39730 32564 39732
rect 32284 39678 32510 39730
rect 32562 39678 32564 39730
rect 32284 39676 32564 39678
rect 32060 39330 32116 39340
rect 31836 38780 32228 38836
rect 31836 37938 31892 38780
rect 32172 38724 32228 38780
rect 32284 38724 32340 39676
rect 32508 39666 32564 39676
rect 33068 39396 33124 39406
rect 32956 39394 33124 39396
rect 32956 39342 33070 39394
rect 33122 39342 33124 39394
rect 32956 39340 33124 39342
rect 32172 38722 32340 38724
rect 32172 38670 32174 38722
rect 32226 38670 32340 38722
rect 32172 38668 32340 38670
rect 32508 38834 32564 38846
rect 32508 38782 32510 38834
rect 32562 38782 32564 38834
rect 32172 38658 32228 38668
rect 31836 37886 31838 37938
rect 31890 37886 31892 37938
rect 31836 37874 31892 37886
rect 31948 38610 32004 38622
rect 31948 38558 31950 38610
rect 32002 38558 32004 38610
rect 31948 38500 32004 38558
rect 31500 35922 31668 35924
rect 31500 35870 31502 35922
rect 31554 35870 31668 35922
rect 31500 35868 31668 35870
rect 31500 35858 31556 35868
rect 31052 34738 31108 34748
rect 31388 35698 31444 35710
rect 31388 35646 31390 35698
rect 31442 35646 31444 35698
rect 30716 34078 30718 34130
rect 30770 34078 30772 34130
rect 30716 34066 30772 34078
rect 30940 34244 30996 34254
rect 30380 33068 30548 33124
rect 30492 31780 30548 33068
rect 30492 31714 30548 31724
rect 30940 33122 30996 34188
rect 31388 34242 31444 35646
rect 31388 34190 31390 34242
rect 31442 34190 31444 34242
rect 31388 34178 31444 34190
rect 31612 35028 31668 35038
rect 31612 34018 31668 34972
rect 31836 34132 31892 34142
rect 31836 34038 31892 34076
rect 31612 33966 31614 34018
rect 31666 33966 31668 34018
rect 31612 33954 31668 33966
rect 31836 33684 31892 33694
rect 31500 33460 31556 33470
rect 31276 33348 31332 33358
rect 31276 33254 31332 33292
rect 30940 33070 30942 33122
rect 30994 33070 30996 33122
rect 30940 31556 30996 33070
rect 31500 33122 31556 33404
rect 31500 33070 31502 33122
rect 31554 33070 31556 33122
rect 31500 33058 31556 33070
rect 31612 33348 31668 33358
rect 31052 32452 31108 32462
rect 31500 32452 31556 32462
rect 31052 32450 31556 32452
rect 31052 32398 31054 32450
rect 31106 32398 31502 32450
rect 31554 32398 31556 32450
rect 31052 32396 31556 32398
rect 31052 32386 31108 32396
rect 31500 31892 31556 32396
rect 31500 31826 31556 31836
rect 31612 31892 31668 33292
rect 31836 33346 31892 33628
rect 31836 33294 31838 33346
rect 31890 33294 31892 33346
rect 31836 33282 31892 33294
rect 31836 32676 31892 32686
rect 31724 32562 31780 32574
rect 31724 32510 31726 32562
rect 31778 32510 31780 32562
rect 31724 32452 31780 32510
rect 31836 32562 31892 32620
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 31724 32386 31780 32396
rect 31836 31892 31892 31902
rect 31612 31890 31892 31892
rect 31612 31838 31838 31890
rect 31890 31838 31892 31890
rect 31612 31836 31892 31838
rect 30156 30706 30212 30716
rect 30380 31500 30996 31556
rect 30156 30324 30212 30334
rect 30156 30210 30212 30268
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 30156 30146 30212 30158
rect 30380 30098 30436 31500
rect 31052 31220 31108 31230
rect 31052 31126 31108 31164
rect 31612 30882 31668 31836
rect 31836 31826 31892 31836
rect 31948 31556 32004 38444
rect 32508 38052 32564 38782
rect 32956 38668 33012 39340
rect 33068 39330 33124 39340
rect 33292 38668 33348 41916
rect 33404 41746 33460 41758
rect 33404 41694 33406 41746
rect 33458 41694 33460 41746
rect 33404 41524 33460 41694
rect 33404 41458 33460 41468
rect 33516 41410 33572 52444
rect 33628 52274 33684 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36316 53954 36372 55916
rect 37660 55298 37716 57148
rect 37996 56868 38052 56878
rect 37996 56774 38052 56812
rect 37660 55246 37662 55298
rect 37714 55246 37716 55298
rect 37660 55234 37716 55246
rect 36316 53902 36318 53954
rect 36370 53902 36372 53954
rect 36316 53890 36372 53902
rect 36092 53842 36148 53854
rect 36092 53790 36094 53842
rect 36146 53790 36148 53842
rect 34524 53732 34580 53742
rect 34524 53638 34580 53676
rect 35980 53730 36036 53742
rect 35980 53678 35982 53730
rect 36034 53678 36036 53730
rect 35980 53172 36036 53678
rect 35980 53106 36036 53116
rect 35644 53060 35700 53070
rect 33628 52222 33630 52274
rect 33682 52222 33684 52274
rect 33628 52210 33684 52222
rect 33740 52946 33796 52958
rect 33740 52894 33742 52946
rect 33794 52894 33796 52946
rect 33740 52276 33796 52894
rect 34412 52948 34468 52958
rect 34412 52854 34468 52892
rect 35644 52946 35700 53004
rect 35644 52894 35646 52946
rect 35698 52894 35700 52946
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 33740 52050 33796 52220
rect 35644 52164 35700 52894
rect 35980 52948 36036 52958
rect 35980 52274 36036 52892
rect 36092 52386 36148 53790
rect 36204 53844 36260 53854
rect 36204 53058 36260 53788
rect 37100 53844 37156 53854
rect 37100 53750 37156 53788
rect 37996 53844 38052 53854
rect 36428 53732 36484 53742
rect 36204 53006 36206 53058
rect 36258 53006 36260 53058
rect 36204 52994 36260 53006
rect 36316 53172 36372 53182
rect 36092 52334 36094 52386
rect 36146 52334 36148 52386
rect 36092 52322 36148 52334
rect 35980 52222 35982 52274
rect 36034 52222 36036 52274
rect 35980 52210 36036 52222
rect 35644 52070 35700 52108
rect 33740 51998 33742 52050
rect 33794 51998 33796 52050
rect 33740 51986 33796 51998
rect 36316 51602 36372 53116
rect 36428 53170 36484 53676
rect 36428 53118 36430 53170
rect 36482 53118 36484 53170
rect 36428 53106 36484 53118
rect 37324 53730 37380 53742
rect 37324 53678 37326 53730
rect 37378 53678 37380 53730
rect 37324 53172 37380 53678
rect 37996 53730 38052 53788
rect 37996 53678 37998 53730
rect 38050 53678 38052 53730
rect 37996 53666 38052 53678
rect 37324 53106 37380 53116
rect 36652 53060 36708 53070
rect 36652 52966 36708 53004
rect 36764 52948 36820 52958
rect 36764 52854 36820 52892
rect 36316 51550 36318 51602
rect 36370 51550 36372 51602
rect 36316 51538 36372 51550
rect 37324 51492 37380 51502
rect 37324 51490 37940 51492
rect 37324 51438 37326 51490
rect 37378 51438 37940 51490
rect 37324 51436 37940 51438
rect 36204 51380 36260 51390
rect 35532 51378 36260 51380
rect 35532 51326 36206 51378
rect 36258 51326 36260 51378
rect 35532 51324 36260 51326
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50706 35252 50718
rect 35196 50654 35198 50706
rect 35250 50654 35252 50706
rect 35084 50594 35140 50606
rect 35084 50542 35086 50594
rect 35138 50542 35140 50594
rect 35084 50428 35140 50542
rect 34860 50372 35140 50428
rect 34076 49922 34132 49934
rect 34076 49870 34078 49922
rect 34130 49870 34132 49922
rect 34076 49812 34132 49870
rect 34188 49812 34244 49822
rect 34076 49756 34188 49812
rect 34188 49746 34244 49756
rect 34860 49698 34916 50372
rect 35084 49812 35140 49822
rect 35196 49812 35252 50654
rect 35420 50036 35476 50046
rect 35532 50036 35588 51324
rect 36204 51314 36260 51324
rect 36764 51378 36820 51390
rect 36764 51326 36766 51378
rect 36818 51326 36820 51378
rect 36764 51268 36820 51326
rect 36316 50708 36372 50718
rect 36764 50708 36820 51212
rect 36316 50706 36820 50708
rect 36316 50654 36318 50706
rect 36370 50654 36820 50706
rect 36316 50652 36820 50654
rect 36316 50642 36372 50652
rect 37324 50428 37380 51436
rect 37884 51380 37940 51436
rect 37996 51380 38052 51390
rect 37884 51378 38052 51380
rect 37884 51326 37998 51378
rect 38050 51326 38052 51378
rect 37884 51324 38052 51326
rect 37996 51314 38052 51324
rect 37772 51268 37828 51278
rect 37772 51174 37828 51212
rect 35420 50034 35588 50036
rect 35420 49982 35422 50034
rect 35474 49982 35588 50034
rect 35420 49980 35588 49982
rect 37212 50372 37380 50428
rect 38108 50428 38164 59724
rect 39228 59108 39284 59118
rect 39004 58996 39060 59006
rect 38556 58548 38612 58558
rect 38556 58434 38612 58492
rect 38556 58382 38558 58434
rect 38610 58382 38612 58434
rect 38556 58370 38612 58382
rect 39004 57762 39060 58940
rect 39228 58546 39284 59052
rect 39228 58494 39230 58546
rect 39282 58494 39284 58546
rect 39228 58482 39284 58494
rect 39004 57710 39006 57762
rect 39058 57710 39060 57762
rect 39004 57698 39060 57710
rect 38220 56756 38276 56766
rect 38220 56082 38276 56700
rect 38220 56030 38222 56082
rect 38274 56030 38276 56082
rect 38220 56018 38276 56030
rect 39004 56084 39060 56094
rect 39004 55990 39060 56028
rect 38332 55188 38388 55198
rect 38332 55094 38388 55132
rect 38556 53508 38612 53518
rect 38444 53452 38556 53508
rect 38444 50428 38500 53452
rect 38556 53442 38612 53452
rect 38892 52164 38948 52174
rect 38668 52162 38948 52164
rect 38668 52110 38894 52162
rect 38946 52110 38948 52162
rect 38668 52108 38948 52110
rect 38668 51490 38724 52108
rect 38892 52098 38948 52108
rect 38668 51438 38670 51490
rect 38722 51438 38724 51490
rect 38668 51426 38724 51438
rect 38556 51268 38612 51278
rect 38612 51212 38724 51268
rect 38556 51202 38612 51212
rect 38556 50706 38612 50718
rect 38556 50654 38558 50706
rect 38610 50654 38612 50706
rect 38556 50428 38612 50654
rect 38108 50372 38276 50428
rect 38444 50372 38612 50428
rect 35420 49970 35476 49980
rect 35140 49756 35252 49812
rect 35084 49718 35140 49756
rect 34860 49646 34862 49698
rect 34914 49646 34916 49698
rect 34860 49476 34916 49646
rect 37212 49698 37268 50372
rect 37660 49924 37716 49934
rect 37660 49830 37716 49868
rect 37212 49646 37214 49698
rect 37266 49646 37268 49698
rect 34860 49410 34916 49420
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 33740 49252 33796 49262
rect 33740 49138 33796 49196
rect 33740 49086 33742 49138
rect 33794 49086 33796 49138
rect 33740 49074 33796 49086
rect 35084 48804 35140 48814
rect 34636 47570 34692 47582
rect 34636 47518 34638 47570
rect 34690 47518 34692 47570
rect 34636 47460 34692 47518
rect 34636 47394 34692 47404
rect 34748 47458 34804 47470
rect 34748 47406 34750 47458
rect 34802 47406 34804 47458
rect 34748 46900 34804 47406
rect 34748 46786 34804 46844
rect 34748 46734 34750 46786
rect 34802 46734 34804 46786
rect 34748 46722 34804 46734
rect 34972 47460 35028 47470
rect 34972 46674 35028 47404
rect 34972 46622 34974 46674
rect 35026 46622 35028 46674
rect 34972 46610 35028 46622
rect 33964 45890 34020 45902
rect 33964 45838 33966 45890
rect 34018 45838 34020 45890
rect 33964 45668 34020 45838
rect 34412 45668 34468 45678
rect 33964 45666 34468 45668
rect 33964 45614 34414 45666
rect 34466 45614 34468 45666
rect 33964 45612 34468 45614
rect 34412 45332 34468 45612
rect 34412 45266 34468 45276
rect 34076 45220 34132 45230
rect 33964 44996 34020 45006
rect 33740 44324 33796 44334
rect 33740 44230 33796 44268
rect 33964 44098 34020 44940
rect 34076 44212 34132 45164
rect 34300 44324 34356 44334
rect 34748 44324 34804 44334
rect 34300 44322 34804 44324
rect 34300 44270 34302 44322
rect 34354 44270 34750 44322
rect 34802 44270 34804 44322
rect 34300 44268 34804 44270
rect 35084 44324 35140 48748
rect 37212 48354 37268 49646
rect 37212 48302 37214 48354
rect 37266 48302 37268 48354
rect 37212 48290 37268 48302
rect 35980 48244 36036 48254
rect 35532 48242 36036 48244
rect 35532 48190 35982 48242
rect 36034 48190 36036 48242
rect 35532 48188 36036 48190
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35420 47684 35476 47694
rect 35420 47590 35476 47628
rect 35532 47236 35588 48188
rect 35980 48178 36036 48188
rect 37100 48242 37156 48254
rect 37100 48190 37102 48242
rect 37154 48190 37156 48242
rect 36652 48130 36708 48142
rect 36652 48078 36654 48130
rect 36706 48078 36708 48130
rect 36652 47684 36708 48078
rect 36652 47618 36708 47628
rect 35308 47180 35588 47236
rect 36428 47460 36484 47470
rect 35308 46898 35364 47180
rect 35308 46846 35310 46898
rect 35362 46846 35364 46898
rect 35308 46834 35364 46846
rect 36092 47124 36148 47134
rect 36092 46898 36148 47068
rect 36092 46846 36094 46898
rect 36146 46846 36148 46898
rect 36092 46834 36148 46846
rect 36428 46898 36484 47404
rect 37100 47236 37156 48190
rect 37436 47684 37492 47694
rect 37436 47570 37492 47628
rect 37436 47518 37438 47570
rect 37490 47518 37492 47570
rect 37436 47506 37492 47518
rect 37996 47572 38052 47582
rect 37996 47478 38052 47516
rect 37100 47170 37156 47180
rect 37660 47458 37716 47470
rect 37660 47406 37662 47458
rect 37714 47406 37716 47458
rect 37660 47236 37716 47406
rect 37660 47170 37716 47180
rect 36428 46846 36430 46898
rect 36482 46846 36484 46898
rect 36428 46834 36484 46846
rect 35868 46786 35924 46798
rect 35868 46734 35870 46786
rect 35922 46734 35924 46786
rect 35756 46674 35812 46686
rect 35756 46622 35758 46674
rect 35810 46622 35812 46674
rect 35756 46452 35812 46622
rect 35868 46676 35924 46734
rect 37436 46786 37492 46798
rect 37436 46734 37438 46786
rect 37490 46734 37492 46786
rect 35868 46610 35924 46620
rect 36652 46676 36708 46686
rect 36652 46582 36708 46620
rect 37436 46676 37492 46734
rect 37100 46562 37156 46574
rect 37100 46510 37102 46562
rect 37154 46510 37156 46562
rect 35756 46386 35812 46396
rect 36316 46452 36372 46462
rect 36316 46358 36372 46396
rect 37100 46452 37156 46510
rect 37100 46386 37156 46396
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 36204 45332 36260 45342
rect 36204 45106 36260 45276
rect 36652 45332 36708 45342
rect 36652 45238 36708 45276
rect 36204 45054 36206 45106
rect 36258 45054 36260 45106
rect 36204 45042 36260 45054
rect 35420 44996 35476 45006
rect 35420 44902 35476 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35308 44324 35364 44334
rect 35084 44322 35364 44324
rect 35084 44270 35310 44322
rect 35362 44270 35364 44322
rect 35084 44268 35364 44270
rect 34300 44258 34356 44268
rect 34748 44258 34804 44268
rect 34076 44118 34132 44156
rect 33964 44046 33966 44098
rect 34018 44046 34020 44098
rect 33964 44034 34020 44046
rect 34636 44100 34692 44110
rect 34636 44006 34692 44044
rect 34860 44100 34916 44110
rect 35308 44100 35364 44268
rect 35644 44100 35700 44110
rect 35308 44098 35700 44100
rect 35308 44046 35646 44098
rect 35698 44046 35700 44098
rect 35308 44044 35700 44046
rect 34860 44006 34916 44044
rect 35644 43876 35700 44044
rect 35644 43810 35700 43820
rect 36764 43988 36820 43998
rect 36652 43650 36708 43662
rect 36652 43598 36654 43650
rect 36706 43598 36708 43650
rect 33740 43540 33796 43550
rect 33796 43484 33908 43540
rect 33740 43474 33796 43484
rect 33628 42530 33684 42542
rect 33628 42478 33630 42530
rect 33682 42478 33684 42530
rect 33628 41524 33684 42478
rect 33740 42084 33796 42094
rect 33740 41970 33796 42028
rect 33740 41918 33742 41970
rect 33794 41918 33796 41970
rect 33740 41906 33796 41918
rect 33740 41748 33796 41758
rect 33740 41654 33796 41692
rect 33628 41458 33684 41468
rect 33516 41358 33518 41410
rect 33570 41358 33572 41410
rect 33516 41346 33572 41358
rect 33516 41188 33572 41198
rect 33516 41094 33572 41132
rect 33852 38668 33908 43484
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34076 42978 34132 42990
rect 34076 42926 34078 42978
rect 34130 42926 34132 42978
rect 34076 42866 34132 42926
rect 34076 42814 34078 42866
rect 34130 42814 34132 42866
rect 34076 42084 34132 42814
rect 36428 42530 36484 42542
rect 36428 42478 36430 42530
rect 36482 42478 36484 42530
rect 36428 42196 36484 42478
rect 36428 42130 36484 42140
rect 34076 41990 34132 42028
rect 35532 42084 35588 42094
rect 35532 41990 35588 42028
rect 35868 41972 35924 41982
rect 36652 41972 36708 43598
rect 35868 41970 36708 41972
rect 35868 41918 35870 41970
rect 35922 41918 36708 41970
rect 35868 41916 36708 41918
rect 34412 41858 34468 41870
rect 34412 41806 34414 41858
rect 34466 41806 34468 41858
rect 34412 41524 34468 41806
rect 34636 41748 34692 41758
rect 34636 41746 34916 41748
rect 34636 41694 34638 41746
rect 34690 41694 34916 41746
rect 34636 41692 34916 41694
rect 34636 41682 34692 41692
rect 34412 41458 34468 41468
rect 34860 41298 34916 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34860 41246 34862 41298
rect 34914 41246 34916 41298
rect 34860 41234 34916 41246
rect 32956 38612 33124 38668
rect 32956 38052 33012 38062
rect 32508 38050 33012 38052
rect 32508 37998 32958 38050
rect 33010 37998 33012 38050
rect 32508 37996 33012 37998
rect 32060 36370 32116 36382
rect 32060 36318 32062 36370
rect 32114 36318 32116 36370
rect 32060 36260 32116 36318
rect 32060 32786 32116 36204
rect 32956 36258 33012 37996
rect 32956 36206 32958 36258
rect 33010 36206 33012 36258
rect 32956 36194 33012 36206
rect 33068 37044 33124 38612
rect 32396 35812 32452 35822
rect 32284 35810 32452 35812
rect 32284 35758 32398 35810
rect 32450 35758 32452 35810
rect 32284 35756 32452 35758
rect 32060 32734 32062 32786
rect 32114 32734 32116 32786
rect 32060 32722 32116 32734
rect 32172 35588 32228 35598
rect 32060 31780 32116 31790
rect 32060 31686 32116 31724
rect 32060 31556 32116 31566
rect 31948 31554 32116 31556
rect 31948 31502 32062 31554
rect 32114 31502 32116 31554
rect 31948 31500 32116 31502
rect 32060 31490 32116 31500
rect 32060 31220 32116 31230
rect 32172 31220 32228 35532
rect 32284 32676 32340 35756
rect 32396 35746 32452 35756
rect 32508 35700 32564 35710
rect 32508 35606 32564 35644
rect 32396 35474 32452 35486
rect 32396 35422 32398 35474
rect 32450 35422 32452 35474
rect 32396 33234 32452 35422
rect 32956 33684 33012 33694
rect 33068 33684 33124 36988
rect 33012 33628 33124 33684
rect 33180 38612 33348 38668
rect 33740 38612 33908 38668
rect 33964 41186 34020 41198
rect 33964 41134 33966 41186
rect 34018 41134 34020 41186
rect 32956 33618 33012 33628
rect 32396 33182 32398 33234
rect 32450 33182 32452 33234
rect 32396 33170 32452 33182
rect 32284 32116 32340 32620
rect 32284 32050 32340 32060
rect 33068 31892 33124 31902
rect 33068 31666 33124 31836
rect 33068 31614 33070 31666
rect 33122 31614 33124 31666
rect 33068 31602 33124 31614
rect 32116 31164 32228 31220
rect 32060 31126 32116 31164
rect 31612 30830 31614 30882
rect 31666 30830 31668 30882
rect 31612 30818 31668 30830
rect 32284 30212 32340 30222
rect 30380 30046 30382 30098
rect 30434 30046 30436 30098
rect 30380 30034 30436 30046
rect 30492 30100 30548 30110
rect 29932 29988 29988 29998
rect 29932 29894 29988 29932
rect 30380 28756 30436 28766
rect 30492 28756 30548 30044
rect 31276 30100 31332 30110
rect 31276 30006 31332 30044
rect 30604 29988 30660 29998
rect 30604 29426 30660 29932
rect 31388 29988 31444 29998
rect 31612 29988 31668 29998
rect 31388 29894 31444 29932
rect 31500 29986 31668 29988
rect 31500 29934 31614 29986
rect 31666 29934 31668 29986
rect 31500 29932 31668 29934
rect 31500 29764 31556 29932
rect 31612 29922 31668 29932
rect 31052 29708 31556 29764
rect 30828 29652 30884 29662
rect 30828 29558 30884 29596
rect 30604 29374 30606 29426
rect 30658 29374 30660 29426
rect 30604 28868 30660 29374
rect 31052 29426 31108 29708
rect 31836 29652 31892 29662
rect 31836 29558 31892 29596
rect 31164 29540 31220 29550
rect 31164 29446 31220 29484
rect 31052 29374 31054 29426
rect 31106 29374 31108 29426
rect 31052 29362 31108 29374
rect 31388 29316 31444 29326
rect 31388 29314 31780 29316
rect 31388 29262 31390 29314
rect 31442 29262 31780 29314
rect 31388 29260 31780 29262
rect 31388 29250 31444 29260
rect 31276 29092 31332 29102
rect 31332 29036 31444 29092
rect 31276 29026 31332 29036
rect 30660 28812 30884 28868
rect 30604 28774 30660 28812
rect 30436 28700 30548 28756
rect 30380 28690 30436 28700
rect 30268 28644 30324 28654
rect 30492 28644 30548 28700
rect 30604 28644 30660 28654
rect 30492 28642 30660 28644
rect 30492 28590 30606 28642
rect 30658 28590 30660 28642
rect 30492 28588 30660 28590
rect 30268 28550 30324 28588
rect 30604 28578 30660 28588
rect 30716 28532 30772 28542
rect 30716 28438 30772 28476
rect 29484 28252 29876 28308
rect 26348 26898 26404 26908
rect 26460 26852 26628 26908
rect 26684 26852 26740 26862
rect 26460 26514 26516 26852
rect 26684 26758 26740 26796
rect 27020 26852 27076 26862
rect 26460 26462 26462 26514
rect 26514 26462 26516 26514
rect 26460 26450 26516 26462
rect 27020 26516 27076 26796
rect 28588 26850 28644 26862
rect 28588 26798 28590 26850
rect 28642 26798 28644 26850
rect 27356 26516 27412 26526
rect 27020 26514 27412 26516
rect 27020 26462 27358 26514
rect 27410 26462 27412 26514
rect 27020 26460 27412 26462
rect 26348 26292 26404 26302
rect 26572 26292 26628 26302
rect 26236 26290 26404 26292
rect 26236 26238 26350 26290
rect 26402 26238 26404 26290
rect 26236 26236 26404 26238
rect 26124 26178 26180 26190
rect 26124 26126 26126 26178
rect 26178 26126 26180 26178
rect 25900 26068 25956 26078
rect 25788 26066 25956 26068
rect 25788 26014 25902 26066
rect 25954 26014 25956 26066
rect 25788 26012 25956 26014
rect 25564 25508 25620 25518
rect 25788 25508 25844 26012
rect 25900 26002 25956 26012
rect 26124 25956 26180 26126
rect 26124 25890 26180 25900
rect 26236 26068 26292 26078
rect 25452 25506 25844 25508
rect 25452 25454 25566 25506
rect 25618 25454 25844 25506
rect 25452 25452 25844 25454
rect 25900 25732 25956 25742
rect 25900 25506 25956 25676
rect 25900 25454 25902 25506
rect 25954 25454 25956 25506
rect 25452 25060 25508 25452
rect 25564 25442 25620 25452
rect 25900 25060 25956 25454
rect 26012 25620 26068 25630
rect 26012 25506 26068 25564
rect 26124 25620 26180 25630
rect 26236 25620 26292 26012
rect 26348 25956 26404 26236
rect 26348 25890 26404 25900
rect 26460 26236 26572 26292
rect 26124 25618 26292 25620
rect 26124 25566 26126 25618
rect 26178 25566 26292 25618
rect 26124 25564 26292 25566
rect 26460 25620 26516 26236
rect 26572 26198 26628 26236
rect 26124 25554 26180 25564
rect 26460 25554 26516 25564
rect 26908 26180 26964 26190
rect 26908 25732 26964 26124
rect 26012 25454 26014 25506
rect 26066 25454 26068 25506
rect 26012 25442 26068 25454
rect 26908 25506 26964 25676
rect 26908 25454 26910 25506
rect 26962 25454 26964 25506
rect 26908 25442 26964 25454
rect 26684 25394 26740 25406
rect 26684 25342 26686 25394
rect 26738 25342 26740 25394
rect 26236 25284 26292 25294
rect 26236 25190 26292 25228
rect 25340 24834 25396 24846
rect 25340 24782 25342 24834
rect 25394 24782 25396 24834
rect 25228 24724 25284 24734
rect 25116 23716 25172 23726
rect 25116 22260 25172 23660
rect 25228 23266 25284 24668
rect 25340 23828 25396 24782
rect 25340 23762 25396 23772
rect 25340 23492 25396 23502
rect 25340 23378 25396 23436
rect 25340 23326 25342 23378
rect 25394 23326 25396 23378
rect 25340 23314 25396 23326
rect 25228 23214 25230 23266
rect 25282 23214 25284 23266
rect 25228 23202 25284 23214
rect 25228 22260 25284 22270
rect 25116 22204 25228 22260
rect 25228 22194 25284 22204
rect 25340 22260 25396 22270
rect 25452 22260 25508 25004
rect 25676 25004 25956 25060
rect 26684 25060 26740 25342
rect 25564 24948 25620 24958
rect 25564 24854 25620 24892
rect 25564 23380 25620 23390
rect 25676 23380 25732 25004
rect 26684 24994 26740 25004
rect 26348 24948 26404 24958
rect 26404 24892 26516 24948
rect 26348 24882 26404 24892
rect 26348 24500 26404 24510
rect 26348 23826 26404 24444
rect 26348 23774 26350 23826
rect 26402 23774 26404 23826
rect 25564 23378 25732 23380
rect 25564 23326 25566 23378
rect 25618 23326 25732 23378
rect 25564 23324 25732 23326
rect 25788 23492 25844 23502
rect 25788 23378 25844 23436
rect 25788 23326 25790 23378
rect 25842 23326 25844 23378
rect 25564 23314 25620 23324
rect 25788 23314 25844 23326
rect 25900 23154 25956 23166
rect 25900 23102 25902 23154
rect 25954 23102 25956 23154
rect 25900 22372 25956 23102
rect 25900 22306 25956 22316
rect 25340 22258 25508 22260
rect 25340 22206 25342 22258
rect 25394 22206 25508 22258
rect 25340 22204 25508 22206
rect 25340 22194 25396 22204
rect 25340 21812 25396 21822
rect 25340 21718 25396 21756
rect 26348 21698 26404 23774
rect 26460 23940 26516 24892
rect 27020 24500 27076 26460
rect 27356 26450 27412 26460
rect 28476 26516 28532 26526
rect 28588 26516 28644 26798
rect 28476 26514 28588 26516
rect 28476 26462 28478 26514
rect 28530 26462 28588 26514
rect 28476 26460 28588 26462
rect 28476 26450 28532 26460
rect 28588 26450 28644 26460
rect 28924 26852 29204 26908
rect 29372 26962 29428 26974
rect 29372 26910 29374 26962
rect 29426 26910 29428 26962
rect 29372 26908 29428 26910
rect 29484 26908 29540 28252
rect 29372 26852 29540 26908
rect 29708 28084 29764 28094
rect 27468 26404 27524 26414
rect 27132 26290 27188 26302
rect 27132 26238 27134 26290
rect 27186 26238 27188 26290
rect 27132 25620 27188 26238
rect 27468 26290 27524 26348
rect 28812 26404 28868 26414
rect 28812 26310 28868 26348
rect 27468 26238 27470 26290
rect 27522 26238 27524 26290
rect 27468 26226 27524 26238
rect 28252 26292 28308 26302
rect 28252 26198 28308 26236
rect 28588 26292 28644 26302
rect 27132 25554 27188 25564
rect 27244 26178 27300 26190
rect 27244 26126 27246 26178
rect 27298 26126 27300 26178
rect 27244 25508 27300 26126
rect 27804 26068 27860 26078
rect 27804 26066 27972 26068
rect 27804 26014 27806 26066
rect 27858 26014 27972 26066
rect 27804 26012 27972 26014
rect 27804 26002 27860 26012
rect 27580 25844 27636 25854
rect 27580 25508 27636 25788
rect 27692 25732 27748 25742
rect 27692 25638 27748 25676
rect 27804 25620 27860 25630
rect 27804 25526 27860 25564
rect 27692 25508 27748 25518
rect 27580 25452 27692 25508
rect 27244 25442 27300 25452
rect 27356 25396 27412 25406
rect 27356 25394 27636 25396
rect 27356 25342 27358 25394
rect 27410 25342 27636 25394
rect 27356 25340 27636 25342
rect 27356 25330 27412 25340
rect 27580 24836 27636 25340
rect 27692 25060 27748 25452
rect 27916 25396 27972 26012
rect 28140 25620 28196 25630
rect 28028 25396 28084 25406
rect 27916 25340 28028 25396
rect 28028 25330 28084 25340
rect 27692 25004 27972 25060
rect 27692 24836 27748 24846
rect 27580 24780 27692 24836
rect 27748 24780 27860 24836
rect 27692 24742 27748 24780
rect 27468 24724 27524 24734
rect 27524 24668 27636 24724
rect 27468 24630 27524 24668
rect 27132 24500 27188 24510
rect 27020 24444 27132 24500
rect 27132 24406 27188 24444
rect 27580 24052 27636 24668
rect 27692 24052 27748 24062
rect 27580 24050 27748 24052
rect 27580 23998 27694 24050
rect 27746 23998 27748 24050
rect 27580 23996 27748 23998
rect 27692 23986 27748 23996
rect 26908 23940 26964 23950
rect 26460 23938 26964 23940
rect 26460 23886 26910 23938
rect 26962 23886 26964 23938
rect 26460 23884 26964 23886
rect 26460 22372 26516 23884
rect 26908 23874 26964 23884
rect 26796 23714 26852 23726
rect 26796 23662 26798 23714
rect 26850 23662 26852 23714
rect 26796 23492 26852 23662
rect 26796 23426 26852 23436
rect 26908 23604 26964 23614
rect 26460 22370 26852 22372
rect 26460 22318 26462 22370
rect 26514 22318 26852 22370
rect 26460 22316 26852 22318
rect 26460 22306 26516 22316
rect 26348 21646 26350 21698
rect 26402 21646 26404 21698
rect 26348 21634 26404 21646
rect 26796 21586 26852 22316
rect 26796 21534 26798 21586
rect 26850 21534 26852 21586
rect 26796 21522 26852 21534
rect 26908 22370 26964 23548
rect 27580 23380 27636 23390
rect 27580 23286 27636 23324
rect 27804 23044 27860 24780
rect 27916 23938 27972 25004
rect 28140 24946 28196 25564
rect 28588 25620 28644 26236
rect 28924 26180 28980 26852
rect 29036 26516 29092 26526
rect 29036 26514 29316 26516
rect 29036 26462 29038 26514
rect 29090 26462 29316 26514
rect 29036 26460 29316 26462
rect 29036 26450 29092 26460
rect 29148 26292 29204 26302
rect 29148 26198 29204 26236
rect 28588 25526 28644 25564
rect 28812 26124 28980 26180
rect 28140 24894 28142 24946
rect 28194 24894 28196 24946
rect 28140 24724 28196 24894
rect 28700 24724 28756 24734
rect 28140 24658 28196 24668
rect 28252 24722 28756 24724
rect 28252 24670 28702 24722
rect 28754 24670 28756 24722
rect 28252 24668 28756 24670
rect 27916 23886 27918 23938
rect 27970 23886 27972 23938
rect 27916 23874 27972 23886
rect 28252 23940 28308 24668
rect 28700 24658 28756 24668
rect 28252 23826 28308 23884
rect 28252 23774 28254 23826
rect 28306 23774 28308 23826
rect 28252 23762 28308 23774
rect 27916 23492 27972 23502
rect 27972 23436 28084 23492
rect 27916 23426 27972 23436
rect 27916 23044 27972 23054
rect 27804 23042 27972 23044
rect 27804 22990 27918 23042
rect 27970 22990 27972 23042
rect 27804 22988 27972 22990
rect 27916 22978 27972 22988
rect 26908 22318 26910 22370
rect 26962 22318 26964 22370
rect 26908 21588 26964 22318
rect 27804 22260 27860 22270
rect 27916 22260 27972 22270
rect 27860 22258 27972 22260
rect 27860 22206 27918 22258
rect 27970 22206 27972 22258
rect 27860 22204 27972 22206
rect 27804 21698 27860 22204
rect 27916 22194 27972 22204
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 27804 21634 27860 21646
rect 27244 21588 27300 21598
rect 26908 21586 27300 21588
rect 26908 21534 27246 21586
rect 27298 21534 27300 21586
rect 26908 21532 27300 21534
rect 27244 21522 27300 21532
rect 28028 20804 28084 23436
rect 28812 23156 28868 26124
rect 29260 26068 29316 26460
rect 29372 26292 29428 26852
rect 29596 26516 29652 26526
rect 29596 26402 29652 26460
rect 29596 26350 29598 26402
rect 29650 26350 29652 26402
rect 29596 26338 29652 26350
rect 29372 26226 29428 26236
rect 29708 26180 29764 28028
rect 30828 28082 30884 28812
rect 31052 28812 31332 28868
rect 30940 28644 30996 28654
rect 31052 28644 31108 28812
rect 30940 28642 31108 28644
rect 30940 28590 30942 28642
rect 30994 28590 31108 28642
rect 30940 28588 31108 28590
rect 31164 28644 31220 28654
rect 30940 28578 30996 28588
rect 31164 28196 31220 28588
rect 30828 28030 30830 28082
rect 30882 28030 30884 28082
rect 30828 28018 30884 28030
rect 30940 28140 31220 28196
rect 30604 27076 30660 27086
rect 30940 27076 30996 28140
rect 30604 27074 30996 27076
rect 30604 27022 30606 27074
rect 30658 27022 30942 27074
rect 30994 27022 30996 27074
rect 30604 27020 30996 27022
rect 30604 27010 30660 27020
rect 30940 27010 30996 27020
rect 31052 27972 31108 27982
rect 29820 26852 29876 26862
rect 29820 26850 29988 26852
rect 29820 26798 29822 26850
rect 29874 26798 29988 26850
rect 29820 26796 29988 26798
rect 29820 26786 29876 26796
rect 29932 26516 29988 26796
rect 30268 26516 30324 26526
rect 29932 26460 30268 26516
rect 30268 26422 30324 26460
rect 30828 26516 30884 26526
rect 30828 26422 30884 26460
rect 29596 26124 29764 26180
rect 30156 26290 30212 26302
rect 30156 26238 30158 26290
rect 30210 26238 30212 26290
rect 29484 26068 29540 26078
rect 29260 26066 29540 26068
rect 29260 26014 29486 26066
rect 29538 26014 29540 26066
rect 29260 26012 29540 26014
rect 28924 25620 28980 25630
rect 28924 25284 28980 25564
rect 29148 25508 29204 25518
rect 29148 25414 29204 25452
rect 29484 25394 29540 26012
rect 29484 25342 29486 25394
rect 29538 25342 29540 25394
rect 29484 25330 29540 25342
rect 28924 25218 28980 25228
rect 29484 25172 29540 25182
rect 28924 24836 28980 24846
rect 28924 24742 28980 24780
rect 29148 24722 29204 24734
rect 29148 24670 29150 24722
rect 29202 24670 29204 24722
rect 29036 24610 29092 24622
rect 29036 24558 29038 24610
rect 29090 24558 29092 24610
rect 29036 24052 29092 24558
rect 29148 24612 29204 24670
rect 29484 24722 29540 25116
rect 29484 24670 29486 24722
rect 29538 24670 29540 24722
rect 29484 24658 29540 24670
rect 29148 24546 29204 24556
rect 29148 24052 29204 24062
rect 29036 24050 29204 24052
rect 29036 23998 29150 24050
rect 29202 23998 29204 24050
rect 29036 23996 29204 23998
rect 29148 23986 29204 23996
rect 29260 23716 29316 23726
rect 29260 23622 29316 23660
rect 28812 23090 28868 23100
rect 28476 22146 28532 22158
rect 28476 22094 28478 22146
rect 28530 22094 28532 22146
rect 28476 21812 28532 22094
rect 28476 21746 28532 21756
rect 29372 20916 29428 20926
rect 27356 20802 28084 20804
rect 27356 20750 28030 20802
rect 28082 20750 28084 20802
rect 27356 20748 28084 20750
rect 27356 20188 27412 20748
rect 28028 20738 28084 20748
rect 29036 20802 29092 20814
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 26796 20132 26852 20142
rect 26684 20076 26796 20132
rect 26572 20020 26628 20030
rect 26572 19926 26628 19964
rect 26236 19348 26292 19358
rect 26236 19254 26292 19292
rect 25004 19170 25060 19180
rect 26572 19236 26628 19246
rect 26684 19236 26740 20076
rect 26796 20038 26852 20076
rect 27244 20132 27412 20188
rect 28252 20578 28308 20590
rect 28252 20526 28254 20578
rect 28306 20526 28308 20578
rect 27244 20020 27300 20132
rect 27244 19926 27300 19964
rect 27468 20130 27524 20142
rect 27468 20078 27470 20130
rect 27522 20078 27524 20130
rect 26572 19234 26740 19236
rect 26572 19182 26574 19234
rect 26626 19182 26740 19234
rect 26572 19180 26740 19182
rect 26796 19348 26852 19358
rect 26796 19234 26852 19292
rect 26796 19182 26798 19234
rect 26850 19182 26852 19234
rect 26572 19170 26628 19180
rect 26796 19170 26852 19182
rect 27132 19122 27188 19134
rect 27132 19070 27134 19122
rect 27186 19070 27188 19122
rect 22988 18620 23268 18676
rect 22988 18450 23044 18620
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 22988 18386 23044 18398
rect 23100 18452 23156 18462
rect 22876 18172 23044 18228
rect 22764 17462 22820 17500
rect 22988 17444 23044 18172
rect 23100 17666 23156 18396
rect 23212 18450 23268 18620
rect 23996 19010 24052 19022
rect 23996 18958 23998 19010
rect 24050 18958 24052 19010
rect 23996 18564 24052 18958
rect 26684 19010 26740 19022
rect 26684 18958 26686 19010
rect 26738 18958 26740 19010
rect 26684 18676 26740 18958
rect 26012 18620 26740 18676
rect 24220 18564 24276 18574
rect 23996 18508 24220 18564
rect 23212 18398 23214 18450
rect 23266 18398 23268 18450
rect 23212 18386 23268 18398
rect 24220 18450 24276 18508
rect 24220 18398 24222 18450
rect 24274 18398 24276 18450
rect 24220 18386 24276 18398
rect 24444 18562 24500 18574
rect 24444 18510 24446 18562
rect 24498 18510 24500 18562
rect 23772 18340 23828 18350
rect 23772 18246 23828 18284
rect 24444 18340 24500 18510
rect 26012 18562 26068 18620
rect 26012 18510 26014 18562
rect 26066 18510 26068 18562
rect 26012 18498 26068 18510
rect 23100 17614 23102 17666
rect 23154 17614 23156 17666
rect 23100 17602 23156 17614
rect 24444 17668 24500 18284
rect 25340 18450 25396 18462
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 24444 17602 24500 17612
rect 25004 18116 25060 18126
rect 22988 17388 23156 17444
rect 22652 17164 23044 17220
rect 22204 16828 22820 16884
rect 20412 16146 20468 16156
rect 21868 16212 21924 16222
rect 19292 15988 19348 15998
rect 19068 15932 19292 15988
rect 19292 15894 19348 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 21868 15538 21924 16156
rect 22428 16212 22484 16222
rect 22428 16118 22484 16156
rect 21868 15486 21870 15538
rect 21922 15486 21924 15538
rect 21868 15474 21924 15486
rect 22428 15202 22484 15214
rect 22428 15150 22430 15202
rect 22482 15150 22484 15202
rect 18732 15092 19348 15148
rect 19068 14532 19124 14542
rect 18844 14308 18900 14318
rect 18844 14306 19012 14308
rect 18844 14254 18846 14306
rect 18898 14254 19012 14306
rect 18844 14252 19012 14254
rect 18844 14242 18900 14252
rect 18732 13860 18788 13870
rect 18732 13766 18788 13804
rect 18844 13748 18900 13758
rect 18844 13654 18900 13692
rect 18956 13746 19012 14252
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13524 19012 13694
rect 18956 13458 19012 13468
rect 19068 13188 19124 14476
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18620 12898 18676 12910
rect 18844 13132 19124 13188
rect 18732 12852 18788 12862
rect 18732 12758 18788 12796
rect 18844 12852 18900 13132
rect 19180 12852 19236 12862
rect 18844 12850 19012 12852
rect 18844 12798 18846 12850
rect 18898 12798 19012 12850
rect 18844 12796 19012 12798
rect 18844 12786 18900 12796
rect 18844 12066 18900 12078
rect 18844 12014 18846 12066
rect 18898 12014 18900 12066
rect 18732 11508 18788 11518
rect 18732 11282 18788 11452
rect 18844 11396 18900 12014
rect 18956 11732 19012 12796
rect 19180 12758 19236 12796
rect 18956 11666 19012 11676
rect 18844 11330 18900 11340
rect 18732 11230 18734 11282
rect 18786 11230 18788 11282
rect 18732 10948 18788 11230
rect 18956 11284 19012 11294
rect 18956 11190 19012 11228
rect 18844 11172 18900 11182
rect 18844 11078 18900 11116
rect 19180 11170 19236 11182
rect 19180 11118 19182 11170
rect 19234 11118 19236 11170
rect 18732 10892 19012 10948
rect 18508 10780 18788 10836
rect 18396 10724 18452 10734
rect 18396 10630 18452 10668
rect 18732 10722 18788 10780
rect 18732 10670 18734 10722
rect 18786 10670 18788 10722
rect 18732 10658 18788 10670
rect 18956 10386 19012 10892
rect 19180 10612 19236 11118
rect 19292 10836 19348 15092
rect 22204 15090 22260 15102
rect 22204 15038 22206 15090
rect 22258 15038 22260 15090
rect 22204 14532 22260 15038
rect 22428 14868 22484 15150
rect 22652 15148 22708 16828
rect 22764 16770 22820 16828
rect 22764 16718 22766 16770
rect 22818 16718 22820 16770
rect 22764 16706 22820 16718
rect 22764 16212 22820 16222
rect 22764 16098 22820 16156
rect 22764 16046 22766 16098
rect 22818 16046 22820 16098
rect 22764 16034 22820 16046
rect 22988 16098 23044 17164
rect 22988 16046 22990 16098
rect 23042 16046 23044 16098
rect 22988 16034 23044 16046
rect 22988 15876 23044 15886
rect 22988 15782 23044 15820
rect 22652 15092 22820 15148
rect 22652 14868 22708 14878
rect 22428 14812 22652 14868
rect 22652 14642 22708 14812
rect 22652 14590 22654 14642
rect 22706 14590 22708 14642
rect 22652 14578 22708 14590
rect 22428 14532 22484 14542
rect 22204 14476 22428 14532
rect 22092 14306 22148 14318
rect 22092 14254 22094 14306
rect 22146 14254 22148 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20748 13972 20804 13982
rect 20748 13878 20804 13916
rect 21308 13916 21588 13972
rect 19852 13860 19908 13870
rect 19852 13746 19908 13804
rect 21084 13860 21140 13870
rect 20188 13748 20244 13758
rect 20860 13748 20916 13758
rect 19852 13694 19854 13746
rect 19906 13694 19908 13746
rect 19404 13634 19460 13646
rect 19404 13582 19406 13634
rect 19458 13582 19460 13634
rect 19404 13524 19460 13582
rect 19404 13458 19460 13468
rect 19852 13412 19908 13694
rect 19852 13346 19908 13356
rect 20076 13746 20244 13748
rect 20076 13694 20190 13746
rect 20242 13694 20244 13746
rect 20076 13692 20244 13694
rect 19964 13188 20020 13198
rect 19628 13186 20020 13188
rect 19628 13134 19966 13186
rect 20018 13134 20020 13186
rect 19628 13132 20020 13134
rect 19516 13074 19572 13086
rect 19516 13022 19518 13074
rect 19570 13022 19572 13074
rect 19404 12740 19460 12750
rect 19404 12646 19460 12684
rect 19516 11618 19572 13022
rect 19516 11566 19518 11618
rect 19570 11566 19572 11618
rect 19516 11554 19572 11566
rect 19628 11618 19684 13132
rect 19964 13122 20020 13132
rect 20076 13188 20132 13692
rect 20188 13682 20244 13692
rect 20524 13746 20916 13748
rect 20524 13694 20862 13746
rect 20914 13694 20916 13746
rect 20524 13692 20916 13694
rect 20412 13524 20468 13534
rect 20412 13430 20468 13468
rect 19852 12964 19908 12974
rect 20076 12964 20132 13132
rect 20300 13412 20356 13422
rect 19852 12962 20132 12964
rect 19852 12910 19854 12962
rect 19906 12910 20132 12962
rect 19852 12908 20132 12910
rect 20188 13076 20244 13086
rect 20300 13076 20356 13356
rect 20524 13186 20580 13692
rect 20860 13682 20916 13692
rect 21084 13746 21140 13804
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13682 21140 13694
rect 21308 13746 21364 13916
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21308 13682 21364 13694
rect 21420 13746 21476 13758
rect 21420 13694 21422 13746
rect 21474 13694 21476 13746
rect 20524 13134 20526 13186
rect 20578 13134 20580 13186
rect 20524 13122 20580 13134
rect 21196 13524 21252 13534
rect 21196 13188 21252 13468
rect 21308 13188 21364 13198
rect 21196 13186 21364 13188
rect 21196 13134 21310 13186
rect 21362 13134 21364 13186
rect 21196 13132 21364 13134
rect 21308 13122 21364 13132
rect 20412 13076 20468 13086
rect 20300 13074 20468 13076
rect 20300 13022 20414 13074
rect 20466 13022 20468 13074
rect 20300 13020 20468 13022
rect 19852 12898 19908 12908
rect 19964 12740 20020 12750
rect 20188 12740 20244 13020
rect 20412 13010 20468 13020
rect 20860 13076 20916 13086
rect 19964 12738 20244 12740
rect 19964 12686 19966 12738
rect 20018 12686 20244 12738
rect 19964 12684 20244 12686
rect 19964 12674 20020 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20860 12402 20916 13020
rect 21420 13074 21476 13694
rect 21532 13524 21588 13916
rect 22092 13860 22148 14254
rect 21756 13748 21812 13758
rect 21756 13654 21812 13692
rect 21980 13524 22036 13534
rect 21532 13522 22036 13524
rect 21532 13470 21982 13522
rect 22034 13470 22036 13522
rect 21532 13468 22036 13470
rect 21420 13022 21422 13074
rect 21474 13022 21476 13074
rect 21420 13010 21476 13022
rect 21644 12962 21700 12974
rect 21644 12910 21646 12962
rect 21698 12910 21700 12962
rect 21644 12852 21700 12910
rect 21644 12786 21700 12796
rect 20860 12350 20862 12402
rect 20914 12350 20916 12402
rect 20860 12338 20916 12350
rect 21196 12066 21252 12078
rect 21196 12014 21198 12066
rect 21250 12014 21252 12066
rect 21196 11956 21252 12014
rect 21196 11890 21252 11900
rect 19628 11566 19630 11618
rect 19682 11566 19684 11618
rect 19628 11554 19684 11566
rect 21308 11732 21364 11742
rect 21308 11282 21364 11676
rect 21308 11230 21310 11282
rect 21362 11230 21364 11282
rect 21308 11218 21364 11230
rect 21532 11394 21588 11406
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 20188 11172 20244 11182
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19292 10770 19348 10780
rect 20188 10612 20244 11116
rect 19180 10546 19236 10556
rect 19964 10556 20244 10612
rect 21532 10724 21588 11342
rect 21980 11284 22036 13468
rect 22092 13188 22148 13804
rect 22204 13748 22260 13758
rect 22204 13634 22260 13692
rect 22428 13746 22484 14476
rect 22652 13860 22708 13870
rect 22652 13766 22708 13804
rect 22428 13694 22430 13746
rect 22482 13694 22484 13746
rect 22428 13682 22484 13694
rect 22764 13746 22820 15092
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22764 13682 22820 13694
rect 22988 13746 23044 13758
rect 22988 13694 22990 13746
rect 23042 13694 23044 13746
rect 22204 13582 22206 13634
rect 22258 13582 22260 13634
rect 22204 13522 22260 13582
rect 22204 13470 22206 13522
rect 22258 13470 22260 13522
rect 22204 13458 22260 13470
rect 22988 13300 23044 13694
rect 23100 13748 23156 17388
rect 23324 15988 23380 15998
rect 24444 15988 24500 15998
rect 23212 15986 23380 15988
rect 23212 15934 23326 15986
rect 23378 15934 23380 15986
rect 23212 15932 23380 15934
rect 23212 14644 23268 15932
rect 23324 15922 23380 15932
rect 24220 15986 24500 15988
rect 24220 15934 24446 15986
rect 24498 15934 24500 15986
rect 24220 15932 24500 15934
rect 23660 15876 23716 15886
rect 23660 15202 23716 15820
rect 24220 15426 24276 15932
rect 24444 15922 24500 15932
rect 24220 15374 24222 15426
rect 24274 15374 24276 15426
rect 24220 15362 24276 15374
rect 24556 15874 24612 15886
rect 24556 15822 24558 15874
rect 24610 15822 24612 15874
rect 23660 15150 23662 15202
rect 23714 15150 23716 15202
rect 23660 15138 23716 15150
rect 23772 15314 23828 15326
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 23212 14578 23268 14588
rect 23548 14530 23604 14542
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23100 13682 23156 13692
rect 23212 14308 23268 14318
rect 23548 14308 23604 14478
rect 23212 14306 23604 14308
rect 23212 14254 23214 14306
rect 23266 14254 23604 14306
rect 23212 14252 23604 14254
rect 23212 13636 23268 14252
rect 23212 13570 23268 13580
rect 23324 13860 23380 13870
rect 23324 13746 23380 13804
rect 23324 13694 23326 13746
rect 23378 13694 23380 13746
rect 22764 13244 23044 13300
rect 22092 13132 22708 13188
rect 22540 12964 22596 12974
rect 22540 12870 22596 12908
rect 22092 12852 22148 12862
rect 22428 12852 22484 12862
rect 22092 12850 22428 12852
rect 22092 12798 22094 12850
rect 22146 12798 22428 12850
rect 22092 12796 22428 12798
rect 22092 12786 22148 12796
rect 22428 12758 22484 12796
rect 22652 11732 22708 13132
rect 22652 11666 22708 11676
rect 22764 12850 22820 13244
rect 23324 12962 23380 13694
rect 23660 13746 23716 13758
rect 23660 13694 23662 13746
rect 23714 13694 23716 13746
rect 23548 13524 23604 13534
rect 23660 13524 23716 13694
rect 23772 13636 23828 15262
rect 24556 15148 24612 15822
rect 24668 15874 24724 15886
rect 24668 15822 24670 15874
rect 24722 15822 24724 15874
rect 24668 15764 24724 15822
rect 24780 15764 24836 15774
rect 24668 15708 24780 15764
rect 24780 15698 24836 15708
rect 24332 15092 24612 15148
rect 24332 14642 24388 15092
rect 24332 14590 24334 14642
rect 24386 14590 24388 14642
rect 24332 14578 24388 14590
rect 24332 14308 24388 14318
rect 23884 13972 23940 13982
rect 24332 13972 24388 14252
rect 23884 13970 24388 13972
rect 23884 13918 23886 13970
rect 23938 13918 24334 13970
rect 24386 13918 24388 13970
rect 23884 13916 24388 13918
rect 23884 13906 23940 13916
rect 24332 13906 24388 13916
rect 23772 13634 24500 13636
rect 23772 13582 23774 13634
rect 23826 13582 24500 13634
rect 23772 13580 24500 13582
rect 23772 13570 23828 13580
rect 23604 13468 23716 13524
rect 23548 13186 23604 13468
rect 23548 13134 23550 13186
rect 23602 13134 23604 13186
rect 23548 13122 23604 13134
rect 23772 13188 23828 13198
rect 23772 13094 23828 13132
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 24220 12964 24276 12974
rect 24220 12870 24276 12908
rect 24444 12962 24500 13580
rect 24668 13524 24724 13534
rect 24444 12910 24446 12962
rect 24498 12910 24500 12962
rect 24444 12898 24500 12910
rect 24556 13188 24612 13198
rect 22764 12798 22766 12850
rect 22818 12798 22820 12850
rect 21980 11218 22036 11228
rect 19180 10388 19236 10398
rect 18956 10334 18958 10386
rect 19010 10334 19012 10386
rect 18956 10322 19012 10334
rect 19068 10386 19236 10388
rect 19068 10334 19182 10386
rect 19234 10334 19236 10386
rect 19068 10332 19236 10334
rect 18844 10052 18900 10062
rect 17948 10050 18564 10052
rect 17948 9998 17950 10050
rect 18002 9998 18564 10050
rect 17948 9996 18564 9998
rect 17948 9986 18004 9996
rect 18172 9826 18228 9838
rect 18172 9774 18174 9826
rect 18226 9774 18228 9826
rect 17948 9716 18004 9726
rect 17836 9660 17948 9716
rect 17948 9650 18004 9660
rect 17500 9214 17502 9266
rect 17554 9214 17556 9266
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 15484 6692 15540 6702
rect 15484 6598 15540 6636
rect 17500 6692 17556 9214
rect 18172 9156 18228 9774
rect 18508 9268 18564 9996
rect 18620 9940 18676 9950
rect 18620 9846 18676 9884
rect 18844 9826 18900 9996
rect 19068 9828 19124 10332
rect 19180 10322 19236 10332
rect 19404 10386 19460 10398
rect 19404 10334 19406 10386
rect 19458 10334 19460 10386
rect 19404 10052 19460 10334
rect 19852 10386 19908 10398
rect 19852 10334 19854 10386
rect 19906 10334 19908 10386
rect 19404 9996 19684 10052
rect 18844 9774 18846 9826
rect 18898 9774 18900 9826
rect 18844 9762 18900 9774
rect 18956 9772 19124 9828
rect 19404 9828 19460 9838
rect 18620 9716 18676 9726
rect 18620 9622 18676 9660
rect 18956 9716 19012 9772
rect 19404 9734 19460 9772
rect 19516 9826 19572 9838
rect 19516 9774 19518 9826
rect 19570 9774 19572 9826
rect 18956 9650 19012 9660
rect 19068 9604 19124 9642
rect 19068 9538 19124 9548
rect 19068 9380 19124 9390
rect 18844 9324 19068 9380
rect 18732 9268 18788 9278
rect 18508 9266 18788 9268
rect 18508 9214 18734 9266
rect 18786 9214 18788 9266
rect 18508 9212 18788 9214
rect 18732 9202 18788 9212
rect 18844 9266 18900 9324
rect 19068 9314 19124 9324
rect 19516 9380 19572 9774
rect 19516 9314 19572 9324
rect 18844 9214 18846 9266
rect 18898 9214 18900 9266
rect 18844 9202 18900 9214
rect 18172 9090 18228 9100
rect 18956 9156 19012 9166
rect 18956 9062 19012 9100
rect 19404 9156 19460 9166
rect 19460 9100 19572 9156
rect 19404 9090 19460 9100
rect 19292 9042 19348 9054
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 18844 7924 18900 7934
rect 18732 7868 18844 7924
rect 18732 7586 18788 7868
rect 18844 7858 18900 7868
rect 19292 7812 19348 8990
rect 19292 7756 19460 7812
rect 19068 7700 19124 7710
rect 18732 7534 18734 7586
rect 18786 7534 18788 7586
rect 18732 7028 18788 7534
rect 18284 6972 18788 7028
rect 17724 6804 17780 6814
rect 17500 6626 17556 6636
rect 17612 6748 17724 6804
rect 16156 6580 16212 6590
rect 16156 6486 16212 6524
rect 17388 6580 17444 6590
rect 17388 6130 17444 6524
rect 17388 6078 17390 6130
rect 17442 6078 17444 6130
rect 17388 6066 17444 6078
rect 17500 6020 17556 6030
rect 17612 6020 17668 6748
rect 17724 6738 17780 6748
rect 18284 6802 18340 6972
rect 18284 6750 18286 6802
rect 18338 6750 18340 6802
rect 18284 6738 18340 6750
rect 18620 6804 18676 6814
rect 18620 6710 18676 6748
rect 17500 6018 17668 6020
rect 17500 5966 17502 6018
rect 17554 5966 17668 6018
rect 17500 5964 17668 5966
rect 18508 6692 18564 6702
rect 18508 6130 18564 6636
rect 18732 6690 18788 6972
rect 18732 6638 18734 6690
rect 18786 6638 18788 6690
rect 18732 6626 18788 6638
rect 18844 7698 19124 7700
rect 18844 7646 19070 7698
rect 19122 7646 19124 7698
rect 18844 7644 19124 7646
rect 18844 7252 18900 7644
rect 19068 7634 19124 7644
rect 19292 7588 19348 7598
rect 19292 7494 19348 7532
rect 18956 7476 19012 7486
rect 18956 7382 19012 7420
rect 18508 6078 18510 6130
rect 18562 6078 18564 6130
rect 17500 5954 17556 5964
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 18508 5236 18564 6078
rect 18844 6130 18900 7196
rect 19068 7028 19124 7038
rect 18956 6580 19012 6590
rect 18956 6486 19012 6524
rect 18844 6078 18846 6130
rect 18898 6078 18900 6130
rect 18844 6066 18900 6078
rect 19068 6018 19124 6972
rect 19404 6692 19460 7756
rect 19516 7476 19572 9100
rect 19628 7924 19684 9996
rect 19852 9716 19908 10334
rect 19964 10164 20020 10556
rect 19964 9938 20020 10108
rect 19964 9886 19966 9938
rect 20018 9886 20020 9938
rect 19964 9874 20020 9886
rect 19852 9650 19908 9660
rect 21420 9604 21476 9614
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 21420 8596 21476 9548
rect 21196 8540 21476 8596
rect 21532 9380 21588 10668
rect 21644 10498 21700 10510
rect 21644 10446 21646 10498
rect 21698 10446 21700 10498
rect 21644 10388 21700 10446
rect 21644 10322 21700 10332
rect 22764 10388 22820 12798
rect 22988 12850 23044 12862
rect 22988 12798 22990 12850
rect 23042 12798 23044 12850
rect 22988 12740 23044 12798
rect 23436 12740 23492 12750
rect 24332 12740 24388 12750
rect 22988 12738 23492 12740
rect 22988 12686 23438 12738
rect 23490 12686 23492 12738
rect 22988 12684 23492 12686
rect 23436 12674 23492 12684
rect 23772 12738 24388 12740
rect 23772 12686 24334 12738
rect 24386 12686 24388 12738
rect 23772 12684 24388 12686
rect 23324 12516 23380 12526
rect 23324 12402 23380 12460
rect 23324 12350 23326 12402
rect 23378 12350 23380 12402
rect 23324 12338 23380 12350
rect 23772 10722 23828 12684
rect 24332 12674 24388 12684
rect 24556 12516 24612 13132
rect 24220 12460 24612 12516
rect 24220 12402 24276 12460
rect 24220 12350 24222 12402
rect 24274 12350 24276 12402
rect 24220 12338 24276 12350
rect 24556 12292 24612 12302
rect 24668 12292 24724 13468
rect 24780 12964 24836 12974
rect 24780 12870 24836 12908
rect 24332 12290 24724 12292
rect 24332 12238 24558 12290
rect 24610 12238 24724 12290
rect 24332 12236 24724 12238
rect 24332 11394 24388 12236
rect 24556 12226 24612 12236
rect 24332 11342 24334 11394
rect 24386 11342 24388 11394
rect 24332 11330 24388 11342
rect 24668 11506 24724 11518
rect 24668 11454 24670 11506
rect 24722 11454 24724 11506
rect 23772 10670 23774 10722
rect 23826 10670 23828 10722
rect 23772 10658 23828 10670
rect 23996 11170 24052 11182
rect 23996 11118 23998 11170
rect 24050 11118 24052 11170
rect 22764 10322 22820 10332
rect 21756 9940 21812 9950
rect 21756 9826 21812 9884
rect 22204 9940 22260 9950
rect 22204 9846 22260 9884
rect 21756 9774 21758 9826
rect 21810 9774 21812 9826
rect 21756 9762 21812 9774
rect 23436 9716 23492 9726
rect 23436 9622 23492 9660
rect 21532 9324 22148 9380
rect 19628 7858 19684 7868
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19628 7476 19684 7486
rect 19516 7474 19684 7476
rect 19516 7422 19630 7474
rect 19682 7422 19684 7474
rect 19516 7420 19684 7422
rect 19516 6914 19572 7420
rect 19628 7410 19684 7420
rect 20188 7362 20244 7374
rect 20188 7310 20190 7362
rect 20242 7310 20244 7362
rect 19964 7252 20020 7262
rect 19964 7158 20020 7196
rect 20188 7252 20244 7310
rect 21084 7364 21140 7374
rect 21084 7270 21140 7308
rect 20748 7252 20804 7262
rect 20188 7196 20748 7252
rect 20188 7028 20244 7196
rect 20748 7158 20804 7196
rect 20188 6962 20244 6972
rect 20524 7028 20580 7038
rect 19516 6862 19518 6914
rect 19570 6862 19572 6914
rect 19516 6850 19572 6862
rect 20188 6804 20244 6814
rect 19292 6578 19348 6590
rect 19292 6526 19294 6578
rect 19346 6526 19348 6578
rect 19292 6468 19348 6526
rect 19292 6402 19348 6412
rect 19068 5966 19070 6018
rect 19122 5966 19124 6018
rect 19068 5954 19124 5966
rect 19404 5906 19460 6636
rect 19404 5854 19406 5906
rect 19458 5854 19460 5906
rect 19404 5842 19460 5854
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 18956 5794 19012 5806
rect 18956 5742 18958 5794
rect 19010 5742 19012 5794
rect 18956 5684 19012 5742
rect 19628 5684 19684 6638
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 18956 5628 19684 5684
rect 18508 4338 18564 5180
rect 20188 5234 20244 6748
rect 20300 6692 20356 6702
rect 20300 6466 20356 6636
rect 20524 6690 20580 6972
rect 20524 6638 20526 6690
rect 20578 6638 20580 6690
rect 20524 6626 20580 6638
rect 20636 6692 20692 6702
rect 20636 6598 20692 6636
rect 20300 6414 20302 6466
rect 20354 6414 20356 6466
rect 20300 6356 20356 6414
rect 20300 6290 20356 6300
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20748 6132 20804 6414
rect 21196 6468 21252 8540
rect 21532 7588 21588 9324
rect 22092 9266 22148 9324
rect 22092 9214 22094 9266
rect 22146 9214 22148 9266
rect 22092 9202 22148 9214
rect 22428 9042 22484 9054
rect 22428 8990 22430 9042
rect 22482 8990 22484 9042
rect 22428 8484 22484 8990
rect 22428 8418 22484 8428
rect 21308 7362 21364 7374
rect 21308 7310 21310 7362
rect 21362 7310 21364 7362
rect 21308 7140 21364 7310
rect 21308 7074 21364 7084
rect 21420 7252 21476 7262
rect 21420 6914 21476 7196
rect 21420 6862 21422 6914
rect 21474 6862 21476 6914
rect 21420 6850 21476 6862
rect 21308 6692 21364 6702
rect 21308 6598 21364 6636
rect 21196 6402 21252 6412
rect 20748 6066 20804 6076
rect 21532 6018 21588 7532
rect 23548 7532 23828 7588
rect 23324 7476 23380 7486
rect 23548 7476 23604 7532
rect 23324 7474 23604 7476
rect 23324 7422 23326 7474
rect 23378 7422 23604 7474
rect 23324 7420 23604 7422
rect 23324 7410 23380 7420
rect 21644 7364 21700 7374
rect 21644 6132 21700 7308
rect 23660 7362 23716 7374
rect 23660 7310 23662 7362
rect 23714 7310 23716 7362
rect 22764 7250 22820 7262
rect 22764 7198 22766 7250
rect 22818 7198 22820 7250
rect 22764 7140 22820 7198
rect 23100 7252 23156 7262
rect 23100 7250 23268 7252
rect 23100 7198 23102 7250
rect 23154 7198 23268 7250
rect 23100 7196 23268 7198
rect 23100 7186 23156 7196
rect 22764 7074 22820 7084
rect 23212 7028 23268 7196
rect 23548 7140 23604 7150
rect 23212 6972 23380 7028
rect 22204 6804 22260 6814
rect 22204 6710 22260 6748
rect 23212 6804 23268 6814
rect 22316 6690 22372 6702
rect 22316 6638 22318 6690
rect 22370 6638 22372 6690
rect 21980 6580 22036 6590
rect 21980 6486 22036 6524
rect 21756 6468 21812 6478
rect 22316 6468 22372 6638
rect 21756 6374 21812 6412
rect 22092 6412 22316 6468
rect 21644 6038 21700 6076
rect 21532 5966 21534 6018
rect 21586 5966 21588 6018
rect 21532 5954 21588 5966
rect 22092 6018 22148 6412
rect 22316 6402 22372 6412
rect 22092 5966 22094 6018
rect 22146 5966 22148 6018
rect 21756 5908 21812 5918
rect 21756 5814 21812 5852
rect 20188 5182 20190 5234
rect 20242 5182 20244 5234
rect 20188 5170 20244 5182
rect 21308 5796 21364 5806
rect 20076 4900 20132 4910
rect 19180 4898 20132 4900
rect 19180 4846 20078 4898
rect 20130 4846 20132 4898
rect 19180 4844 20132 4846
rect 19180 4450 19236 4844
rect 20076 4834 20132 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19180 4398 19182 4450
rect 19234 4398 19236 4450
rect 19180 4386 19236 4398
rect 18508 4286 18510 4338
rect 18562 4286 18564 4338
rect 18508 4274 18564 4286
rect 21308 4226 21364 5740
rect 22092 5796 22148 5966
rect 22092 5730 22148 5740
rect 21420 5236 21476 5246
rect 21476 5180 21700 5236
rect 21420 5142 21476 5180
rect 21308 4174 21310 4226
rect 21362 4174 21364 4226
rect 21308 4162 21364 4174
rect 21644 4338 21700 5180
rect 23212 5234 23268 6748
rect 23324 6692 23380 6972
rect 23548 6914 23604 7084
rect 23548 6862 23550 6914
rect 23602 6862 23604 6914
rect 23548 6850 23604 6862
rect 23324 6020 23380 6636
rect 23436 6690 23492 6702
rect 23436 6638 23438 6690
rect 23490 6638 23492 6690
rect 23436 6132 23492 6638
rect 23660 6468 23716 7310
rect 23660 6402 23716 6412
rect 23772 7364 23828 7532
rect 23660 6132 23716 6142
rect 23436 6130 23716 6132
rect 23436 6078 23662 6130
rect 23714 6078 23716 6130
rect 23436 6076 23716 6078
rect 23660 6066 23716 6076
rect 23772 6130 23828 7308
rect 23884 7250 23940 7262
rect 23884 7198 23886 7250
rect 23938 7198 23940 7250
rect 23884 7028 23940 7198
rect 23884 6962 23940 6972
rect 23884 6468 23940 6478
rect 23884 6374 23940 6412
rect 23772 6078 23774 6130
rect 23826 6078 23828 6130
rect 23772 6066 23828 6078
rect 23996 6356 24052 11118
rect 24556 10612 24612 10622
rect 24556 10518 24612 10556
rect 24668 10164 24724 11454
rect 24332 7476 24388 7486
rect 24668 7476 24724 10108
rect 25004 9940 25060 18060
rect 25340 17444 25396 18398
rect 27132 18452 27188 19070
rect 27468 18676 27524 20078
rect 27468 18610 27524 18620
rect 27692 20132 27748 20142
rect 27132 18386 27188 18396
rect 25340 17378 25396 17388
rect 27580 17108 27636 17118
rect 27580 17014 27636 17052
rect 27692 16882 27748 20076
rect 27916 20018 27972 20030
rect 27916 19966 27918 20018
rect 27970 19966 27972 20018
rect 27916 17444 27972 19966
rect 28252 20020 28308 20526
rect 29036 20188 29092 20750
rect 29372 20802 29428 20860
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 29372 20738 29428 20750
rect 29260 20578 29316 20590
rect 29260 20526 29262 20578
rect 29314 20526 29316 20578
rect 29260 20188 29316 20526
rect 29596 20468 29652 26124
rect 30156 25508 30212 26238
rect 30268 26068 30324 26078
rect 30268 25974 30324 26012
rect 30156 25442 30212 25452
rect 30940 25396 30996 25406
rect 31052 25396 31108 27916
rect 31276 27858 31332 28812
rect 31388 27972 31444 29036
rect 31724 28756 31780 29260
rect 31948 28756 32004 28766
rect 31724 28754 32004 28756
rect 31724 28702 31950 28754
rect 32002 28702 32004 28754
rect 31724 28700 32004 28702
rect 31948 28690 32004 28700
rect 31388 27906 31444 27916
rect 31836 28532 31892 28542
rect 31276 27806 31278 27858
rect 31330 27806 31332 27858
rect 31276 27794 31332 27806
rect 31500 27860 31556 27870
rect 31500 27766 31556 27804
rect 31612 27748 31668 27758
rect 31612 27746 31780 27748
rect 31612 27694 31614 27746
rect 31666 27694 31780 27746
rect 31612 27692 31780 27694
rect 31612 27682 31668 27692
rect 31724 27186 31780 27692
rect 31724 27134 31726 27186
rect 31778 27134 31780 27186
rect 31724 27122 31780 27134
rect 31836 26516 31892 28476
rect 32060 27972 32116 27982
rect 32060 27878 32116 27916
rect 31836 26450 31892 26460
rect 30940 25394 31108 25396
rect 30940 25342 30942 25394
rect 30994 25342 31108 25394
rect 30940 25340 31108 25342
rect 30940 25330 30996 25340
rect 29708 25282 29764 25294
rect 29708 25230 29710 25282
rect 29762 25230 29764 25282
rect 29708 24612 29764 25230
rect 31276 25282 31332 25294
rect 31276 25230 31278 25282
rect 31330 25230 31332 25282
rect 29932 25172 29988 25182
rect 29932 24946 29988 25116
rect 29932 24894 29934 24946
rect 29986 24894 29988 24946
rect 29932 24882 29988 24894
rect 31276 24948 31332 25230
rect 32284 25172 32340 30156
rect 33180 30212 33236 38612
rect 33516 37268 33572 37278
rect 33516 37174 33572 37212
rect 33292 36482 33348 36494
rect 33292 36430 33294 36482
rect 33346 36430 33348 36482
rect 33292 36148 33348 36430
rect 33292 36082 33348 36092
rect 33628 35586 33684 35598
rect 33628 35534 33630 35586
rect 33682 35534 33684 35586
rect 33628 34132 33684 35534
rect 33628 33346 33684 34076
rect 33628 33294 33630 33346
rect 33682 33294 33684 33346
rect 33628 33282 33684 33294
rect 33740 35026 33796 38612
rect 33964 37940 34020 41134
rect 34636 41186 34692 41198
rect 35532 41188 35588 41198
rect 34636 41134 34638 41186
rect 34690 41134 34692 41186
rect 34188 41076 34244 41086
rect 34188 40404 34244 41020
rect 34636 40516 34692 41134
rect 34972 41186 35588 41188
rect 34972 41134 35534 41186
rect 35586 41134 35588 41186
rect 34972 41132 35588 41134
rect 34748 41076 34804 41086
rect 34748 40982 34804 41020
rect 34972 40962 35028 41132
rect 34972 40910 34974 40962
rect 35026 40910 35028 40962
rect 34860 40516 34916 40526
rect 34636 40514 34916 40516
rect 34636 40462 34862 40514
rect 34914 40462 34916 40514
rect 34636 40460 34916 40462
rect 34188 40402 34692 40404
rect 34188 40350 34190 40402
rect 34242 40350 34692 40402
rect 34188 40348 34692 40350
rect 34188 40338 34244 40348
rect 34636 39730 34692 40348
rect 34636 39678 34638 39730
rect 34690 39678 34692 39730
rect 34076 38834 34132 38846
rect 34076 38782 34078 38834
rect 34130 38782 34132 38834
rect 34076 38500 34132 38782
rect 34076 38434 34132 38444
rect 34300 38722 34356 38734
rect 34300 38670 34302 38722
rect 34354 38670 34356 38722
rect 33964 37874 34020 37884
rect 33852 37266 33908 37278
rect 33852 37214 33854 37266
rect 33906 37214 33908 37266
rect 33852 35700 33908 37214
rect 34300 37268 34356 38670
rect 34300 37202 34356 37212
rect 34412 38050 34468 38062
rect 34412 37998 34414 38050
rect 34466 37998 34468 38050
rect 34412 37380 34468 37998
rect 34076 37156 34132 37166
rect 33964 35700 34020 35710
rect 33852 35644 33964 35700
rect 33740 34974 33742 35026
rect 33794 34974 33796 35026
rect 33740 32788 33796 34974
rect 33852 34018 33908 34030
rect 33852 33966 33854 34018
rect 33906 33966 33908 34018
rect 33852 33348 33908 33966
rect 33852 33282 33908 33292
rect 33964 32788 34020 35644
rect 34076 34354 34132 37100
rect 34188 35588 34244 35598
rect 34188 35494 34244 35532
rect 34076 34302 34078 34354
rect 34130 34302 34132 34354
rect 34076 34290 34132 34302
rect 34188 34130 34244 34142
rect 34188 34078 34190 34130
rect 34242 34078 34244 34130
rect 34188 33796 34244 34078
rect 34412 34020 34468 37324
rect 34412 33954 34468 33964
rect 34524 37828 34580 37838
rect 34524 33796 34580 37772
rect 34636 37380 34692 39678
rect 34860 39618 34916 40460
rect 34972 40516 35028 40910
rect 35084 40964 35140 40974
rect 35084 40870 35140 40908
rect 35532 40516 35588 41132
rect 35756 41186 35812 41198
rect 35756 41134 35758 41186
rect 35810 41134 35812 41186
rect 35644 40964 35700 40974
rect 35756 40964 35812 41134
rect 35700 40908 35812 40964
rect 35644 40898 35700 40908
rect 35644 40516 35700 40526
rect 35532 40514 35700 40516
rect 35532 40462 35646 40514
rect 35698 40462 35700 40514
rect 35532 40460 35700 40462
rect 34972 40450 35028 40460
rect 35644 40450 35700 40460
rect 35756 40402 35812 40908
rect 35756 40350 35758 40402
rect 35810 40350 35812 40402
rect 35756 40338 35812 40350
rect 35868 40290 35924 41916
rect 36092 41188 36148 41198
rect 36092 41094 36148 41132
rect 35868 40238 35870 40290
rect 35922 40238 35924 40290
rect 35868 40226 35924 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 39732 35252 39742
rect 35196 39638 35252 39676
rect 34860 39566 34862 39618
rect 34914 39566 34916 39618
rect 34636 37314 34692 37324
rect 34748 38834 34804 38846
rect 34748 38782 34750 38834
rect 34802 38782 34804 38834
rect 34748 38724 34804 38782
rect 34748 35028 34804 38668
rect 34860 38722 34916 39566
rect 34860 38670 34862 38722
rect 34914 38670 34916 38722
rect 34860 38658 34916 38670
rect 36540 38946 36596 38958
rect 36540 38894 36542 38946
rect 36594 38894 36596 38946
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38276 35588 38286
rect 36540 38276 36596 38894
rect 36764 38948 36820 43932
rect 37100 43538 37156 43550
rect 37100 43486 37102 43538
rect 37154 43486 37156 43538
rect 37100 42978 37156 43486
rect 37436 43540 37492 46620
rect 37660 46676 37716 46686
rect 37548 46564 37604 46574
rect 37548 45892 37604 46508
rect 37548 45798 37604 45836
rect 37660 43762 37716 46620
rect 38220 46340 38276 50372
rect 38556 49924 38612 50372
rect 38556 49858 38612 49868
rect 38668 49810 38724 51212
rect 39340 50428 39396 63868
rect 39452 63858 39508 63868
rect 39452 62580 39508 62590
rect 39452 62466 39508 62524
rect 39452 62414 39454 62466
rect 39506 62414 39508 62466
rect 39452 62402 39508 62414
rect 40124 62188 40180 65212
rect 41356 64818 41412 64830
rect 41356 64766 41358 64818
rect 41410 64766 41412 64818
rect 41356 64708 41412 64766
rect 41692 64708 41748 64718
rect 41356 64706 41748 64708
rect 41356 64654 41694 64706
rect 41746 64654 41748 64706
rect 41356 64652 41748 64654
rect 41692 64642 41748 64652
rect 41580 64148 41636 64158
rect 41580 64054 41636 64092
rect 41244 63138 41300 63150
rect 41244 63086 41246 63138
rect 41298 63086 41300 63138
rect 41020 63028 41076 63038
rect 41020 62934 41076 62972
rect 41244 62356 41300 63086
rect 41804 63028 41860 65324
rect 42028 64148 42084 65324
rect 42700 64930 42756 65436
rect 44380 65492 44436 65502
rect 44828 65492 44884 65502
rect 44380 65490 44996 65492
rect 44380 65438 44382 65490
rect 44434 65438 44830 65490
rect 44882 65438 44996 65490
rect 44380 65436 44996 65438
rect 43708 65380 43764 65390
rect 42700 64878 42702 64930
rect 42754 64878 42756 64930
rect 42700 64866 42756 64878
rect 43596 65378 43764 65380
rect 43596 65326 43710 65378
rect 43762 65326 43764 65378
rect 43596 65324 43764 65326
rect 42028 64146 42196 64148
rect 42028 64094 42030 64146
rect 42082 64094 42196 64146
rect 42028 64092 42196 64094
rect 42028 64082 42084 64092
rect 41804 62962 41860 62972
rect 41916 62916 41972 62926
rect 41916 62466 41972 62860
rect 41916 62414 41918 62466
rect 41970 62414 41972 62466
rect 41916 62402 41972 62414
rect 41244 62262 41300 62300
rect 39788 62132 40180 62188
rect 41020 62244 41076 62254
rect 41020 62150 41076 62188
rect 39452 59106 39508 59118
rect 39452 59054 39454 59106
rect 39506 59054 39508 59106
rect 39452 58996 39508 59054
rect 39452 58930 39508 58940
rect 39564 55188 39620 55198
rect 39564 54738 39620 55132
rect 39788 54964 39844 62132
rect 42028 61460 42084 61470
rect 41020 61348 41076 61358
rect 40012 61010 40068 61022
rect 40012 60958 40014 61010
rect 40066 60958 40068 61010
rect 39900 60788 39956 60798
rect 40012 60788 40068 60958
rect 40236 60788 40292 60798
rect 40012 60732 40236 60788
rect 39900 60694 39956 60732
rect 40236 60722 40292 60732
rect 41020 60674 41076 61292
rect 41020 60622 41022 60674
rect 41074 60622 41076 60674
rect 39900 60564 39956 60574
rect 39900 59218 39956 60508
rect 40236 60004 40292 60014
rect 41020 60004 41076 60622
rect 41356 60786 41412 60798
rect 41356 60734 41358 60786
rect 41410 60734 41412 60786
rect 41244 60004 41300 60014
rect 41020 60002 41300 60004
rect 41020 59950 41246 60002
rect 41298 59950 41300 60002
rect 41020 59948 41300 59950
rect 40012 59780 40068 59790
rect 40236 59780 40292 59948
rect 40012 59778 40292 59780
rect 40012 59726 40014 59778
rect 40066 59726 40292 59778
rect 40012 59724 40292 59726
rect 40012 59714 40068 59724
rect 39900 59166 39902 59218
rect 39954 59166 39956 59218
rect 39900 59154 39956 59166
rect 39788 54908 40180 54964
rect 39564 54686 39566 54738
rect 39618 54686 39620 54738
rect 39564 54674 39620 54686
rect 39788 54684 40068 54740
rect 39452 54628 39508 54638
rect 39452 54292 39508 54572
rect 39788 54626 39844 54684
rect 39788 54574 39790 54626
rect 39842 54574 39844 54626
rect 39788 54562 39844 54574
rect 39900 54514 39956 54526
rect 39900 54462 39902 54514
rect 39954 54462 39956 54514
rect 39452 54236 39844 54292
rect 39564 53732 39620 53742
rect 39452 53620 39508 53630
rect 39452 52274 39508 53564
rect 39452 52222 39454 52274
rect 39506 52222 39508 52274
rect 39452 52210 39508 52222
rect 39564 53506 39620 53676
rect 39788 53730 39844 54236
rect 39900 53842 39956 54462
rect 39900 53790 39902 53842
rect 39954 53790 39956 53842
rect 39900 53778 39956 53790
rect 39788 53678 39790 53730
rect 39842 53678 39844 53730
rect 39788 53666 39844 53678
rect 40012 53730 40068 54684
rect 40012 53678 40014 53730
rect 40066 53678 40068 53730
rect 39564 53454 39566 53506
rect 39618 53454 39620 53506
rect 39564 50428 39620 53454
rect 40012 53396 40068 53678
rect 40012 53330 40068 53340
rect 40124 52052 40180 54908
rect 40236 53732 40292 59724
rect 40684 59778 40740 59790
rect 40684 59726 40686 59778
rect 40738 59726 40740 59778
rect 40684 59556 40740 59726
rect 40796 59780 40852 59790
rect 40796 59686 40852 59724
rect 40908 59778 40964 59790
rect 40908 59726 40910 59778
rect 40962 59726 40964 59778
rect 40684 59490 40740 59500
rect 40348 59332 40404 59342
rect 40908 59332 40964 59726
rect 40348 59330 40964 59332
rect 40348 59278 40350 59330
rect 40402 59278 40910 59330
rect 40962 59278 40964 59330
rect 40348 59276 40964 59278
rect 40348 59266 40404 59276
rect 40908 59266 40964 59276
rect 41020 59108 41076 59118
rect 41020 59014 41076 59052
rect 41020 58548 41076 58558
rect 40460 55410 40516 55422
rect 40460 55358 40462 55410
rect 40514 55358 40516 55410
rect 40460 55076 40516 55358
rect 40460 55010 40516 55020
rect 40796 55186 40852 55198
rect 40796 55134 40798 55186
rect 40850 55134 40852 55186
rect 40796 54628 40852 55134
rect 40796 54562 40852 54572
rect 41020 54738 41076 58492
rect 41020 54686 41022 54738
rect 41074 54686 41076 54738
rect 41020 54068 41076 54686
rect 41020 54002 41076 54012
rect 41132 58324 41188 59948
rect 41244 59938 41300 59948
rect 41244 59556 41300 59566
rect 41244 59220 41300 59500
rect 41244 59126 41300 59164
rect 41356 58546 41412 60734
rect 41468 60564 41524 60574
rect 41468 60470 41524 60508
rect 41916 60564 41972 60574
rect 41468 59780 41524 59790
rect 41468 59330 41524 59724
rect 41468 59278 41470 59330
rect 41522 59278 41524 59330
rect 41468 59266 41524 59278
rect 41804 59444 41860 59454
rect 41916 59444 41972 60508
rect 42028 59892 42084 61404
rect 42140 60116 42196 64092
rect 43372 63924 43428 63934
rect 43372 63830 43428 63868
rect 43036 63700 43092 63710
rect 43372 63700 43428 63710
rect 43596 63700 43652 65324
rect 43708 65314 43764 65324
rect 44380 65380 44436 65436
rect 44828 65426 44884 65436
rect 44380 65314 44436 65324
rect 44940 64820 44996 65436
rect 45612 65380 45668 65390
rect 45500 65378 45668 65380
rect 45500 65326 45614 65378
rect 45666 65326 45668 65378
rect 45500 65324 45668 65326
rect 45388 64820 45444 64830
rect 44940 64818 45444 64820
rect 44940 64766 44942 64818
rect 44994 64766 45390 64818
rect 45442 64766 45444 64818
rect 44940 64764 45444 64766
rect 44940 64754 44996 64764
rect 45388 64754 45444 64764
rect 44940 64148 44996 64158
rect 44828 64036 44884 64046
rect 43036 63698 43316 63700
rect 43036 63646 43038 63698
rect 43090 63646 43316 63698
rect 43036 63644 43316 63646
rect 43036 63634 43092 63644
rect 42252 63026 42308 63038
rect 42252 62974 42254 63026
rect 42306 62974 42308 63026
rect 42252 62244 42308 62974
rect 42252 62178 42308 62188
rect 42476 62914 42532 62926
rect 42476 62862 42478 62914
rect 42530 62862 42532 62914
rect 42476 62356 42532 62862
rect 42924 62916 42980 62926
rect 42924 62822 42980 62860
rect 43260 62466 43316 63644
rect 43372 63698 43652 63700
rect 43372 63646 43374 63698
rect 43426 63646 43652 63698
rect 43372 63644 43652 63646
rect 43820 63924 43876 63934
rect 43372 63634 43428 63644
rect 43484 63140 43540 63150
rect 43484 63046 43540 63084
rect 43260 62414 43262 62466
rect 43314 62414 43316 62466
rect 43260 62402 43316 62414
rect 42700 62356 42756 62366
rect 42476 62300 42700 62356
rect 42476 62242 42532 62300
rect 42700 62290 42756 62300
rect 42812 62356 42868 62366
rect 43484 62356 43540 62366
rect 42812 62354 43204 62356
rect 42812 62302 42814 62354
rect 42866 62302 43204 62354
rect 42812 62300 43204 62302
rect 42812 62290 42868 62300
rect 42476 62190 42478 62242
rect 42530 62190 42532 62242
rect 42476 62178 42532 62190
rect 43148 62188 43204 62300
rect 43484 62262 43540 62300
rect 43596 62244 43652 62254
rect 43148 62132 43428 62188
rect 43372 61794 43428 62132
rect 43372 61742 43374 61794
rect 43426 61742 43428 61794
rect 43372 61730 43428 61742
rect 43372 61572 43428 61582
rect 43596 61572 43652 62188
rect 43372 61570 43652 61572
rect 43372 61518 43374 61570
rect 43426 61518 43652 61570
rect 43372 61516 43652 61518
rect 42700 61012 42756 61022
rect 43372 61012 43428 61516
rect 43708 61460 43764 61470
rect 43708 61366 43764 61404
rect 42700 61010 43428 61012
rect 42700 60958 42702 61010
rect 42754 60958 43428 61010
rect 42700 60956 43428 60958
rect 42700 60946 42756 60956
rect 42476 60786 42532 60798
rect 42476 60734 42478 60786
rect 42530 60734 42532 60786
rect 42476 60564 42532 60734
rect 42476 60498 42532 60508
rect 42812 60562 42868 60574
rect 42812 60510 42814 60562
rect 42866 60510 42868 60562
rect 42476 60116 42532 60126
rect 42140 60114 42532 60116
rect 42140 60062 42478 60114
rect 42530 60062 42532 60114
rect 42140 60060 42532 60062
rect 42028 59836 42308 59892
rect 41916 59388 42084 59444
rect 41804 59220 41860 59388
rect 41916 59220 41972 59230
rect 41804 59218 41972 59220
rect 41804 59166 41918 59218
rect 41970 59166 41972 59218
rect 41804 59164 41972 59166
rect 42028 59220 42084 59388
rect 42252 59442 42308 59836
rect 42252 59390 42254 59442
rect 42306 59390 42308 59442
rect 42252 59378 42308 59390
rect 42364 59332 42420 59342
rect 42364 59238 42420 59276
rect 42140 59220 42196 59230
rect 42028 59218 42196 59220
rect 42028 59166 42142 59218
rect 42194 59166 42196 59218
rect 42028 59164 42196 59166
rect 41916 58996 41972 59164
rect 42140 59154 42196 59164
rect 41916 58930 41972 58940
rect 41356 58494 41358 58546
rect 41410 58494 41412 58546
rect 41356 58482 41412 58494
rect 41804 58548 41860 58558
rect 41804 58454 41860 58492
rect 42364 58548 42420 58558
rect 42476 58548 42532 60060
rect 42812 59444 42868 60510
rect 42812 59378 42868 59388
rect 43036 59332 43092 59342
rect 43092 59276 43204 59332
rect 43036 59238 43092 59276
rect 42420 58492 42532 58548
rect 42588 59220 42644 59230
rect 42924 59220 42980 59230
rect 42588 59218 42980 59220
rect 42588 59166 42590 59218
rect 42642 59166 42926 59218
rect 42978 59166 42980 59218
rect 42588 59164 42980 59166
rect 42364 58482 42420 58492
rect 42588 58324 42644 59164
rect 42924 59154 42980 59164
rect 43148 58658 43204 59276
rect 43260 59220 43316 59230
rect 43260 59126 43316 59164
rect 43820 59220 43876 63868
rect 44044 63140 44100 63150
rect 44044 63046 44100 63084
rect 44156 63028 44212 63038
rect 44156 62934 44212 62972
rect 44380 62916 44436 62926
rect 44380 62914 44772 62916
rect 44380 62862 44382 62914
rect 44434 62862 44772 62914
rect 44380 62860 44772 62862
rect 44380 62850 44436 62860
rect 44044 62580 44100 62590
rect 44044 62578 44660 62580
rect 44044 62526 44046 62578
rect 44098 62526 44660 62578
rect 44044 62524 44660 62526
rect 44044 62514 44100 62524
rect 43932 62356 43988 62366
rect 43932 62262 43988 62300
rect 44156 62354 44212 62366
rect 44156 62302 44158 62354
rect 44210 62302 44212 62354
rect 44156 61460 44212 62302
rect 44604 62356 44660 62524
rect 44716 62578 44772 62860
rect 44716 62526 44718 62578
rect 44770 62526 44772 62578
rect 44716 62514 44772 62526
rect 44828 62356 44884 63980
rect 44940 63140 44996 64092
rect 45164 63924 45220 63934
rect 45164 63250 45220 63868
rect 45500 63252 45556 65324
rect 45612 65314 45668 65324
rect 45164 63198 45166 63250
rect 45218 63198 45220 63250
rect 45164 63186 45220 63198
rect 45388 63196 45556 63252
rect 45612 64260 45668 64270
rect 44940 63046 44996 63084
rect 45052 63028 45108 63038
rect 45052 62934 45108 62972
rect 45276 62916 45332 62926
rect 45276 62468 45332 62860
rect 45276 62402 45332 62412
rect 44604 62354 44884 62356
rect 44604 62302 44606 62354
rect 44658 62302 44884 62354
rect 44604 62300 44884 62302
rect 44940 62356 44996 62366
rect 44604 62290 44660 62300
rect 44940 62262 44996 62300
rect 45052 62354 45108 62366
rect 45052 62302 45054 62354
rect 45106 62302 45108 62354
rect 45052 62188 45108 62302
rect 45388 62356 45444 63196
rect 45612 63140 45668 64204
rect 46060 64036 46116 64074
rect 46060 63970 46116 63980
rect 45948 63924 46004 63934
rect 45948 63830 46004 63868
rect 46172 63476 46228 66108
rect 47404 66274 47460 66286
rect 47404 66222 47406 66274
rect 47458 66222 47460 66274
rect 46508 65380 46564 65390
rect 46508 64260 46564 65324
rect 46172 63420 46452 63476
rect 45500 63084 45668 63140
rect 46060 63140 46116 63150
rect 45500 63026 45556 63084
rect 46060 63046 46116 63084
rect 45836 63028 45892 63038
rect 45500 62974 45502 63026
rect 45554 62974 45556 63026
rect 45500 62962 45556 62974
rect 45612 63026 45892 63028
rect 45612 62974 45838 63026
rect 45890 62974 45892 63026
rect 45612 62972 45892 62974
rect 45612 62804 45668 62972
rect 45500 62748 45668 62804
rect 45500 62578 45556 62748
rect 45836 62692 45892 62972
rect 45836 62636 46340 62692
rect 45500 62526 45502 62578
rect 45554 62526 45556 62578
rect 45500 62514 45556 62526
rect 45612 62580 45668 62590
rect 45612 62578 46116 62580
rect 45612 62526 45614 62578
rect 45666 62526 46116 62578
rect 45612 62524 46116 62526
rect 45612 62514 45668 62524
rect 46060 62468 46116 62524
rect 46060 62402 46116 62412
rect 45724 62356 45780 62366
rect 45948 62356 46004 62366
rect 45388 62300 45668 62356
rect 44156 61394 44212 61404
rect 44940 62132 45108 62188
rect 45612 62188 45668 62300
rect 45780 62354 46004 62356
rect 45780 62302 45950 62354
rect 46002 62302 46004 62354
rect 45780 62300 46004 62302
rect 45724 62262 45780 62300
rect 45948 62290 46004 62300
rect 46284 62354 46340 62636
rect 46284 62302 46286 62354
rect 46338 62302 46340 62354
rect 46284 62290 46340 62302
rect 46172 62244 46228 62254
rect 46060 62242 46228 62244
rect 46060 62190 46174 62242
rect 46226 62190 46228 62242
rect 46060 62188 46228 62190
rect 46396 62188 46452 63420
rect 46508 63140 46564 64204
rect 46956 64260 47012 64270
rect 46956 64146 47012 64204
rect 46956 64094 46958 64146
rect 47010 64094 47012 64146
rect 46956 64082 47012 64094
rect 46956 63922 47012 63934
rect 46956 63870 46958 63922
rect 47010 63870 47012 63922
rect 46508 63138 46900 63140
rect 46508 63086 46510 63138
rect 46562 63086 46900 63138
rect 46508 63084 46900 63086
rect 46508 63074 46564 63084
rect 46508 62468 46564 62478
rect 46508 62354 46564 62412
rect 46508 62302 46510 62354
rect 46562 62302 46564 62354
rect 46508 62290 46564 62302
rect 46844 62356 46900 63084
rect 46956 62580 47012 63870
rect 47292 63140 47348 63150
rect 47180 62916 47236 62926
rect 47180 62822 47236 62860
rect 47180 62580 47236 62590
rect 46956 62578 47236 62580
rect 46956 62526 47182 62578
rect 47234 62526 47236 62578
rect 46956 62524 47236 62526
rect 47180 62514 47236 62524
rect 47292 62466 47348 63084
rect 47292 62414 47294 62466
rect 47346 62414 47348 62466
rect 47292 62402 47348 62414
rect 46956 62356 47012 62366
rect 46844 62354 47012 62356
rect 46844 62302 46958 62354
rect 47010 62302 47012 62354
rect 46844 62300 47012 62302
rect 46956 62290 47012 62300
rect 47404 62188 47460 66222
rect 47516 64930 47572 67172
rect 48412 66500 48468 66510
rect 48412 66406 48468 66444
rect 49084 66500 49140 69200
rect 49084 66434 49140 66444
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 51100 65604 51156 69200
rect 52220 66500 52276 66510
rect 52220 66406 52276 66444
rect 53116 66500 53172 69200
rect 53116 66434 53172 66444
rect 51100 65538 51156 65548
rect 51212 66274 51268 66286
rect 51212 66222 51214 66274
rect 51266 66222 51268 66274
rect 48860 65490 48916 65502
rect 48860 65438 48862 65490
rect 48914 65438 48916 65490
rect 47740 65380 47796 65390
rect 47740 65286 47796 65324
rect 47516 64878 47518 64930
rect 47570 64878 47572 64930
rect 47516 64866 47572 64878
rect 47516 64372 47572 64382
rect 47572 64316 47684 64372
rect 47516 64306 47572 64316
rect 45612 62132 46116 62188
rect 46172 62178 46228 62188
rect 46284 62132 46452 62188
rect 47180 62132 47460 62188
rect 44940 61346 44996 62132
rect 44940 61294 44942 61346
rect 44994 61294 44996 61346
rect 44268 60228 44324 60238
rect 44268 60134 44324 60172
rect 44940 60004 44996 61294
rect 44940 59938 44996 59948
rect 44156 59890 44212 59902
rect 44156 59838 44158 59890
rect 44210 59838 44212 59890
rect 44156 59444 44212 59838
rect 44156 59378 44212 59388
rect 43820 59154 43876 59164
rect 45276 59220 45332 59258
rect 45276 59154 45332 59164
rect 45724 59220 45780 59230
rect 45724 59126 45780 59164
rect 44940 58994 44996 59006
rect 44940 58942 44942 58994
rect 44994 58942 44996 58994
rect 43148 58606 43150 58658
rect 43202 58606 43204 58658
rect 43148 58594 43204 58606
rect 43260 58772 43316 58782
rect 40236 53618 40292 53676
rect 40236 53566 40238 53618
rect 40290 53566 40292 53618
rect 40236 53554 40292 53566
rect 40908 53620 40964 53630
rect 40908 53172 40964 53564
rect 41020 53508 41076 53518
rect 41020 53414 41076 53452
rect 41020 53172 41076 53182
rect 40908 53170 41076 53172
rect 40908 53118 41022 53170
rect 41074 53118 41076 53170
rect 40908 53116 41076 53118
rect 41020 53106 41076 53116
rect 40124 51986 40180 51996
rect 41020 51490 41076 51502
rect 41020 51438 41022 51490
rect 41074 51438 41076 51490
rect 40908 51156 40964 51166
rect 40684 51154 40964 51156
rect 40684 51102 40910 51154
rect 40962 51102 40964 51154
rect 40684 51100 40964 51102
rect 40684 50706 40740 51100
rect 40908 51090 40964 51100
rect 41020 50820 41076 51438
rect 41020 50754 41076 50764
rect 40684 50654 40686 50706
rect 40738 50654 40740 50706
rect 40684 50642 40740 50654
rect 39228 50372 39396 50428
rect 39452 50372 39620 50428
rect 39228 49924 39284 50372
rect 39228 49858 39284 49868
rect 39340 50036 39396 50046
rect 39340 49922 39396 49980
rect 39340 49870 39342 49922
rect 39394 49870 39396 49922
rect 39340 49858 39396 49870
rect 38668 49758 38670 49810
rect 38722 49758 38724 49810
rect 38668 49746 38724 49758
rect 38444 47460 38500 47470
rect 38444 47366 38500 47404
rect 39004 47458 39060 47470
rect 39004 47406 39006 47458
rect 39058 47406 39060 47458
rect 38556 47236 38612 47246
rect 38556 47142 38612 47180
rect 39004 47124 39060 47406
rect 39004 47058 39060 47068
rect 39116 47346 39172 47358
rect 39116 47294 39118 47346
rect 39170 47294 39172 47346
rect 38892 46676 38948 46686
rect 39116 46676 39172 47294
rect 38948 46620 39172 46676
rect 38892 46582 38948 46620
rect 38220 46274 38276 46284
rect 37996 45890 38052 45902
rect 37996 45838 37998 45890
rect 38050 45838 38052 45890
rect 37996 45668 38052 45838
rect 38892 45890 38948 45902
rect 38892 45838 38894 45890
rect 38946 45838 38948 45890
rect 37996 45602 38052 45612
rect 38444 45668 38500 45678
rect 38444 45330 38500 45612
rect 38444 45278 38446 45330
rect 38498 45278 38500 45330
rect 38444 45266 38500 45278
rect 38892 45332 38948 45838
rect 38892 44324 38948 45276
rect 38892 44258 38948 44268
rect 37660 43710 37662 43762
rect 37714 43710 37716 43762
rect 37660 43698 37716 43710
rect 37884 44098 37940 44110
rect 37884 44046 37886 44098
rect 37938 44046 37940 44098
rect 37436 43484 37716 43540
rect 37100 42926 37102 42978
rect 37154 42926 37156 42978
rect 37100 42914 37156 42926
rect 37548 42756 37604 42766
rect 37324 42754 37604 42756
rect 37324 42702 37550 42754
rect 37602 42702 37604 42754
rect 37324 42700 37604 42702
rect 37212 42642 37268 42654
rect 37212 42590 37214 42642
rect 37266 42590 37268 42642
rect 37100 42530 37156 42542
rect 37100 42478 37102 42530
rect 37154 42478 37156 42530
rect 36876 41972 36932 41982
rect 37100 41972 37156 42478
rect 36876 41970 37156 41972
rect 36876 41918 36878 41970
rect 36930 41918 37156 41970
rect 36876 41916 37156 41918
rect 36876 41748 36932 41916
rect 37212 41860 37268 42590
rect 36876 41682 36932 41692
rect 36988 41858 37268 41860
rect 36988 41806 37214 41858
rect 37266 41806 37268 41858
rect 36988 41804 37268 41806
rect 36988 41298 37044 41804
rect 37212 41794 37268 41804
rect 36988 41246 36990 41298
rect 37042 41246 37044 41298
rect 36988 41234 37044 41246
rect 36764 38882 36820 38892
rect 37100 41186 37156 41198
rect 37100 41134 37102 41186
rect 37154 41134 37156 41186
rect 37100 39732 37156 41134
rect 35532 38274 36596 38276
rect 35532 38222 35534 38274
rect 35586 38222 36596 38274
rect 35532 38220 36596 38222
rect 35532 38210 35588 38220
rect 35084 37938 35140 37950
rect 35084 37886 35086 37938
rect 35138 37886 35140 37938
rect 35084 36148 35140 37886
rect 35644 37940 35700 37950
rect 35644 37938 36260 37940
rect 35644 37886 35646 37938
rect 35698 37886 36260 37938
rect 35644 37884 36260 37886
rect 35644 37874 35700 37884
rect 35532 37826 35588 37838
rect 35532 37774 35534 37826
rect 35586 37774 35588 37826
rect 35532 37604 35588 37774
rect 35532 37538 35588 37548
rect 35756 37380 35812 37390
rect 35756 37286 35812 37324
rect 35644 37268 35700 37278
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35644 36706 35700 37212
rect 35980 37266 36036 37278
rect 35980 37214 35982 37266
rect 36034 37214 36036 37266
rect 35980 37044 36036 37214
rect 35980 36978 36036 36988
rect 35644 36654 35646 36706
rect 35698 36654 35700 36706
rect 35644 36642 35700 36654
rect 35532 36594 35588 36606
rect 35532 36542 35534 36594
rect 35586 36542 35588 36594
rect 35420 36484 35476 36494
rect 35420 36390 35476 36428
rect 35084 36082 35140 36092
rect 34748 34962 34804 34972
rect 34972 35810 35028 35822
rect 34972 35758 34974 35810
rect 35026 35758 35028 35810
rect 34636 34244 34692 34254
rect 34636 34242 34804 34244
rect 34636 34190 34638 34242
rect 34690 34190 34804 34242
rect 34636 34188 34804 34190
rect 34636 34178 34692 34188
rect 34188 33740 34692 33796
rect 34188 33572 34244 33582
rect 34076 32788 34132 32798
rect 33740 32732 33908 32788
rect 33964 32786 34132 32788
rect 33964 32734 34078 32786
rect 34130 32734 34132 32786
rect 33964 32732 34132 32734
rect 33180 30146 33236 30156
rect 33628 32452 33684 32462
rect 33516 28644 33572 28654
rect 33628 28644 33684 32396
rect 33572 28588 33684 28644
rect 33516 28578 33572 28588
rect 33852 28084 33908 32732
rect 34076 32722 34132 32732
rect 33964 32562 34020 32574
rect 33964 32510 33966 32562
rect 34018 32510 34020 32562
rect 33964 32340 34020 32510
rect 34188 32564 34244 33516
rect 34300 33348 34356 33358
rect 34300 33254 34356 33292
rect 34188 32562 34356 32564
rect 34188 32510 34190 32562
rect 34242 32510 34356 32562
rect 34188 32508 34356 32510
rect 34188 32498 34244 32508
rect 33964 32284 34244 32340
rect 34076 32116 34132 32126
rect 34076 30210 34132 32060
rect 34076 30158 34078 30210
rect 34130 30158 34132 30210
rect 34076 28754 34132 30158
rect 34076 28702 34078 28754
rect 34130 28702 34132 28754
rect 34076 28690 34132 28702
rect 34188 31778 34244 32284
rect 34300 32004 34356 32508
rect 34300 31938 34356 31948
rect 34524 32450 34580 32462
rect 34524 32398 34526 32450
rect 34578 32398 34580 32450
rect 34188 31726 34190 31778
rect 34242 31726 34244 31778
rect 34188 28420 34244 31726
rect 34300 31780 34356 31790
rect 34524 31780 34580 32398
rect 34356 31724 34580 31780
rect 34300 31686 34356 31724
rect 34636 30210 34692 33740
rect 34748 32452 34804 34188
rect 34972 34132 35028 35758
rect 35532 35700 35588 36542
rect 36092 36482 36148 36494
rect 36092 36430 36094 36482
rect 36146 36430 36148 36482
rect 36092 36372 36148 36430
rect 36092 36306 36148 36316
rect 35980 36148 36036 36158
rect 35868 35700 35924 35710
rect 35532 35698 35924 35700
rect 35532 35646 35870 35698
rect 35922 35646 35924 35698
rect 35532 35644 35924 35646
rect 35868 35364 35924 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35868 35298 35924 35308
rect 35196 35242 35460 35252
rect 35756 35028 35812 35038
rect 35756 34934 35812 34972
rect 34972 33572 35028 34076
rect 34972 33506 35028 33516
rect 35084 34804 35140 34814
rect 35084 33346 35140 34748
rect 35980 34242 36036 36092
rect 36204 35028 36260 37884
rect 36540 36484 36596 38220
rect 36876 38834 36932 38846
rect 36876 38782 36878 38834
rect 36930 38782 36932 38834
rect 36876 37828 36932 38782
rect 37100 38836 37156 39676
rect 37100 38770 37156 38780
rect 37324 38668 37380 42700
rect 37548 42690 37604 42700
rect 37660 42530 37716 43484
rect 37772 43538 37828 43550
rect 37772 43486 37774 43538
rect 37826 43486 37828 43538
rect 37772 42756 37828 43486
rect 37884 43428 37940 44046
rect 39452 43708 39508 50372
rect 41020 50036 41076 50046
rect 41020 49942 41076 49980
rect 41132 49476 41188 58268
rect 42476 58268 42644 58324
rect 43148 58436 43204 58446
rect 43148 58322 43204 58380
rect 43260 58436 43316 58716
rect 44828 58546 44884 58558
rect 44828 58494 44830 58546
rect 44882 58494 44884 58546
rect 44828 58436 44884 58494
rect 43260 58434 43428 58436
rect 43260 58382 43262 58434
rect 43314 58382 43428 58434
rect 43260 58380 43428 58382
rect 43260 58370 43316 58380
rect 43148 58270 43150 58322
rect 43202 58270 43204 58322
rect 42140 57650 42196 57662
rect 42140 57598 42142 57650
rect 42194 57598 42196 57650
rect 42140 56868 42196 57598
rect 42364 56980 42420 56990
rect 42476 56980 42532 58268
rect 43148 57764 43204 58270
rect 43260 57764 43316 57774
rect 42700 57762 43316 57764
rect 42700 57710 43262 57762
rect 43314 57710 43316 57762
rect 42700 57708 43316 57710
rect 42588 57540 42644 57550
rect 42588 57446 42644 57484
rect 42700 57204 42756 57708
rect 43260 57698 43316 57708
rect 43148 57540 43204 57550
rect 43372 57540 43428 58380
rect 44828 58370 44884 58380
rect 44940 57874 44996 58942
rect 45276 58994 45332 59006
rect 45276 58942 45278 58994
rect 45330 58942 45332 58994
rect 45276 58548 45332 58942
rect 45276 58482 45332 58492
rect 44940 57822 44942 57874
rect 44994 57822 44996 57874
rect 44940 57810 44996 57822
rect 43204 57484 43428 57540
rect 43596 57652 43652 57662
rect 43148 57446 43204 57484
rect 42364 56978 42532 56980
rect 42364 56926 42366 56978
rect 42418 56926 42532 56978
rect 42364 56924 42532 56926
rect 42588 57148 42756 57204
rect 42364 56914 42420 56924
rect 42252 56868 42308 56878
rect 42140 56812 42252 56868
rect 42252 56774 42308 56812
rect 42476 56756 42532 56766
rect 42588 56756 42644 57148
rect 42700 57036 43540 57092
rect 42700 56978 42756 57036
rect 42700 56926 42702 56978
rect 42754 56926 42756 56978
rect 42700 56914 42756 56926
rect 42476 56754 42644 56756
rect 42476 56702 42478 56754
rect 42530 56702 42644 56754
rect 42476 56700 42644 56702
rect 42924 56866 42980 56878
rect 42924 56814 42926 56866
rect 42978 56814 42980 56866
rect 42924 56756 42980 56814
rect 42476 56690 42532 56700
rect 41692 55972 41748 55982
rect 41580 55412 41636 55422
rect 41580 55318 41636 55356
rect 41468 55298 41524 55310
rect 41468 55246 41470 55298
rect 41522 55246 41524 55298
rect 41468 55076 41524 55246
rect 41468 55010 41524 55020
rect 41580 54740 41636 54750
rect 41244 54738 41636 54740
rect 41244 54686 41582 54738
rect 41634 54686 41636 54738
rect 41244 54684 41636 54686
rect 41244 53732 41300 54684
rect 41580 54674 41636 54684
rect 41692 54738 41748 55916
rect 42924 55972 42980 56700
rect 42924 55906 42980 55916
rect 43148 55522 43204 57036
rect 43260 56756 43316 56766
rect 43260 56662 43316 56700
rect 43484 56754 43540 57036
rect 43596 57090 43652 57596
rect 44492 57652 44548 57662
rect 44492 57558 44548 57596
rect 43596 57038 43598 57090
rect 43650 57038 43652 57090
rect 43596 57026 43652 57038
rect 43484 56702 43486 56754
rect 43538 56702 43540 56754
rect 43484 56690 43540 56702
rect 45500 55972 45556 55982
rect 45500 55878 45556 55916
rect 43148 55470 43150 55522
rect 43202 55470 43204 55522
rect 43148 55458 43204 55470
rect 45612 55858 45668 55870
rect 45612 55806 45614 55858
rect 45666 55806 45668 55858
rect 42140 55412 42196 55422
rect 42140 55318 42196 55356
rect 45612 55410 45668 55806
rect 45612 55358 45614 55410
rect 45666 55358 45668 55410
rect 45612 55346 45668 55358
rect 42364 55300 42420 55310
rect 42812 55300 42868 55310
rect 42252 55298 42868 55300
rect 42252 55246 42366 55298
rect 42418 55246 42814 55298
rect 42866 55246 42868 55298
rect 42252 55244 42868 55246
rect 41692 54686 41694 54738
rect 41746 54686 41748 54738
rect 41692 54674 41748 54686
rect 41804 54740 41860 54750
rect 41804 54646 41860 54684
rect 41468 54514 41524 54526
rect 41468 54462 41470 54514
rect 41522 54462 41524 54514
rect 41468 53956 41524 54462
rect 42028 54516 42084 54526
rect 42252 54516 42308 55244
rect 42364 55234 42420 55244
rect 42812 55234 42868 55244
rect 44268 55300 44324 55310
rect 42364 55076 42420 55086
rect 42364 54626 42420 55020
rect 43036 55074 43092 55086
rect 43036 55022 43038 55074
rect 43090 55022 43092 55074
rect 43036 54852 43092 55022
rect 42476 54796 43092 54852
rect 44268 55074 44324 55244
rect 44940 55300 44996 55310
rect 44940 55206 44996 55244
rect 44268 55022 44270 55074
rect 44322 55022 44324 55074
rect 42476 54740 42532 54796
rect 42476 54646 42532 54684
rect 42364 54574 42366 54626
rect 42418 54574 42420 54626
rect 42364 54562 42420 54574
rect 42028 54514 42308 54516
rect 42028 54462 42030 54514
rect 42082 54462 42308 54514
rect 42028 54460 42308 54462
rect 41468 53900 41748 53956
rect 41244 53676 41524 53732
rect 41244 53618 41300 53676
rect 41244 53566 41246 53618
rect 41298 53566 41300 53618
rect 41244 53554 41300 53566
rect 41468 53620 41524 53676
rect 41580 53620 41636 53630
rect 41468 53618 41636 53620
rect 41468 53566 41582 53618
rect 41634 53566 41636 53618
rect 41468 53564 41636 53566
rect 41580 53554 41636 53564
rect 41692 53618 41748 53900
rect 42028 53844 42084 54460
rect 42028 53778 42084 53788
rect 42476 54068 42532 54078
rect 41692 53566 41694 53618
rect 41746 53566 41748 53618
rect 41356 53506 41412 53518
rect 41356 53454 41358 53506
rect 41410 53454 41412 53506
rect 41356 53396 41412 53454
rect 41356 53330 41412 53340
rect 41692 52500 41748 53566
rect 41580 52444 41748 52500
rect 42476 52946 42532 54012
rect 44268 54068 44324 55022
rect 46284 54964 46340 62132
rect 47068 60002 47124 60014
rect 47068 59950 47070 60002
rect 47122 59950 47124 60002
rect 47068 59444 47124 59950
rect 47068 59378 47124 59388
rect 46956 58548 47012 58558
rect 46956 58454 47012 58492
rect 47068 57428 47124 57438
rect 47068 56978 47124 57372
rect 47068 56926 47070 56978
rect 47122 56926 47124 56978
rect 47068 56914 47124 56926
rect 46956 56308 47012 56318
rect 47180 56308 47236 62132
rect 46732 56306 47236 56308
rect 46732 56254 46958 56306
rect 47010 56254 47236 56306
rect 46732 56252 47236 56254
rect 47628 56308 47684 64316
rect 47740 63476 47796 63486
rect 47740 63250 47796 63420
rect 47740 63198 47742 63250
rect 47794 63198 47796 63250
rect 47740 63140 47796 63198
rect 47740 63074 47796 63084
rect 48860 62580 48916 65438
rect 49532 65380 49588 65390
rect 49532 65378 50260 65380
rect 49532 65326 49534 65378
rect 49586 65326 50260 65378
rect 49532 65324 50260 65326
rect 49532 65314 49588 65324
rect 50204 64930 50260 65324
rect 50204 64878 50206 64930
rect 50258 64878 50260 64930
rect 50204 64866 50260 64878
rect 48860 62354 48916 62524
rect 49420 64706 49476 64718
rect 49420 64654 49422 64706
rect 49474 64654 49476 64706
rect 49420 62356 49476 64654
rect 50316 64594 50372 64606
rect 50316 64542 50318 64594
rect 50370 64542 50372 64594
rect 50316 64148 50372 64542
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 51212 64260 51268 66222
rect 55020 66274 55076 66286
rect 55020 66222 55022 66274
rect 55074 66222 55076 66274
rect 52332 65492 52388 65502
rect 51660 65380 51716 65390
rect 50556 64250 50820 64260
rect 50988 64204 51268 64260
rect 51324 65378 51716 65380
rect 51324 65326 51662 65378
rect 51714 65326 51716 65378
rect 51324 65324 51716 65326
rect 50428 64148 50484 64158
rect 50316 64146 50484 64148
rect 50316 64094 50430 64146
rect 50482 64094 50484 64146
rect 50316 64092 50484 64094
rect 50428 64082 50484 64092
rect 50876 64036 50932 64046
rect 50764 64034 50932 64036
rect 50764 63982 50878 64034
rect 50930 63982 50932 64034
rect 50764 63980 50932 63982
rect 49532 63924 49588 63934
rect 49532 63830 49588 63868
rect 49644 63922 49700 63934
rect 49644 63870 49646 63922
rect 49698 63870 49700 63922
rect 49644 63140 49700 63870
rect 49980 63922 50036 63934
rect 49980 63870 49982 63922
rect 50034 63870 50036 63922
rect 49980 63252 50036 63870
rect 49980 63186 50036 63196
rect 50092 63922 50148 63934
rect 50092 63870 50094 63922
rect 50146 63870 50148 63922
rect 49644 63074 49700 63084
rect 48860 62302 48862 62354
rect 48914 62302 48916 62354
rect 48860 62290 48916 62302
rect 49084 62300 49476 62356
rect 49084 62188 49140 62300
rect 49532 62244 49588 62254
rect 48972 62132 49140 62188
rect 49196 62242 49588 62244
rect 49196 62190 49534 62242
rect 49586 62190 49588 62242
rect 49196 62188 49588 62190
rect 48860 61908 48916 61918
rect 48860 60786 48916 61852
rect 48860 60734 48862 60786
rect 48914 60734 48916 60786
rect 48860 60228 48916 60734
rect 48860 60162 48916 60172
rect 47740 59892 47796 59902
rect 47740 59890 48132 59892
rect 47740 59838 47742 59890
rect 47794 59838 48132 59890
rect 47740 59836 48132 59838
rect 47740 59826 47796 59836
rect 48076 59442 48132 59836
rect 48972 59668 49028 62132
rect 49196 61794 49252 62188
rect 49532 62178 49588 62188
rect 50092 62244 50148 63870
rect 49196 61742 49198 61794
rect 49250 61742 49252 61794
rect 49196 61730 49252 61742
rect 49084 61460 49140 61470
rect 49084 61458 49700 61460
rect 49084 61406 49086 61458
rect 49138 61406 49700 61458
rect 49084 61404 49700 61406
rect 49084 61394 49140 61404
rect 48860 59612 49028 59668
rect 49084 61012 49140 61022
rect 48076 59390 48078 59442
rect 48130 59390 48132 59442
rect 48076 59378 48132 59390
rect 48300 59444 48356 59454
rect 48188 59332 48244 59342
rect 48188 59238 48244 59276
rect 48188 58548 48244 58558
rect 48300 58548 48356 59388
rect 48860 59442 48916 59612
rect 48860 59390 48862 59442
rect 48914 59390 48916 59442
rect 47740 58546 48356 58548
rect 47740 58494 48190 58546
rect 48242 58494 48356 58546
rect 47740 58492 48356 58494
rect 48636 59220 48692 59230
rect 47740 58434 47796 58492
rect 48188 58482 48244 58492
rect 47740 58382 47742 58434
rect 47794 58382 47796 58434
rect 47740 58370 47796 58382
rect 48188 57428 48244 57438
rect 48076 57372 48188 57428
rect 46396 55972 46452 55982
rect 46452 55916 46676 55972
rect 46396 55906 46452 55916
rect 45948 54908 46340 54964
rect 44268 53732 44324 54012
rect 44268 53666 44324 53676
rect 45500 54740 45556 54750
rect 45948 54740 46004 54908
rect 45500 54738 46004 54740
rect 45500 54686 45502 54738
rect 45554 54686 45950 54738
rect 46002 54686 46004 54738
rect 45500 54684 46004 54686
rect 45500 53620 45556 54684
rect 45948 54674 46004 54684
rect 46620 54738 46676 55916
rect 46732 55412 46788 56252
rect 46956 56242 47012 56252
rect 47628 56242 47684 56252
rect 47964 56308 48020 56318
rect 47068 56082 47124 56094
rect 47068 56030 47070 56082
rect 47122 56030 47124 56082
rect 47068 55636 47124 56030
rect 46732 55346 46788 55356
rect 46844 55580 47124 55636
rect 47180 56082 47236 56094
rect 47180 56030 47182 56082
rect 47234 56030 47236 56082
rect 46620 54686 46622 54738
rect 46674 54686 46676 54738
rect 46620 54674 46676 54686
rect 46060 54628 46116 54638
rect 46060 54514 46116 54572
rect 46844 54628 46900 55580
rect 47180 55524 47236 56030
rect 46844 54562 46900 54572
rect 46956 55468 47236 55524
rect 47628 56082 47684 56094
rect 47628 56030 47630 56082
rect 47682 56030 47684 56082
rect 46956 55188 47012 55468
rect 47628 55412 47684 56030
rect 47852 55970 47908 55982
rect 47852 55918 47854 55970
rect 47906 55918 47908 55970
rect 47740 55412 47796 55422
rect 47628 55410 47796 55412
rect 47628 55358 47742 55410
rect 47794 55358 47796 55410
rect 47628 55356 47796 55358
rect 46060 54462 46062 54514
rect 46114 54462 46116 54514
rect 45500 53554 45556 53564
rect 45836 53732 45892 53742
rect 45836 53170 45892 53676
rect 45836 53118 45838 53170
rect 45890 53118 45892 53170
rect 45836 53106 45892 53118
rect 42476 52894 42478 52946
rect 42530 52894 42532 52946
rect 41580 51378 41636 52444
rect 42476 51604 42532 52894
rect 43260 52834 43316 52846
rect 43260 52782 43262 52834
rect 43314 52782 43316 52834
rect 43260 52274 43316 52782
rect 43260 52222 43262 52274
rect 43314 52222 43316 52274
rect 43260 52210 43316 52222
rect 43820 52836 43876 52846
rect 43820 52162 43876 52780
rect 45388 52834 45444 52846
rect 45388 52782 45390 52834
rect 45442 52782 45444 52834
rect 45388 52724 45444 52782
rect 45612 52724 45668 52734
rect 45388 52722 45668 52724
rect 45388 52670 45614 52722
rect 45666 52670 45668 52722
rect 45388 52668 45668 52670
rect 45612 52658 45668 52668
rect 43820 52110 43822 52162
rect 43874 52110 43876 52162
rect 43820 52098 43876 52110
rect 45500 52276 45556 52286
rect 43148 52052 43204 52062
rect 43148 51958 43204 51996
rect 44156 52052 44212 52062
rect 43372 51938 43428 51950
rect 43372 51886 43374 51938
rect 43426 51886 43428 51938
rect 42476 51538 42532 51548
rect 43260 51604 43316 51614
rect 43260 51510 43316 51548
rect 41692 51492 41748 51502
rect 41692 51490 41860 51492
rect 41692 51438 41694 51490
rect 41746 51438 41860 51490
rect 41692 51436 41860 51438
rect 41692 51426 41748 51436
rect 41580 51326 41582 51378
rect 41634 51326 41636 51378
rect 41244 51156 41300 51166
rect 41244 51062 41300 51100
rect 41468 50596 41524 50606
rect 41468 50502 41524 50540
rect 41580 50428 41636 51326
rect 41804 51268 41860 51436
rect 43260 51380 43316 51390
rect 41804 51202 41860 51212
rect 42252 51268 42308 51278
rect 42252 51174 42308 51212
rect 41692 51156 41748 51166
rect 41692 51062 41748 51100
rect 41804 50820 41860 50830
rect 41804 50726 41860 50764
rect 41916 50594 41972 50606
rect 41916 50542 41918 50594
rect 41970 50542 41972 50594
rect 41916 50428 41972 50542
rect 41356 50372 41636 50428
rect 41804 50372 41972 50428
rect 42140 50594 42196 50606
rect 42140 50542 42142 50594
rect 42194 50542 42196 50594
rect 41356 50034 41412 50372
rect 41356 49982 41358 50034
rect 41410 49982 41412 50034
rect 41356 49970 41412 49982
rect 41244 49810 41300 49822
rect 41244 49758 41246 49810
rect 41298 49758 41300 49810
rect 41244 49588 41300 49758
rect 41468 49812 41524 49822
rect 41468 49718 41524 49756
rect 41804 49698 41860 50372
rect 42140 50036 42196 50542
rect 42140 49970 42196 49980
rect 42252 50594 42308 50606
rect 42252 50542 42254 50594
rect 42306 50542 42308 50594
rect 41804 49646 41806 49698
rect 41858 49646 41860 49698
rect 41804 49588 41860 49646
rect 41244 49532 41860 49588
rect 41916 49922 41972 49934
rect 41916 49870 41918 49922
rect 41970 49870 41972 49922
rect 41132 49420 41412 49476
rect 41132 47234 41188 47246
rect 41132 47182 41134 47234
rect 41186 47182 41188 47234
rect 39900 46788 39956 46798
rect 39900 46694 39956 46732
rect 41020 46786 41076 46798
rect 41020 46734 41022 46786
rect 41074 46734 41076 46786
rect 41020 46564 41076 46734
rect 41132 46788 41188 47182
rect 41244 46788 41300 46798
rect 41132 46786 41300 46788
rect 41132 46734 41246 46786
rect 41298 46734 41300 46786
rect 41132 46732 41300 46734
rect 41244 46722 41300 46732
rect 39564 46452 39620 46462
rect 39564 46002 39620 46396
rect 40908 46452 40964 46462
rect 40908 46358 40964 46396
rect 39564 45950 39566 46002
rect 39618 45950 39620 46002
rect 39564 45938 39620 45950
rect 40796 44324 40852 44334
rect 40796 44230 40852 44268
rect 41020 43708 41076 46508
rect 38556 43650 38612 43662
rect 39452 43652 39844 43708
rect 38556 43598 38558 43650
rect 38610 43598 38612 43650
rect 38220 43428 38276 43438
rect 37884 43426 38276 43428
rect 37884 43374 38222 43426
rect 38274 43374 38276 43426
rect 37884 43372 38276 43374
rect 37772 42690 37828 42700
rect 38108 42754 38164 43372
rect 38220 43362 38276 43372
rect 38108 42702 38110 42754
rect 38162 42702 38164 42754
rect 37660 42478 37662 42530
rect 37714 42478 37716 42530
rect 37660 42466 37716 42478
rect 38108 42196 38164 42702
rect 38556 42642 38612 43598
rect 39676 43538 39732 43550
rect 39676 43486 39678 43538
rect 39730 43486 39732 43538
rect 39676 42980 39732 43486
rect 39340 42924 39732 42980
rect 38556 42590 38558 42642
rect 38610 42590 38612 42642
rect 38164 42140 38276 42196
rect 38108 42130 38164 42140
rect 38220 41972 38276 42140
rect 38556 41972 38612 42590
rect 39228 42756 39284 42766
rect 39340 42756 39396 42924
rect 39228 42754 39396 42756
rect 39228 42702 39230 42754
rect 39282 42702 39396 42754
rect 39228 42700 39396 42702
rect 39452 42756 39508 42766
rect 39228 42084 39284 42700
rect 39228 42018 39284 42028
rect 38780 41972 38836 41982
rect 38276 41916 38500 41972
rect 38556 41970 38836 41972
rect 38556 41918 38782 41970
rect 38834 41918 38836 41970
rect 38556 41916 38836 41918
rect 38220 41906 38276 41916
rect 38108 41860 38164 41870
rect 38108 41766 38164 41804
rect 38444 41300 38500 41916
rect 38556 41300 38612 41310
rect 38444 41298 38612 41300
rect 38444 41246 38558 41298
rect 38610 41246 38612 41298
rect 38444 41244 38612 41246
rect 38556 41234 38612 41244
rect 37660 41188 37716 41198
rect 37660 41094 37716 41132
rect 38108 40516 38164 40526
rect 37884 40404 37940 40414
rect 37772 40402 37940 40404
rect 37772 40350 37886 40402
rect 37938 40350 37940 40402
rect 37772 40348 37940 40350
rect 37548 39508 37604 39518
rect 37772 39508 37828 40348
rect 37884 40338 37940 40348
rect 37548 39506 37828 39508
rect 37548 39454 37550 39506
rect 37602 39454 37828 39506
rect 37548 39452 37828 39454
rect 38108 40290 38164 40460
rect 38780 40514 38836 41916
rect 38892 41972 38948 41982
rect 38892 41858 38948 41916
rect 38892 41806 38894 41858
rect 38946 41806 38948 41858
rect 38892 41794 38948 41806
rect 39452 41858 39508 42700
rect 39452 41806 39454 41858
rect 39506 41806 39508 41858
rect 39452 41794 39508 41806
rect 38780 40462 38782 40514
rect 38834 40462 38836 40514
rect 38780 40450 38836 40462
rect 38108 40238 38110 40290
rect 38162 40238 38164 40290
rect 36876 37762 36932 37772
rect 36988 38612 37380 38668
rect 37436 38834 37492 38846
rect 37436 38782 37438 38834
rect 37490 38782 37492 38834
rect 36876 36708 36932 36718
rect 36988 36708 37044 38612
rect 37436 38052 37492 38782
rect 37548 38724 37604 39452
rect 37548 38658 37604 38668
rect 37884 39394 37940 39406
rect 37884 39342 37886 39394
rect 37938 39342 37940 39394
rect 37324 37996 37492 38052
rect 37884 38164 37940 39342
rect 38108 38946 38164 40238
rect 38108 38894 38110 38946
rect 38162 38894 38164 38946
rect 38108 38882 38164 38894
rect 39004 38948 39060 38958
rect 39004 38854 39060 38892
rect 39676 38834 39732 38846
rect 39676 38782 39678 38834
rect 39730 38782 39732 38834
rect 39228 38722 39284 38734
rect 39228 38670 39230 38722
rect 39282 38670 39284 38722
rect 37212 37940 37268 37950
rect 37212 37846 37268 37884
rect 37100 37492 37156 37530
rect 37100 37426 37156 37436
rect 36876 36706 37044 36708
rect 36876 36654 36878 36706
rect 36930 36654 37044 36706
rect 36876 36652 37044 36654
rect 37212 37378 37268 37390
rect 37212 37326 37214 37378
rect 37266 37326 37268 37378
rect 36876 36642 36932 36652
rect 37100 36484 37156 36494
rect 36540 36482 37156 36484
rect 36540 36430 37102 36482
rect 37154 36430 37156 36482
rect 36540 36428 37156 36430
rect 37100 36418 37156 36428
rect 37212 36484 37268 37326
rect 37324 36932 37380 37996
rect 37436 37828 37492 37838
rect 37436 37156 37492 37772
rect 37772 37380 37828 37390
rect 37772 37286 37828 37324
rect 37436 37100 37604 37156
rect 37324 36866 37380 36876
rect 37268 36428 37492 36484
rect 37212 36418 37268 36428
rect 36204 34914 36260 34972
rect 36204 34862 36206 34914
rect 36258 34862 36260 34914
rect 36204 34850 36260 34862
rect 36540 36148 36596 36158
rect 36540 35588 36596 36092
rect 35980 34190 35982 34242
rect 36034 34190 36036 34242
rect 35980 34178 36036 34190
rect 36540 34130 36596 35532
rect 37212 35810 37268 35822
rect 37212 35758 37214 35810
rect 37266 35758 37268 35810
rect 36988 35364 37044 35374
rect 36540 34078 36542 34130
rect 36594 34078 36596 34130
rect 36540 34066 36596 34078
rect 36764 34132 36820 34142
rect 36764 34038 36820 34076
rect 36876 34020 36932 34030
rect 36988 34020 37044 35308
rect 37212 35140 37268 35758
rect 37436 35810 37492 36428
rect 37548 36482 37604 37100
rect 37772 37044 37828 37054
rect 37548 36430 37550 36482
rect 37602 36430 37604 36482
rect 37548 36418 37604 36430
rect 37660 36932 37716 36942
rect 37660 36482 37716 36876
rect 37660 36430 37662 36482
rect 37714 36430 37716 36482
rect 37660 35922 37716 36430
rect 37660 35870 37662 35922
rect 37714 35870 37716 35922
rect 37660 35858 37716 35870
rect 37436 35758 37438 35810
rect 37490 35758 37492 35810
rect 37436 35746 37492 35758
rect 37548 35140 37604 35150
rect 37212 35084 37548 35140
rect 37212 34916 37268 34926
rect 37212 34914 37380 34916
rect 37212 34862 37214 34914
rect 37266 34862 37380 34914
rect 37212 34860 37380 34862
rect 37212 34850 37268 34860
rect 37100 34804 37156 34814
rect 37100 34242 37156 34748
rect 37100 34190 37102 34242
rect 37154 34190 37156 34242
rect 37100 34178 37156 34190
rect 36988 33964 37156 34020
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35084 33294 35086 33346
rect 35138 33294 35140 33346
rect 35084 33282 35140 33294
rect 34972 33124 35028 33134
rect 34748 31892 34804 32396
rect 34860 32676 34916 32686
rect 34860 32116 34916 32620
rect 34972 32562 35028 33068
rect 34972 32510 34974 32562
rect 35026 32510 35028 32562
rect 34972 32498 35028 32510
rect 36204 33122 36260 33134
rect 36204 33070 36206 33122
rect 36258 33070 36260 33122
rect 36204 32452 36260 33070
rect 36204 32228 36260 32396
rect 36876 32450 36932 33964
rect 36988 33346 37044 33358
rect 36988 33294 36990 33346
rect 37042 33294 37044 33346
rect 36988 32676 37044 33294
rect 37100 33124 37156 33964
rect 37100 33030 37156 33068
rect 37324 34018 37380 34860
rect 37324 33966 37326 34018
rect 37378 33966 37380 34018
rect 36988 32610 37044 32620
rect 37212 32788 37268 32798
rect 37212 32564 37268 32732
rect 36876 32398 36878 32450
rect 36930 32398 36932 32450
rect 36876 32386 36932 32398
rect 37100 32562 37268 32564
rect 37100 32510 37214 32562
rect 37266 32510 37268 32562
rect 37100 32508 37268 32510
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 36204 32162 36260 32172
rect 35196 32106 35460 32116
rect 34860 32050 34916 32060
rect 34748 31798 34804 31836
rect 35308 32004 35364 32014
rect 35196 31668 35252 31678
rect 34860 31612 35196 31668
rect 34860 31218 34916 31612
rect 35196 31574 35252 31612
rect 34860 31166 34862 31218
rect 34914 31166 34916 31218
rect 34860 30772 34916 31166
rect 35308 31106 35364 31948
rect 35756 32004 35812 32014
rect 35756 31910 35812 31948
rect 37100 31890 37156 32508
rect 37212 32498 37268 32508
rect 37212 32004 37268 32014
rect 37324 32004 37380 33966
rect 37436 34130 37492 34142
rect 37436 34078 37438 34130
rect 37490 34078 37492 34130
rect 37436 34020 37492 34078
rect 37436 33954 37492 33964
rect 37436 32564 37492 32574
rect 37548 32564 37604 35084
rect 37660 35028 37716 35038
rect 37772 35028 37828 36988
rect 37884 36594 37940 38108
rect 38780 38164 38836 38174
rect 38108 38050 38164 38062
rect 38108 37998 38110 38050
rect 38162 37998 38164 38050
rect 37996 37938 38052 37950
rect 37996 37886 37998 37938
rect 38050 37886 38052 37938
rect 37996 37492 38052 37886
rect 37996 37426 38052 37436
rect 37884 36542 37886 36594
rect 37938 36542 37940 36594
rect 37884 36530 37940 36542
rect 37996 37266 38052 37278
rect 37996 37214 37998 37266
rect 38050 37214 38052 37266
rect 37996 36372 38052 37214
rect 37660 35026 37828 35028
rect 37660 34974 37662 35026
rect 37714 34974 37828 35026
rect 37660 34972 37828 34974
rect 37884 35700 37940 35710
rect 37996 35700 38052 36316
rect 38108 35924 38164 37998
rect 38668 37940 38724 37950
rect 38668 36708 38724 37884
rect 38780 37380 38836 38108
rect 39004 37940 39060 37950
rect 38780 37044 38836 37324
rect 38892 37938 39060 37940
rect 38892 37886 39006 37938
rect 39058 37886 39060 37938
rect 38892 37884 39060 37886
rect 38892 37268 38948 37884
rect 39004 37874 39060 37884
rect 39228 37716 39284 38670
rect 39676 38612 39732 38782
rect 39676 38546 39732 38556
rect 39004 37660 39284 37716
rect 39004 37490 39060 37660
rect 39004 37438 39006 37490
rect 39058 37438 39060 37490
rect 39004 37426 39060 37438
rect 39564 37380 39620 37390
rect 39564 37286 39620 37324
rect 39676 37378 39732 37390
rect 39676 37326 39678 37378
rect 39730 37326 39732 37378
rect 39228 37268 39284 37278
rect 38892 37266 39284 37268
rect 38892 37214 39230 37266
rect 39282 37214 39284 37266
rect 38892 37212 39284 37214
rect 39228 37156 39284 37212
rect 39228 37090 39284 37100
rect 39676 37156 39732 37326
rect 39676 37090 39732 37100
rect 38892 37044 38948 37054
rect 38780 37042 38948 37044
rect 38780 36990 38894 37042
rect 38946 36990 38948 37042
rect 38780 36988 38948 36990
rect 38892 36978 38948 36988
rect 38668 36652 39060 36708
rect 38556 36484 38612 36494
rect 38556 36390 38612 36428
rect 38220 36370 38276 36382
rect 38220 36318 38222 36370
rect 38274 36318 38276 36370
rect 38220 36148 38276 36318
rect 38220 36082 38276 36092
rect 38220 35924 38276 35934
rect 38108 35922 38276 35924
rect 38108 35870 38222 35922
rect 38274 35870 38276 35922
rect 38108 35868 38276 35870
rect 38220 35858 38276 35868
rect 39004 35922 39060 36652
rect 39004 35870 39006 35922
rect 39058 35870 39060 35922
rect 39004 35858 39060 35870
rect 39228 36484 39284 36494
rect 39228 35922 39284 36428
rect 39228 35870 39230 35922
rect 39282 35870 39284 35922
rect 39228 35858 39284 35870
rect 37884 35698 38052 35700
rect 37884 35646 37886 35698
rect 37938 35646 38052 35698
rect 37884 35644 38052 35646
rect 38332 35810 38388 35822
rect 38332 35758 38334 35810
rect 38386 35758 38388 35810
rect 37660 34962 37716 34972
rect 37492 32508 37604 32564
rect 37660 32564 37716 32574
rect 37884 32564 37940 35644
rect 38332 35364 38388 35758
rect 38332 35298 38388 35308
rect 38556 35698 38612 35710
rect 38556 35646 38558 35698
rect 38610 35646 38612 35698
rect 38332 35140 38388 35150
rect 38556 35140 38612 35646
rect 38892 35700 38948 35710
rect 39340 35700 39396 35710
rect 38892 35698 39508 35700
rect 38892 35646 38894 35698
rect 38946 35646 39342 35698
rect 39394 35646 39508 35698
rect 38892 35644 39508 35646
rect 38892 35634 38948 35644
rect 39340 35634 39396 35644
rect 38388 35084 38612 35140
rect 38332 35074 38388 35084
rect 38220 35028 38276 35038
rect 38220 34934 38276 34972
rect 38332 34914 38388 34926
rect 38332 34862 38334 34914
rect 38386 34862 38388 34914
rect 37996 34802 38052 34814
rect 37996 34750 37998 34802
rect 38050 34750 38052 34802
rect 37996 34132 38052 34750
rect 38332 34692 38388 34862
rect 38780 34692 38836 34702
rect 38332 34690 38836 34692
rect 38332 34638 38782 34690
rect 38834 34638 38836 34690
rect 38332 34636 38836 34638
rect 37996 34066 38052 34076
rect 38332 34132 38388 34142
rect 38332 34018 38388 34076
rect 38332 33966 38334 34018
rect 38386 33966 38388 34018
rect 38332 33954 38388 33966
rect 38444 33348 38500 33358
rect 38332 33346 38500 33348
rect 38332 33294 38446 33346
rect 38498 33294 38500 33346
rect 38332 33292 38500 33294
rect 38108 33236 38164 33246
rect 38108 33142 38164 33180
rect 38108 32788 38164 32798
rect 38108 32694 38164 32732
rect 37716 32508 37940 32564
rect 37436 32498 37492 32508
rect 37660 32450 37716 32508
rect 37660 32398 37662 32450
rect 37714 32398 37716 32450
rect 37660 32386 37716 32398
rect 37268 31948 37380 32004
rect 37212 31938 37268 31948
rect 37884 31892 37940 31902
rect 37100 31838 37102 31890
rect 37154 31838 37156 31890
rect 37100 31826 37156 31838
rect 37548 31836 37884 31892
rect 35420 31780 35476 31790
rect 35420 31686 35476 31724
rect 35868 31780 35924 31790
rect 35868 31218 35924 31724
rect 37548 31778 37604 31836
rect 37884 31798 37940 31836
rect 37548 31726 37550 31778
rect 37602 31726 37604 31778
rect 37548 31714 37604 31726
rect 37996 31780 38052 31790
rect 37996 31686 38052 31724
rect 35868 31166 35870 31218
rect 35922 31166 35924 31218
rect 35868 31154 35924 31166
rect 35308 31054 35310 31106
rect 35362 31054 35364 31106
rect 35308 31042 35364 31054
rect 34860 30706 34916 30716
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34636 30158 34638 30210
rect 34690 30158 34692 30210
rect 34524 29988 34580 29998
rect 34636 29988 34692 30158
rect 37100 30210 37156 30222
rect 37100 30158 37102 30210
rect 37154 30158 37156 30210
rect 35420 30100 35476 30110
rect 34580 29932 34692 29988
rect 35084 29988 35140 29998
rect 35420 29988 35476 30044
rect 35084 29986 35476 29988
rect 35084 29934 35086 29986
rect 35138 29934 35476 29986
rect 35084 29932 35476 29934
rect 35756 29986 35812 29998
rect 35756 29934 35758 29986
rect 35810 29934 35812 29986
rect 34524 29922 34580 29932
rect 35084 29764 35140 29932
rect 35084 29698 35140 29708
rect 35644 29428 35700 29438
rect 35756 29428 35812 29934
rect 35644 29426 35812 29428
rect 35644 29374 35646 29426
rect 35698 29374 35812 29426
rect 35644 29372 35812 29374
rect 35644 29362 35700 29372
rect 35196 29036 35460 29046
rect 34524 28980 34580 28990
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34412 28420 34468 28430
rect 34188 28418 34468 28420
rect 34188 28366 34414 28418
rect 34466 28366 34468 28418
rect 34188 28364 34468 28366
rect 33852 28018 33908 28028
rect 32508 27860 32564 27870
rect 32508 27766 32564 27804
rect 33852 27188 33908 27198
rect 34412 27188 34468 28364
rect 34524 28196 34580 28924
rect 34860 28754 34916 28766
rect 34860 28702 34862 28754
rect 34914 28702 34916 28754
rect 34860 28644 34916 28702
rect 34860 28578 34916 28588
rect 35308 28642 35364 28654
rect 35308 28590 35310 28642
rect 35362 28590 35364 28642
rect 34524 28082 34580 28140
rect 34524 28030 34526 28082
rect 34578 28030 34580 28082
rect 34524 28018 34580 28030
rect 33852 27186 34468 27188
rect 33852 27134 33854 27186
rect 33906 27134 34468 27186
rect 33852 27132 34468 27134
rect 34972 27860 35028 27870
rect 34972 27746 35028 27804
rect 34972 27694 34974 27746
rect 35026 27694 35028 27746
rect 33852 27122 33908 27132
rect 34972 26908 35028 27694
rect 35308 27636 35364 28590
rect 35308 27570 35364 27580
rect 35756 27858 35812 29372
rect 36428 29652 36484 29662
rect 35980 29314 36036 29326
rect 35980 29262 35982 29314
rect 36034 29262 36036 29314
rect 35868 29204 35924 29214
rect 35980 29204 36036 29262
rect 35924 29148 36036 29204
rect 35868 28756 35924 29148
rect 35868 28642 35924 28700
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35868 28578 35924 28590
rect 36428 28754 36484 29596
rect 36988 29652 37044 29662
rect 36988 29538 37044 29596
rect 36988 29486 36990 29538
rect 37042 29486 37044 29538
rect 36988 29474 37044 29486
rect 36876 29428 36932 29438
rect 36876 29334 36932 29372
rect 36428 28702 36430 28754
rect 36482 28702 36484 28754
rect 36092 28196 36148 28206
rect 36092 28082 36148 28140
rect 36092 28030 36094 28082
rect 36146 28030 36148 28082
rect 36092 28018 36148 28030
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34412 26852 34468 26862
rect 34972 26852 35140 26908
rect 34412 26516 34468 26796
rect 33964 26514 34468 26516
rect 33964 26462 34414 26514
rect 34466 26462 34468 26514
rect 33964 26460 34468 26462
rect 33292 26404 33348 26414
rect 32396 25956 32452 25966
rect 32396 25506 32452 25900
rect 33292 25620 33348 26348
rect 33964 26402 34020 26460
rect 34412 26450 34468 26460
rect 33964 26350 33966 26402
rect 34018 26350 34020 26402
rect 33964 26338 34020 26350
rect 33852 26068 33908 26078
rect 33852 26066 34020 26068
rect 33852 26014 33854 26066
rect 33906 26014 34020 26066
rect 33852 26012 34020 26014
rect 33852 26002 33908 26012
rect 32732 25564 33348 25620
rect 32396 25454 32398 25506
rect 32450 25454 32452 25506
rect 32396 25442 32452 25454
rect 32620 25508 32676 25518
rect 32620 25394 32676 25452
rect 32732 25506 32788 25564
rect 32732 25454 32734 25506
rect 32786 25454 32788 25506
rect 32732 25442 32788 25454
rect 33292 25506 33348 25564
rect 33852 25732 33908 25742
rect 33852 25618 33908 25676
rect 33852 25566 33854 25618
rect 33906 25566 33908 25618
rect 33852 25554 33908 25566
rect 33292 25454 33294 25506
rect 33346 25454 33348 25506
rect 32620 25342 32622 25394
rect 32674 25342 32676 25394
rect 32620 25330 32676 25342
rect 32956 25396 33012 25406
rect 32956 25302 33012 25340
rect 33180 25284 33236 25294
rect 33180 25190 33236 25228
rect 32284 25106 32340 25116
rect 31388 24948 31444 24958
rect 31276 24946 31556 24948
rect 31276 24894 31390 24946
rect 31442 24894 31556 24946
rect 31276 24892 31556 24894
rect 31388 24882 31444 24892
rect 29708 24546 29764 24556
rect 31500 24162 31556 24892
rect 32956 24722 33012 24734
rect 32956 24670 32958 24722
rect 33010 24670 33012 24722
rect 31836 24610 31892 24622
rect 31836 24558 31838 24610
rect 31890 24558 31892 24610
rect 31500 24110 31502 24162
rect 31554 24110 31556 24162
rect 31500 24098 31556 24110
rect 31724 24500 31780 24510
rect 31836 24500 31892 24558
rect 31780 24444 31892 24500
rect 31612 23828 31668 23838
rect 29932 23716 29988 23726
rect 29988 23660 30100 23716
rect 29932 23650 29988 23660
rect 30044 23266 30100 23660
rect 30044 23214 30046 23266
rect 30098 23214 30100 23266
rect 30044 23202 30100 23214
rect 30716 23380 30772 23390
rect 30716 23154 30772 23324
rect 30716 23102 30718 23154
rect 30770 23102 30772 23154
rect 30716 23044 30772 23102
rect 30716 22978 30772 22988
rect 31612 22596 31668 23772
rect 31164 22540 31668 22596
rect 30156 20916 30212 20926
rect 30156 20822 30212 20860
rect 30716 20804 30772 20814
rect 30940 20804 30996 20814
rect 30716 20802 30940 20804
rect 30716 20750 30718 20802
rect 30770 20750 30940 20802
rect 30716 20748 30940 20750
rect 30716 20738 30772 20748
rect 29708 20690 29764 20702
rect 29708 20638 29710 20690
rect 29762 20638 29764 20690
rect 29708 20580 29764 20638
rect 29708 20524 30100 20580
rect 29596 20412 29876 20468
rect 29036 20122 29092 20132
rect 29148 20132 29316 20188
rect 28252 19954 28308 19964
rect 28588 20020 28644 20030
rect 29148 20020 29204 20132
rect 28588 20018 29204 20020
rect 28588 19966 28590 20018
rect 28642 19966 29204 20018
rect 28588 19964 29204 19966
rect 28588 19954 28644 19964
rect 28476 18676 28532 18686
rect 28476 18582 28532 18620
rect 29372 18676 29428 18686
rect 28700 18562 28756 18574
rect 28700 18510 28702 18562
rect 28754 18510 28756 18562
rect 28588 18452 28644 18462
rect 28588 18358 28644 18396
rect 28140 18338 28196 18350
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18228 28196 18286
rect 28700 18228 28756 18510
rect 29036 18450 29092 18462
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 28924 18340 28980 18350
rect 29036 18340 29092 18398
rect 28980 18284 29092 18340
rect 28924 18274 28980 18284
rect 28140 18172 28756 18228
rect 27916 17378 27972 17388
rect 28364 17444 28420 17454
rect 28364 17350 28420 17388
rect 28700 17220 28756 18172
rect 28700 17154 28756 17164
rect 28812 17668 28868 17678
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27692 16098 27748 16830
rect 27692 16046 27694 16098
rect 27746 16046 27748 16098
rect 27692 16034 27748 16046
rect 28028 17106 28084 17118
rect 28028 17054 28030 17106
rect 28082 17054 28084 17106
rect 27468 15988 27524 15998
rect 27468 15894 27524 15932
rect 25228 15874 25284 15886
rect 25228 15822 25230 15874
rect 25282 15822 25284 15874
rect 25228 15764 25284 15822
rect 25228 15698 25284 15708
rect 27916 15874 27972 15886
rect 27916 15822 27918 15874
rect 27970 15822 27972 15874
rect 27916 15540 27972 15822
rect 27356 15484 27972 15540
rect 27356 15426 27412 15484
rect 27356 15374 27358 15426
rect 27410 15374 27412 15426
rect 27356 15362 27412 15374
rect 26684 15314 26740 15326
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15204 26740 15262
rect 26684 15148 26964 15204
rect 26908 15092 27076 15148
rect 26796 14868 26852 14878
rect 26460 14644 26516 14654
rect 25228 12964 25284 12974
rect 25228 12740 25284 12908
rect 25228 12674 25284 12684
rect 25340 10612 25396 10622
rect 25340 10518 25396 10556
rect 25004 9874 25060 9884
rect 25340 10388 25396 10398
rect 24892 9828 24948 9838
rect 24780 9826 24948 9828
rect 24780 9774 24894 9826
rect 24946 9774 24948 9826
rect 24780 9772 24948 9774
rect 24780 7698 24836 9772
rect 24892 9762 24948 9772
rect 25340 9826 25396 10332
rect 25340 9774 25342 9826
rect 25394 9774 25396 9826
rect 25340 9762 25396 9774
rect 26460 9714 26516 14588
rect 26796 14530 26852 14812
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26796 14466 26852 14478
rect 27020 13748 27076 15092
rect 27580 14644 27636 14654
rect 27580 14550 27636 14588
rect 27132 14308 27188 14318
rect 27132 14214 27188 14252
rect 27916 13860 27972 13870
rect 28028 13860 28084 17054
rect 28140 17108 28196 17118
rect 28140 16994 28196 17052
rect 28812 17108 28868 17612
rect 28812 17052 29316 17108
rect 28140 16942 28142 16994
rect 28194 16942 28196 16994
rect 28140 16930 28196 16942
rect 28700 16996 28756 17006
rect 28812 16996 28868 17052
rect 28700 16994 28868 16996
rect 28700 16942 28702 16994
rect 28754 16942 28868 16994
rect 28700 16940 28868 16942
rect 28700 16930 28756 16940
rect 28252 16882 28308 16894
rect 28252 16830 28254 16882
rect 28306 16830 28308 16882
rect 28252 16772 28308 16830
rect 28924 16882 28980 16894
rect 28924 16830 28926 16882
rect 28978 16830 28980 16882
rect 28252 16706 28308 16716
rect 28812 16772 28868 16782
rect 28812 16678 28868 16716
rect 28140 15988 28196 15998
rect 28140 15894 28196 15932
rect 28364 15988 28420 15998
rect 28364 15894 28420 15932
rect 28476 14756 28532 14766
rect 27916 13858 28084 13860
rect 27916 13806 27918 13858
rect 27970 13806 28084 13858
rect 27916 13804 28084 13806
rect 28140 14308 28196 14318
rect 27916 13794 27972 13804
rect 27132 13748 27188 13758
rect 27020 13746 27188 13748
rect 27020 13694 27134 13746
rect 27186 13694 27188 13746
rect 27020 13692 27188 13694
rect 26684 12740 26740 12750
rect 26684 12290 26740 12684
rect 27020 12404 27076 12414
rect 26684 12238 26686 12290
rect 26738 12238 26740 12290
rect 26684 12226 26740 12238
rect 26796 12402 27076 12404
rect 26796 12350 27022 12402
rect 27074 12350 27076 12402
rect 26796 12348 27076 12350
rect 26796 11506 26852 12348
rect 27020 12338 27076 12348
rect 27020 12178 27076 12190
rect 27020 12126 27022 12178
rect 27074 12126 27076 12178
rect 27020 12068 27076 12126
rect 27020 12002 27076 12012
rect 26796 11454 26798 11506
rect 26850 11454 26852 11506
rect 26796 11442 26852 11454
rect 27132 11508 27188 13692
rect 27468 12740 27524 12750
rect 27468 12646 27524 12684
rect 27692 12292 27748 12302
rect 27580 12290 27748 12292
rect 27580 12238 27694 12290
rect 27746 12238 27748 12290
rect 27580 12236 27748 12238
rect 26684 10836 26740 10846
rect 26684 10834 27076 10836
rect 26684 10782 26686 10834
rect 26738 10782 27076 10834
rect 26684 10780 27076 10782
rect 26684 10770 26740 10780
rect 27020 10722 27076 10780
rect 27020 10670 27022 10722
rect 27074 10670 27076 10722
rect 26908 10610 26964 10622
rect 26908 10558 26910 10610
rect 26962 10558 26964 10610
rect 26684 9938 26740 9950
rect 26684 9886 26686 9938
rect 26738 9886 26740 9938
rect 26684 9828 26740 9886
rect 26460 9662 26462 9714
rect 26514 9662 26516 9714
rect 26460 9650 26516 9662
rect 26572 9772 26684 9828
rect 24780 7646 24782 7698
rect 24834 7646 24836 7698
rect 24780 7634 24836 7646
rect 25452 8484 25508 8494
rect 24332 7474 24724 7476
rect 24332 7422 24334 7474
rect 24386 7422 24724 7474
rect 24332 7420 24724 7422
rect 24332 7410 24388 7420
rect 24108 7252 24164 7262
rect 24108 7158 24164 7196
rect 24444 7028 24500 7038
rect 24332 6804 24388 6814
rect 24332 6710 24388 6748
rect 24444 6690 24500 6972
rect 24444 6638 24446 6690
rect 24498 6638 24500 6690
rect 23996 6130 24052 6300
rect 24108 6580 24164 6590
rect 24108 6244 24164 6524
rect 24108 6178 24164 6188
rect 24444 6580 24500 6638
rect 25116 6692 25172 6702
rect 24780 6580 24836 6590
rect 24444 6578 24836 6580
rect 24444 6526 24782 6578
rect 24834 6526 24836 6578
rect 24444 6524 24836 6526
rect 23996 6078 23998 6130
rect 24050 6078 24052 6130
rect 23996 6066 24052 6078
rect 23324 5964 23604 6020
rect 23548 5906 23604 5964
rect 23548 5854 23550 5906
rect 23602 5854 23604 5906
rect 23548 5842 23604 5854
rect 23212 5182 23214 5234
rect 23266 5182 23268 5234
rect 23212 5170 23268 5182
rect 23100 4900 23156 4910
rect 22428 4898 23156 4900
rect 22428 4846 23102 4898
rect 23154 4846 23156 4898
rect 22428 4844 23156 4846
rect 22428 4450 22484 4844
rect 23100 4834 23156 4844
rect 22428 4398 22430 4450
rect 22482 4398 22484 4450
rect 22428 4386 22484 4398
rect 21644 4286 21646 4338
rect 21698 4286 21700 4338
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 21644 3666 21700 4286
rect 24444 4228 24500 6524
rect 24780 6514 24836 6524
rect 25004 6580 25060 6590
rect 25004 6486 25060 6524
rect 25116 6466 25172 6636
rect 25452 6690 25508 8428
rect 26572 8484 26628 9772
rect 26684 9762 26740 9772
rect 26348 7476 26404 7486
rect 26348 7382 26404 7420
rect 26572 7474 26628 8428
rect 26908 9604 26964 10558
rect 27020 10276 27076 10670
rect 27132 10612 27188 11452
rect 27244 12178 27300 12190
rect 27244 12126 27246 12178
rect 27298 12126 27300 12178
rect 27244 10834 27300 12126
rect 27468 12178 27524 12190
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27468 12068 27524 12126
rect 27468 12002 27524 12012
rect 27468 11508 27524 11518
rect 27468 11394 27524 11452
rect 27468 11342 27470 11394
rect 27522 11342 27524 11394
rect 27468 11330 27524 11342
rect 27244 10782 27246 10834
rect 27298 10782 27300 10834
rect 27244 10770 27300 10782
rect 27132 10546 27188 10556
rect 27020 10210 27076 10220
rect 27468 10498 27524 10510
rect 27468 10446 27470 10498
rect 27522 10446 27524 10498
rect 27468 9940 27524 10446
rect 27468 9874 27524 9884
rect 27580 10164 27636 12236
rect 27692 12226 27748 12236
rect 27804 12178 27860 12190
rect 27804 12126 27806 12178
rect 27858 12126 27860 12178
rect 27804 12068 27860 12126
rect 27804 12002 27860 12012
rect 28140 11620 28196 14252
rect 28476 13076 28532 14700
rect 28924 13860 28980 16830
rect 29260 16098 29316 17052
rect 29372 16884 29428 18620
rect 29708 17444 29764 17454
rect 29708 16884 29764 17388
rect 29820 16996 29876 20412
rect 30044 19346 30100 20524
rect 30044 19294 30046 19346
rect 30098 19294 30100 19346
rect 30044 19282 30100 19294
rect 30492 20020 30548 20030
rect 29932 19010 29988 19022
rect 29932 18958 29934 19010
rect 29986 18958 29988 19010
rect 29932 18788 29988 18958
rect 30156 19012 30212 19022
rect 30268 19012 30324 19022
rect 30156 19010 30268 19012
rect 30156 18958 30158 19010
rect 30210 18958 30268 19010
rect 30156 18956 30268 18958
rect 30156 18946 30212 18956
rect 29932 18722 29988 18732
rect 29820 16940 30212 16996
rect 29372 16882 29652 16884
rect 29372 16830 29374 16882
rect 29426 16830 29652 16882
rect 29372 16828 29652 16830
rect 29372 16818 29428 16828
rect 29260 16046 29262 16098
rect 29314 16046 29316 16098
rect 29260 16034 29316 16046
rect 29372 15988 29428 15998
rect 29596 15988 29652 16828
rect 29708 16882 29876 16884
rect 29708 16830 29710 16882
rect 29762 16830 29876 16882
rect 29708 16828 29876 16830
rect 29708 16818 29764 16828
rect 29708 15988 29764 15998
rect 29596 15986 29764 15988
rect 29596 15934 29710 15986
rect 29762 15934 29764 15986
rect 29596 15932 29764 15934
rect 29372 15894 29428 15932
rect 29708 15922 29764 15932
rect 29484 15874 29540 15886
rect 29484 15822 29486 15874
rect 29538 15822 29540 15874
rect 29484 15202 29540 15822
rect 29484 15150 29486 15202
rect 29538 15150 29540 15202
rect 29484 15148 29540 15150
rect 29820 15204 29876 16828
rect 29932 15204 29988 15214
rect 29820 15202 29988 15204
rect 29820 15150 29934 15202
rect 29986 15150 29988 15202
rect 29820 15148 29988 15150
rect 29484 15092 29652 15148
rect 28924 13794 28980 13804
rect 28476 13010 28532 13020
rect 29484 12964 29540 12974
rect 28252 12068 28308 12078
rect 28252 11974 28308 12012
rect 28252 11620 28308 11630
rect 28140 11564 28252 11620
rect 28252 11394 28308 11564
rect 29260 11508 29316 11518
rect 29484 11508 29540 12908
rect 29316 11452 29540 11508
rect 29260 11414 29316 11452
rect 28252 11342 28254 11394
rect 28306 11342 28308 11394
rect 28252 11330 28308 11342
rect 29596 11284 29652 15092
rect 29932 13636 29988 15148
rect 29932 12964 29988 13580
rect 30044 13860 30100 13870
rect 30044 13634 30100 13804
rect 30044 13582 30046 13634
rect 30098 13582 30100 13634
rect 30044 13570 30100 13582
rect 29932 12898 29988 12908
rect 30156 12180 30212 16940
rect 30268 16324 30324 18956
rect 30380 19010 30436 19022
rect 30380 18958 30382 19010
rect 30434 18958 30436 19010
rect 30380 18676 30436 18958
rect 30380 18610 30436 18620
rect 30492 17668 30548 19964
rect 30716 19906 30772 19918
rect 30716 19854 30718 19906
rect 30770 19854 30772 19906
rect 30716 19012 30772 19854
rect 30940 19012 30996 20748
rect 31052 20020 31108 20030
rect 31052 19926 31108 19964
rect 30716 18946 30772 18956
rect 30828 19010 30996 19012
rect 30828 18958 30942 19010
rect 30994 18958 30996 19010
rect 30828 18956 30996 18958
rect 30492 17574 30548 17612
rect 30716 17442 30772 17454
rect 30716 17390 30718 17442
rect 30770 17390 30772 17442
rect 30716 17108 30772 17390
rect 30828 17444 30884 18956
rect 30940 18946 30996 18956
rect 31164 17892 31220 22540
rect 31388 20690 31444 20702
rect 31388 20638 31390 20690
rect 31442 20638 31444 20690
rect 31276 20244 31332 20254
rect 31388 20244 31444 20638
rect 31276 20242 31444 20244
rect 31276 20190 31278 20242
rect 31330 20190 31444 20242
rect 31276 20188 31444 20190
rect 31276 20178 31332 20188
rect 31612 20132 31668 20142
rect 31612 20038 31668 20076
rect 31388 20020 31444 20030
rect 31388 19926 31444 19964
rect 31724 19796 31780 24444
rect 32060 23828 32116 23838
rect 32060 23734 32116 23772
rect 31948 23492 32004 23502
rect 31948 21700 32004 23436
rect 31948 20244 32004 21644
rect 31836 20188 32004 20244
rect 32956 20188 33012 24670
rect 33292 24722 33348 25454
rect 33516 25508 33572 25518
rect 33516 25060 33572 25452
rect 33628 25284 33684 25294
rect 33684 25228 33796 25284
rect 33628 25218 33684 25228
rect 33516 25004 33684 25060
rect 33292 24670 33294 24722
rect 33346 24670 33348 24722
rect 33292 24658 33348 24670
rect 33628 24722 33684 25004
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 33740 23938 33796 25228
rect 33740 23886 33742 23938
rect 33794 23886 33796 23938
rect 33740 23874 33796 23886
rect 33404 23714 33460 23726
rect 33404 23662 33406 23714
rect 33458 23662 33460 23714
rect 33404 23492 33460 23662
rect 33404 23426 33460 23436
rect 33628 23380 33684 23390
rect 33964 23380 34020 26012
rect 34188 25732 34244 25742
rect 34188 25618 34244 25676
rect 34188 25566 34190 25618
rect 34242 25566 34244 25618
rect 34188 25554 34244 25566
rect 34972 25732 35028 25742
rect 34636 25508 34692 25518
rect 34636 25394 34692 25452
rect 34972 25506 35028 25676
rect 34972 25454 34974 25506
rect 35026 25454 35028 25506
rect 34972 25442 35028 25454
rect 34636 25342 34638 25394
rect 34690 25342 34692 25394
rect 34636 25330 34692 25342
rect 34076 25284 34132 25294
rect 34076 25190 34132 25228
rect 34188 24836 34244 24846
rect 34188 24722 34244 24780
rect 34188 24670 34190 24722
rect 34242 24670 34244 24722
rect 34188 24658 34244 24670
rect 34076 23380 34132 23390
rect 33628 23378 34132 23380
rect 33628 23326 33630 23378
rect 33682 23326 34078 23378
rect 34130 23326 34132 23378
rect 33628 23324 34132 23326
rect 31836 20020 31892 20188
rect 32060 20132 32116 20142
rect 32396 20132 32452 20142
rect 32060 20038 32116 20076
rect 32284 20130 32452 20132
rect 32284 20078 32398 20130
rect 32450 20078 32452 20130
rect 32284 20076 32452 20078
rect 31836 19954 31892 19964
rect 31948 20018 32004 20030
rect 31948 19966 31950 20018
rect 32002 19966 32004 20018
rect 31724 19740 31892 19796
rect 31500 19124 31556 19134
rect 31052 17836 31220 17892
rect 31388 18340 31444 18350
rect 30940 17780 30996 17790
rect 30940 17666 30996 17724
rect 30940 17614 30942 17666
rect 30994 17614 30996 17666
rect 30940 17602 30996 17614
rect 30828 17378 30884 17388
rect 30380 17052 30772 17108
rect 30380 16994 30436 17052
rect 30380 16942 30382 16994
rect 30434 16942 30436 16994
rect 30380 16930 30436 16942
rect 31052 16436 31108 17836
rect 31388 17780 31444 18284
rect 31388 17714 31444 17724
rect 31164 17668 31220 17678
rect 31164 17574 31220 17612
rect 31500 17666 31556 19068
rect 31500 17614 31502 17666
rect 31554 17614 31556 17666
rect 31500 17602 31556 17614
rect 31612 17668 31668 17678
rect 31612 17574 31668 17612
rect 31724 17442 31780 17454
rect 31724 17390 31726 17442
rect 31778 17390 31780 17442
rect 31500 17220 31556 17230
rect 31052 16380 31220 16436
rect 30268 16268 31108 16324
rect 30492 13636 30548 13646
rect 30492 13542 30548 13580
rect 30156 12086 30212 12124
rect 30268 12850 30324 12862
rect 30268 12798 30270 12850
rect 30322 12798 30324 12850
rect 30268 11844 30324 12798
rect 30940 12066 30996 12078
rect 30940 12014 30942 12066
rect 30994 12014 30996 12066
rect 30604 11844 30660 11854
rect 30268 11788 30604 11844
rect 30604 11778 30660 11788
rect 29708 11620 29764 11630
rect 29708 11506 29764 11564
rect 29708 11454 29710 11506
rect 29762 11454 29764 11506
rect 29708 11442 29764 11454
rect 30156 11508 30212 11518
rect 29596 11228 29764 11284
rect 27580 9826 27636 10108
rect 27580 9774 27582 9826
rect 27634 9774 27636 9826
rect 27580 9762 27636 9774
rect 27916 11170 27972 11182
rect 27916 11118 27918 11170
rect 27970 11118 27972 11170
rect 27580 9604 27636 9614
rect 26908 9602 27636 9604
rect 26908 9550 27582 9602
rect 27634 9550 27636 9602
rect 26908 9548 27636 9550
rect 26908 8258 26964 9548
rect 27580 9538 27636 9548
rect 26908 8206 26910 8258
rect 26962 8206 26964 8258
rect 26572 7422 26574 7474
rect 26626 7422 26628 7474
rect 26572 7410 26628 7422
rect 26684 8034 26740 8046
rect 26684 7982 26686 8034
rect 26738 7982 26740 8034
rect 26684 7588 26740 7982
rect 26796 8034 26852 8046
rect 26796 7982 26798 8034
rect 26850 7982 26852 8034
rect 26796 7812 26852 7982
rect 26908 8036 26964 8206
rect 27356 8260 27412 8270
rect 27356 8166 27412 8204
rect 27916 8148 27972 11118
rect 29596 10498 29652 10510
rect 29596 10446 29598 10498
rect 29650 10446 29652 10498
rect 29596 9940 29652 10446
rect 29596 9874 29652 9884
rect 28028 9828 28084 9838
rect 28028 9734 28084 9772
rect 28588 9716 28644 9726
rect 28588 9622 28644 9660
rect 29708 9492 29764 11228
rect 30156 11172 30212 11452
rect 30604 11172 30660 11182
rect 30940 11172 30996 12014
rect 30156 11170 30996 11172
rect 30156 11118 30606 11170
rect 30658 11118 30996 11170
rect 30156 11116 30996 11118
rect 30156 10612 30212 11116
rect 30604 11106 30660 11116
rect 30268 10612 30324 10622
rect 30940 10612 30996 10622
rect 30156 10610 30324 10612
rect 30156 10558 30270 10610
rect 30322 10558 30324 10610
rect 30156 10556 30324 10558
rect 29932 9716 29988 9726
rect 29932 9622 29988 9660
rect 30044 9604 30100 9614
rect 30044 9510 30100 9548
rect 29708 9426 29764 9436
rect 28028 8148 28084 8158
rect 27916 8092 28028 8148
rect 26908 7970 26964 7980
rect 26796 7756 26964 7812
rect 26796 7588 26852 7598
rect 26684 7586 26852 7588
rect 26684 7534 26798 7586
rect 26850 7534 26852 7586
rect 26684 7532 26852 7534
rect 25788 7364 25844 7374
rect 25788 7270 25844 7308
rect 25452 6638 25454 6690
rect 25506 6638 25508 6690
rect 25452 6626 25508 6638
rect 25900 7252 25956 7262
rect 25900 6916 25956 7196
rect 26124 7252 26180 7262
rect 26684 7252 26740 7532
rect 26796 7522 26852 7532
rect 26124 7250 26740 7252
rect 26124 7198 26126 7250
rect 26178 7198 26740 7250
rect 26124 7196 26740 7198
rect 26796 7364 26852 7374
rect 26124 7186 26180 7196
rect 25900 6690 25956 6860
rect 26796 6914 26852 7308
rect 26796 6862 26798 6914
rect 26850 6862 26852 6914
rect 26796 6850 26852 6862
rect 26908 6914 26964 7756
rect 27020 7474 27076 7486
rect 27020 7422 27022 7474
rect 27074 7422 27076 7474
rect 27020 7364 27076 7422
rect 27020 7298 27076 7308
rect 27244 7476 27300 7486
rect 26908 6862 26910 6914
rect 26962 6862 26964 6914
rect 26908 6850 26964 6862
rect 27244 6916 27300 7420
rect 27692 7364 27748 7374
rect 27692 7270 27748 7308
rect 27244 6850 27300 6860
rect 25900 6638 25902 6690
rect 25954 6638 25956 6690
rect 25900 6626 25956 6638
rect 26236 6692 26292 6702
rect 26236 6578 26292 6636
rect 26236 6526 26238 6578
rect 26290 6526 26292 6578
rect 25116 6414 25118 6466
rect 25170 6414 25172 6466
rect 25116 6402 25172 6414
rect 26124 6466 26180 6478
rect 26124 6414 26126 6466
rect 26178 6414 26180 6466
rect 26124 5234 26180 6414
rect 26236 6244 26292 6526
rect 27244 6692 27300 6702
rect 27244 6578 27300 6636
rect 27580 6692 27636 6702
rect 28028 6692 28084 8092
rect 29820 8036 29876 8046
rect 29820 7586 29876 7980
rect 30268 7812 30324 10556
rect 30716 10610 30996 10612
rect 30716 10558 30942 10610
rect 30994 10558 30996 10610
rect 30716 10556 30996 10558
rect 30492 9940 30548 9950
rect 30492 9846 30548 9884
rect 30716 9714 30772 10556
rect 30940 10546 30996 10556
rect 30716 9662 30718 9714
rect 30770 9662 30772 9714
rect 30716 9650 30772 9662
rect 31052 9716 31108 16268
rect 31164 10948 31220 16380
rect 31500 15314 31556 17164
rect 31724 16324 31780 17390
rect 31724 16258 31780 16268
rect 31724 15876 31780 15886
rect 31836 15876 31892 19740
rect 31948 19124 32004 19966
rect 31948 19058 32004 19068
rect 32172 20018 32228 20030
rect 32172 19966 32174 20018
rect 32226 19966 32228 20018
rect 31780 15820 31892 15876
rect 31948 18788 32004 18798
rect 31724 15810 31780 15820
rect 31500 15262 31502 15314
rect 31554 15262 31556 15314
rect 31500 15250 31556 15262
rect 31724 15204 31780 15214
rect 31724 15110 31780 15148
rect 31948 13860 32004 18732
rect 32172 18452 32228 19966
rect 32172 18386 32228 18396
rect 32284 18228 32340 20076
rect 32396 20066 32452 20076
rect 32620 20132 33012 20188
rect 33068 23042 33124 23054
rect 33068 22990 33070 23042
rect 33122 22990 33124 23042
rect 32172 17668 32228 17678
rect 32284 17668 32340 18172
rect 32172 17666 32340 17668
rect 32172 17614 32174 17666
rect 32226 17614 32340 17666
rect 32172 17612 32340 17614
rect 32172 17602 32228 17612
rect 32508 16772 32564 16782
rect 32508 16678 32564 16716
rect 32172 16212 32228 16222
rect 32172 16118 32228 16156
rect 32508 16098 32564 16110
rect 32508 16046 32510 16098
rect 32562 16046 32564 16098
rect 32508 15204 32564 16046
rect 32508 15138 32564 15148
rect 32060 15092 32116 15102
rect 32060 14998 32116 15036
rect 31724 13804 32004 13860
rect 31612 12628 31668 12638
rect 31500 11844 31556 11854
rect 31500 11170 31556 11788
rect 31612 11394 31668 12572
rect 31612 11342 31614 11394
rect 31666 11342 31668 11394
rect 31612 11330 31668 11342
rect 31724 11172 31780 13804
rect 32172 13748 32228 13758
rect 31836 13636 31892 13646
rect 32060 13636 32116 13646
rect 31892 13634 32116 13636
rect 31892 13582 32062 13634
rect 32114 13582 32116 13634
rect 31892 13580 32116 13582
rect 31836 13570 31892 13580
rect 32060 13570 32116 13580
rect 32060 12964 32116 12974
rect 32060 11956 32116 12908
rect 32172 12852 32228 13692
rect 32172 12786 32228 12796
rect 32396 13634 32452 13646
rect 32396 13582 32398 13634
rect 32450 13582 32452 13634
rect 32396 13074 32452 13582
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 32396 12852 32452 13022
rect 32396 12786 32452 12796
rect 32508 13522 32564 13534
rect 32508 13470 32510 13522
rect 32562 13470 32564 13522
rect 32508 12628 32564 13470
rect 32620 12964 32676 20132
rect 33068 18788 33124 22990
rect 33180 23044 33236 23054
rect 33180 22484 33236 22988
rect 33628 22708 33684 23324
rect 34076 23314 34132 23324
rect 33852 22932 33908 22942
rect 33628 22642 33684 22652
rect 33740 22876 33852 22932
rect 33180 22482 33572 22484
rect 33180 22430 33182 22482
rect 33234 22430 33572 22482
rect 33180 22428 33572 22430
rect 33180 22418 33236 22428
rect 33516 22370 33572 22428
rect 33516 22318 33518 22370
rect 33570 22318 33572 22370
rect 33516 22306 33572 22318
rect 33740 22148 33796 22876
rect 33852 22866 33908 22876
rect 35084 22932 35140 26852
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 25620 35476 25630
rect 35420 25396 35476 25564
rect 35420 25302 35476 25340
rect 35756 25282 35812 27806
rect 36204 25732 36260 25742
rect 36204 25618 36260 25676
rect 36204 25566 36206 25618
rect 36258 25566 36260 25618
rect 36204 25554 36260 25566
rect 36428 25396 36484 28702
rect 36988 28756 37044 28766
rect 36988 28420 37044 28700
rect 37100 28644 37156 30158
rect 37772 30100 37828 30110
rect 37212 30098 37828 30100
rect 37212 30046 37774 30098
rect 37826 30046 37828 30098
rect 37212 30044 37828 30046
rect 37212 29650 37268 30044
rect 37772 30034 37828 30044
rect 37212 29598 37214 29650
rect 37266 29598 37268 29650
rect 37212 29586 37268 29598
rect 37772 29876 37828 29886
rect 37436 29426 37492 29438
rect 37436 29374 37438 29426
rect 37490 29374 37492 29426
rect 37100 28578 37156 28588
rect 37324 28642 37380 28654
rect 37324 28590 37326 28642
rect 37378 28590 37380 28642
rect 37100 28420 37156 28430
rect 36988 28418 37156 28420
rect 36988 28366 37102 28418
rect 37154 28366 37156 28418
rect 36988 28364 37156 28366
rect 37100 28354 37156 28364
rect 37100 28196 37156 28206
rect 37324 28196 37380 28590
rect 37156 28140 37380 28196
rect 37436 28196 37492 29374
rect 37772 28530 37828 29820
rect 37884 29428 37940 29438
rect 37884 28754 37940 29372
rect 37884 28702 37886 28754
rect 37938 28702 37940 28754
rect 37884 28690 37940 28702
rect 37772 28478 37774 28530
rect 37826 28478 37828 28530
rect 37772 28466 37828 28478
rect 37100 28130 37156 28140
rect 37436 26908 37492 28140
rect 37996 28418 38052 28430
rect 37996 28366 37998 28418
rect 38050 28366 38052 28418
rect 37772 27746 37828 27758
rect 37772 27694 37774 27746
rect 37826 27694 37828 27746
rect 37772 27636 37828 27694
rect 37772 27570 37828 27580
rect 36988 26852 37492 26908
rect 37996 27074 38052 28366
rect 37996 27022 37998 27074
rect 38050 27022 38052 27074
rect 36204 25340 36484 25396
rect 36764 26178 36820 26190
rect 36764 26126 36766 26178
rect 36818 26126 36820 26178
rect 35756 25230 35758 25282
rect 35810 25230 35812 25282
rect 35420 24724 35476 24734
rect 35420 24630 35476 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35756 23938 35812 25230
rect 36092 25284 36148 25294
rect 36092 24834 36148 25228
rect 36092 24782 36094 24834
rect 36146 24782 36148 24834
rect 36092 24770 36148 24782
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35756 23874 35812 23886
rect 35980 24612 36036 24622
rect 35980 23826 36036 24556
rect 35980 23774 35982 23826
rect 36034 23774 36036 23826
rect 35980 23762 36036 23774
rect 35084 22866 35140 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22484 35588 22494
rect 34300 22260 34356 22270
rect 34300 22258 34468 22260
rect 34300 22206 34302 22258
rect 34354 22206 34468 22258
rect 34300 22204 34468 22206
rect 34300 22194 34356 22204
rect 33068 18722 33124 18732
rect 33292 22092 33796 22148
rect 33180 17444 33236 17454
rect 33180 17106 33236 17388
rect 33180 17054 33182 17106
rect 33234 17054 33236 17106
rect 33180 17042 33236 17054
rect 32732 16098 32788 16110
rect 32732 16046 32734 16098
rect 32786 16046 32788 16098
rect 32732 15876 32788 16046
rect 32732 14644 32788 15820
rect 33180 15876 33236 15886
rect 33180 15782 33236 15820
rect 32732 14578 32788 14588
rect 33068 13748 33124 13786
rect 33068 13682 33124 13692
rect 33068 13524 33124 13534
rect 32620 12898 32676 12908
rect 32732 13522 33124 13524
rect 32732 13470 33070 13522
rect 33122 13470 33124 13522
rect 32732 13468 33124 13470
rect 32508 12562 32564 12572
rect 32732 12180 32788 13468
rect 33068 13458 33124 13468
rect 33292 13300 33348 22092
rect 33628 21812 33684 21822
rect 33628 21718 33684 21756
rect 34412 21810 34468 22204
rect 34412 21758 34414 21810
rect 34466 21758 34468 21810
rect 34412 21746 34468 21758
rect 35532 21810 35588 22428
rect 35532 21758 35534 21810
rect 35586 21758 35588 21810
rect 35532 21746 35588 21758
rect 33964 21698 34020 21710
rect 33964 21646 33966 21698
rect 34018 21646 34020 21698
rect 33964 21588 34020 21646
rect 34524 21700 34580 21710
rect 34188 21588 34244 21598
rect 33964 21586 34244 21588
rect 33964 21534 34190 21586
rect 34242 21534 34244 21586
rect 33964 21532 34244 21534
rect 33516 20914 33572 20926
rect 33516 20862 33518 20914
rect 33570 20862 33572 20914
rect 33516 18452 33572 20862
rect 33964 20804 34020 20814
rect 33964 20710 34020 20748
rect 33740 19460 33796 19470
rect 33740 19236 33796 19404
rect 34188 19460 34244 21532
rect 34524 21586 34580 21644
rect 36092 21698 36148 21710
rect 36092 21646 36094 21698
rect 36146 21646 36148 21698
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34524 21522 34580 21534
rect 34860 21588 34916 21598
rect 34860 21494 34916 21532
rect 35084 21586 35140 21598
rect 35084 21534 35086 21586
rect 35138 21534 35140 21586
rect 34188 19394 34244 19404
rect 34524 19348 34580 19358
rect 34300 19236 34356 19246
rect 34524 19236 34580 19292
rect 33740 19234 34244 19236
rect 33740 19182 33742 19234
rect 33794 19182 34244 19234
rect 33740 19180 34244 19182
rect 33740 19170 33796 19180
rect 34188 19124 34244 19180
rect 34300 19234 34580 19236
rect 34300 19182 34302 19234
rect 34354 19182 34580 19234
rect 34300 19180 34580 19182
rect 34300 19170 34356 19180
rect 33516 18228 33572 18396
rect 33628 19012 33684 19022
rect 33628 18564 33684 18956
rect 33852 18676 33908 18686
rect 33852 18582 33908 18620
rect 33628 18450 33684 18508
rect 33628 18398 33630 18450
rect 33682 18398 33684 18450
rect 33628 18386 33684 18398
rect 34188 18450 34244 19068
rect 34188 18398 34190 18450
rect 34242 18398 34244 18450
rect 34188 18386 34244 18398
rect 33516 18172 33796 18228
rect 33628 16770 33684 16782
rect 33628 16718 33630 16770
rect 33682 16718 33684 16770
rect 33628 16212 33684 16718
rect 33628 16098 33684 16156
rect 33628 16046 33630 16098
rect 33682 16046 33684 16098
rect 33628 16034 33684 16046
rect 33740 16100 33796 18172
rect 34188 16772 34244 16782
rect 33964 16100 34020 16110
rect 33740 16098 34020 16100
rect 33740 16046 33966 16098
rect 34018 16046 34020 16098
rect 33740 16044 34020 16046
rect 33964 16034 34020 16044
rect 33964 15874 34020 15886
rect 33964 15822 33966 15874
rect 34018 15822 34020 15874
rect 33852 15204 33908 15214
rect 33404 15092 33460 15102
rect 33460 15036 33572 15092
rect 33404 15026 33460 15036
rect 33404 13522 33460 13534
rect 33404 13470 33406 13522
rect 33458 13470 33460 13522
rect 33404 13412 33460 13470
rect 33404 13346 33460 13356
rect 31948 11900 32116 11956
rect 32284 12124 32788 12180
rect 32844 13244 33348 13300
rect 31948 11788 32004 11900
rect 31836 11732 31892 11742
rect 31948 11732 32228 11788
rect 31836 11506 31892 11676
rect 31836 11454 31838 11506
rect 31890 11454 31892 11506
rect 31836 11442 31892 11454
rect 32060 11394 32116 11406
rect 32060 11342 32062 11394
rect 32114 11342 32116 11394
rect 32060 11284 32116 11342
rect 32060 11218 32116 11228
rect 31500 11118 31502 11170
rect 31554 11118 31556 11170
rect 31500 11106 31556 11118
rect 31612 11116 31780 11172
rect 31164 10834 31220 10892
rect 31164 10782 31166 10834
rect 31218 10782 31220 10834
rect 31164 10770 31220 10782
rect 31276 10612 31332 10622
rect 31276 10610 31556 10612
rect 31276 10558 31278 10610
rect 31330 10558 31556 10610
rect 31276 10556 31556 10558
rect 31276 10546 31332 10556
rect 31164 9940 31220 9950
rect 31164 9826 31220 9884
rect 31164 9774 31166 9826
rect 31218 9774 31220 9826
rect 31164 9762 31220 9774
rect 31388 9828 31444 9838
rect 31052 9650 31108 9660
rect 30380 9602 30436 9614
rect 30380 9550 30382 9602
rect 30434 9550 30436 9602
rect 30380 8596 30436 9550
rect 30604 9604 30660 9614
rect 30604 9510 30660 9548
rect 31388 9266 31444 9772
rect 31388 9214 31390 9266
rect 31442 9214 31444 9266
rect 31388 9202 31444 9214
rect 31500 9714 31556 10556
rect 31500 9662 31502 9714
rect 31554 9662 31556 9714
rect 31052 9154 31108 9166
rect 31052 9102 31054 9154
rect 31106 9102 31108 9154
rect 31052 8596 31108 9102
rect 30380 8540 31108 8596
rect 30604 8146 30660 8540
rect 30604 8094 30606 8146
rect 30658 8094 30660 8146
rect 30268 7756 30548 7812
rect 29820 7534 29822 7586
rect 29874 7534 29876 7586
rect 29820 7522 29876 7534
rect 27580 6690 28084 6692
rect 27580 6638 27582 6690
rect 27634 6638 28030 6690
rect 28082 6638 28084 6690
rect 27580 6636 28084 6638
rect 27580 6626 27636 6636
rect 28028 6626 28084 6636
rect 28140 7476 28196 7486
rect 27244 6526 27246 6578
rect 27298 6526 27300 6578
rect 27244 6514 27300 6526
rect 26460 6468 26516 6478
rect 26460 6374 26516 6412
rect 27692 6468 27748 6478
rect 26236 6178 26292 6188
rect 27580 5796 27636 5806
rect 27692 5796 27748 6412
rect 27580 5794 27748 5796
rect 27580 5742 27582 5794
rect 27634 5742 27748 5794
rect 27580 5740 27748 5742
rect 27580 5730 27636 5740
rect 26124 5182 26126 5234
rect 26178 5182 26180 5234
rect 26124 5170 26180 5182
rect 26012 4898 26068 4910
rect 26012 4846 26014 4898
rect 26066 4846 26068 4898
rect 26012 4450 26068 4846
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 25340 4340 25396 4350
rect 25340 4246 25396 4284
rect 24556 4228 24612 4238
rect 24444 4226 24612 4228
rect 24444 4174 24558 4226
rect 24610 4174 24612 4226
rect 24444 4172 24612 4174
rect 24556 4162 24612 4172
rect 28140 4226 28196 7420
rect 30492 7474 30548 7756
rect 30492 7422 30494 7474
rect 30546 7422 30548 7474
rect 30492 6692 30548 7422
rect 30380 6636 30492 6692
rect 29372 6580 29428 6590
rect 29372 5908 29428 6524
rect 30156 6466 30212 6478
rect 30156 6414 30158 6466
rect 30210 6414 30212 6466
rect 30156 6244 30212 6414
rect 30156 6178 30212 6188
rect 28588 4564 28644 4574
rect 28588 4470 28644 4508
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 28140 4162 28196 4174
rect 29372 4226 29428 5852
rect 30380 5906 30436 6636
rect 30492 6626 30548 6636
rect 30492 6466 30548 6478
rect 30492 6414 30494 6466
rect 30546 6414 30548 6466
rect 30492 6244 30548 6414
rect 30492 6178 30548 6188
rect 30380 5854 30382 5906
rect 30434 5854 30436 5906
rect 29708 5794 29764 5806
rect 29708 5742 29710 5794
rect 29762 5742 29764 5794
rect 29708 5348 29764 5742
rect 29708 5282 29764 5292
rect 30380 4564 30436 5854
rect 30604 5796 30660 8094
rect 30940 8372 30996 8382
rect 30940 8258 30996 8316
rect 30940 8206 30942 8258
rect 30994 8206 30996 8258
rect 30716 8036 30772 8046
rect 30716 7942 30772 7980
rect 30940 7700 30996 8206
rect 31500 8258 31556 9662
rect 31500 8206 31502 8258
rect 31554 8206 31556 8258
rect 31164 8146 31220 8158
rect 31164 8094 31166 8146
rect 31218 8094 31220 8146
rect 31164 8036 31220 8094
rect 31164 7970 31220 7980
rect 31500 7924 31556 8206
rect 31612 8260 31668 11116
rect 31724 10948 31780 10958
rect 31724 10834 31780 10892
rect 31724 10782 31726 10834
rect 31778 10782 31780 10834
rect 31724 10770 31780 10782
rect 31836 9828 31892 9838
rect 31836 9734 31892 9772
rect 32172 9828 32228 11732
rect 32284 11394 32340 12124
rect 32732 11618 32788 11630
rect 32732 11566 32734 11618
rect 32786 11566 32788 11618
rect 32284 11342 32286 11394
rect 32338 11342 32340 11394
rect 32284 11330 32340 11342
rect 32620 11396 32676 11406
rect 32732 11396 32788 11566
rect 32620 11394 32788 11396
rect 32620 11342 32622 11394
rect 32674 11342 32788 11394
rect 32620 11340 32788 11342
rect 32620 11330 32676 11340
rect 32844 11172 32900 13244
rect 33516 13188 33572 15036
rect 33740 14308 33796 14318
rect 33740 13748 33796 14252
rect 33740 13682 33796 13692
rect 33852 13746 33908 15148
rect 33964 15202 34020 15822
rect 34188 15764 34244 16716
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 34188 15708 34356 15764
rect 33964 15150 33966 15202
rect 34018 15150 34020 15202
rect 33964 15138 34020 15150
rect 34076 15314 34132 15326
rect 34076 15262 34078 15314
rect 34130 15262 34132 15314
rect 33852 13694 33854 13746
rect 33906 13694 33908 13746
rect 33068 13132 33684 13188
rect 32956 12964 33012 12974
rect 32956 12180 33012 12908
rect 33068 12402 33124 13132
rect 33628 13074 33684 13132
rect 33628 13022 33630 13074
rect 33682 13022 33684 13074
rect 33628 13010 33684 13022
rect 33068 12350 33070 12402
rect 33122 12350 33124 12402
rect 33068 12338 33124 12350
rect 33292 12962 33348 12974
rect 33292 12910 33294 12962
rect 33346 12910 33348 12962
rect 33292 12852 33348 12910
rect 32956 11508 33012 12124
rect 33292 12178 33348 12796
rect 33516 12962 33572 12974
rect 33516 12910 33518 12962
rect 33570 12910 33572 12962
rect 33516 12404 33572 12910
rect 33516 12402 33684 12404
rect 33516 12350 33518 12402
rect 33570 12350 33684 12402
rect 33516 12348 33684 12350
rect 33516 12338 33572 12348
rect 33292 12126 33294 12178
rect 33346 12126 33348 12178
rect 33180 12066 33236 12078
rect 33180 12014 33182 12066
rect 33234 12014 33236 12066
rect 33180 11618 33236 12014
rect 33180 11566 33182 11618
rect 33234 11566 33236 11618
rect 33180 11554 33236 11566
rect 33068 11508 33124 11518
rect 32956 11506 33124 11508
rect 32956 11454 33070 11506
rect 33122 11454 33124 11506
rect 32956 11452 33124 11454
rect 33068 11442 33124 11452
rect 32284 11116 32900 11172
rect 32284 9940 32340 11116
rect 33292 11060 33348 12126
rect 33516 11732 33572 11742
rect 33516 11506 33572 11676
rect 33516 11454 33518 11506
rect 33570 11454 33572 11506
rect 33516 11396 33572 11454
rect 33516 11330 33572 11340
rect 33292 10994 33348 11004
rect 32284 9846 32340 9884
rect 32844 10052 32900 10062
rect 33628 10052 33684 12348
rect 33852 10164 33908 13694
rect 34076 13412 34132 15262
rect 34188 13972 34244 13982
rect 34188 13878 34244 13916
rect 34300 13858 34356 15708
rect 34524 15148 34580 19180
rect 34636 19012 34692 19022
rect 34636 18918 34692 18956
rect 34972 19012 35028 19022
rect 34972 18918 35028 18956
rect 35084 18676 35140 21534
rect 35644 21588 35700 21598
rect 35644 21494 35700 21532
rect 35756 21588 35812 21598
rect 36092 21588 36148 21646
rect 35756 21586 36148 21588
rect 35756 21534 35758 21586
rect 35810 21534 36148 21586
rect 35756 21532 36148 21534
rect 35756 21522 35812 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35420 19124 35476 19134
rect 35420 19030 35476 19068
rect 35980 19012 36036 19022
rect 35084 18610 35140 18620
rect 35868 19010 36036 19012
rect 35868 18958 35982 19010
rect 36034 18958 36036 19010
rect 35868 18956 36036 18958
rect 34748 18452 34804 18462
rect 34748 17668 34804 18396
rect 35308 18452 35364 18462
rect 35868 18452 35924 18956
rect 35980 18946 36036 18956
rect 36092 18900 36148 21532
rect 36092 18834 36148 18844
rect 35308 18450 35588 18452
rect 35308 18398 35310 18450
rect 35362 18398 35588 18450
rect 35308 18396 35588 18398
rect 35308 18386 35364 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 18396
rect 35868 18386 35924 18396
rect 35980 18564 36036 18574
rect 35980 18450 36036 18508
rect 35980 18398 35982 18450
rect 36034 18398 36036 18450
rect 35980 18386 36036 18398
rect 35308 17836 35532 17892
rect 35084 17668 35140 17678
rect 34748 17666 35140 17668
rect 34748 17614 35086 17666
rect 35138 17614 35140 17666
rect 34748 17612 35140 17614
rect 35084 17444 35140 17612
rect 35084 17378 35140 17388
rect 35308 16772 35364 17836
rect 35532 17798 35588 17836
rect 35532 17668 35588 17678
rect 36204 17668 36260 25340
rect 36764 25060 36820 26126
rect 36988 25506 37044 26852
rect 37996 26516 38052 27022
rect 38108 28196 38164 28206
rect 38108 27970 38164 28140
rect 38108 27918 38110 27970
rect 38162 27918 38164 27970
rect 38108 27860 38164 27918
rect 38108 26964 38164 27804
rect 38220 27970 38276 27982
rect 38220 27918 38222 27970
rect 38274 27918 38276 27970
rect 38220 27300 38276 27918
rect 38220 27234 38276 27244
rect 38220 26964 38276 26974
rect 38108 26962 38276 26964
rect 38108 26910 38222 26962
rect 38274 26910 38276 26962
rect 38108 26908 38276 26910
rect 38220 26898 38276 26908
rect 38332 26740 38388 33292
rect 38444 33282 38500 33292
rect 38444 32562 38500 32574
rect 38444 32510 38446 32562
rect 38498 32510 38500 32562
rect 38444 31780 38500 32510
rect 38444 31714 38500 31724
rect 38556 31668 38612 34636
rect 38780 34626 38836 34636
rect 38780 34468 38836 34478
rect 38780 34132 38836 34412
rect 39228 34132 39284 34142
rect 38780 34130 39396 34132
rect 38780 34078 38782 34130
rect 38834 34078 39230 34130
rect 39282 34078 39396 34130
rect 38780 34076 39396 34078
rect 38780 34066 38836 34076
rect 39228 34066 39284 34076
rect 39116 33460 39172 33470
rect 38892 33348 38948 33358
rect 38892 33254 38948 33292
rect 39116 33234 39172 33404
rect 39116 33182 39118 33234
rect 39170 33182 39172 33234
rect 39116 33170 39172 33182
rect 39340 32786 39396 34076
rect 39340 32734 39342 32786
rect 39394 32734 39396 32786
rect 39340 32722 39396 32734
rect 39452 32788 39508 35644
rect 39676 34020 39732 34030
rect 39788 34020 39844 43652
rect 40124 43652 40180 43662
rect 41020 43652 41188 43708
rect 40124 42866 40180 43596
rect 41020 43540 41076 43550
rect 41020 43446 41076 43484
rect 40348 43428 40404 43438
rect 40348 43334 40404 43372
rect 40124 42814 40126 42866
rect 40178 42814 40180 42866
rect 40124 42802 40180 42814
rect 41020 42532 41076 42542
rect 41132 42532 41188 43652
rect 41356 43540 41412 49420
rect 41916 49028 41972 49870
rect 42252 49812 42308 50542
rect 42812 50596 42868 50606
rect 42812 50428 42868 50540
rect 42812 50372 42980 50428
rect 42140 49700 42196 49710
rect 41692 49026 41972 49028
rect 41692 48974 41918 49026
rect 41970 48974 41972 49026
rect 41692 48972 41972 48974
rect 41692 48466 41748 48972
rect 41916 48962 41972 48972
rect 42028 49644 42140 49700
rect 42028 49026 42084 49644
rect 42140 49606 42196 49644
rect 42252 49364 42308 49756
rect 42140 49308 42308 49364
rect 42140 49138 42196 49308
rect 42140 49086 42142 49138
rect 42194 49086 42196 49138
rect 42140 49074 42196 49086
rect 42028 48974 42030 49026
rect 42082 48974 42084 49026
rect 41692 48414 41694 48466
rect 41746 48414 41748 48466
rect 41692 48402 41748 48414
rect 41580 48132 41636 48142
rect 41580 46004 41636 48076
rect 41692 47572 41748 47582
rect 41692 47460 41748 47516
rect 42028 47460 42084 48974
rect 42252 49028 42308 49038
rect 42812 49028 42868 49038
rect 42252 49026 42868 49028
rect 42252 48974 42254 49026
rect 42306 48974 42814 49026
rect 42866 48974 42868 49026
rect 42252 48972 42868 48974
rect 42252 48962 42308 48972
rect 42364 48802 42420 48814
rect 42364 48750 42366 48802
rect 42418 48750 42420 48802
rect 42364 48356 42420 48750
rect 42476 48466 42532 48972
rect 42812 48962 42868 48972
rect 42476 48414 42478 48466
rect 42530 48414 42532 48466
rect 42476 48402 42532 48414
rect 42364 48262 42420 48300
rect 42588 48132 42644 48142
rect 42476 48018 42532 48030
rect 42476 47966 42478 48018
rect 42530 47966 42532 48018
rect 41692 47458 42084 47460
rect 41692 47406 41694 47458
rect 41746 47406 42084 47458
rect 41692 47404 42084 47406
rect 42140 47572 42196 47582
rect 41692 47394 41748 47404
rect 41692 46564 41748 46574
rect 41692 46470 41748 46508
rect 41692 46004 41748 46014
rect 41580 46002 41748 46004
rect 41580 45950 41694 46002
rect 41746 45950 41748 46002
rect 41580 45948 41748 45950
rect 41692 45938 41748 45948
rect 42140 46002 42196 47516
rect 42476 47458 42532 47966
rect 42476 47406 42478 47458
rect 42530 47406 42532 47458
rect 42476 47394 42532 47406
rect 42588 47346 42644 48076
rect 42924 47572 42980 50372
rect 43148 48916 43204 48926
rect 43260 48916 43316 51324
rect 43372 49700 43428 51886
rect 43708 51604 43764 51614
rect 43708 51378 43764 51548
rect 43708 51326 43710 51378
rect 43762 51326 43764 51378
rect 43708 51314 43764 51326
rect 43372 49634 43428 49644
rect 43596 51268 43652 51278
rect 43148 48914 43316 48916
rect 43148 48862 43150 48914
rect 43202 48862 43316 48914
rect 43148 48860 43316 48862
rect 43148 48850 43204 48860
rect 43036 48802 43092 48814
rect 43036 48750 43038 48802
rect 43090 48750 43092 48802
rect 43036 48244 43092 48750
rect 43036 48178 43092 48188
rect 43260 48242 43316 48860
rect 43372 48356 43428 48366
rect 43372 48262 43428 48300
rect 43260 48190 43262 48242
rect 43314 48190 43316 48242
rect 42924 47506 42980 47516
rect 42588 47294 42590 47346
rect 42642 47294 42644 47346
rect 42588 47282 42644 47294
rect 43260 46788 43316 48190
rect 43484 48244 43540 48254
rect 43484 47236 43540 48188
rect 43596 48020 43652 51212
rect 44156 50596 44212 51996
rect 44380 51268 44436 51278
rect 44380 51266 44996 51268
rect 44380 51214 44382 51266
rect 44434 51214 44996 51266
rect 44380 51212 44996 51214
rect 44380 51202 44436 51212
rect 44940 50706 44996 51212
rect 44940 50654 44942 50706
rect 44994 50654 44996 50706
rect 44940 50642 44996 50654
rect 44156 50530 44212 50540
rect 44828 50596 44884 50606
rect 44828 50502 44884 50540
rect 45500 50594 45556 52220
rect 45500 50542 45502 50594
rect 45554 50542 45556 50594
rect 45500 50530 45556 50542
rect 45836 50596 45892 50606
rect 45836 50502 45892 50540
rect 46060 50596 46116 54462
rect 46396 54516 46452 54526
rect 46396 54422 46452 54460
rect 46620 54514 46676 54526
rect 46620 54462 46622 54514
rect 46674 54462 46676 54514
rect 46620 53172 46676 54462
rect 46956 54516 47012 55132
rect 46956 54450 47012 54460
rect 46844 54404 46900 54414
rect 46844 54310 46900 54348
rect 47180 54404 47236 54414
rect 47740 54404 47796 55356
rect 47180 54402 47796 54404
rect 47180 54350 47182 54402
rect 47234 54350 47796 54402
rect 47180 54348 47796 54350
rect 47852 54404 47908 55918
rect 47180 54338 47236 54348
rect 47852 53844 47908 54348
rect 47516 53284 47572 53294
rect 46172 53170 46676 53172
rect 46172 53118 46622 53170
rect 46674 53118 46676 53170
rect 46172 53116 46676 53118
rect 46172 52722 46228 53116
rect 46620 53106 46676 53116
rect 46844 53172 46900 53182
rect 46900 53116 47012 53172
rect 46844 53078 46900 53116
rect 46396 52948 46452 52958
rect 46396 52854 46452 52892
rect 46732 52948 46788 52958
rect 46508 52836 46564 52846
rect 46732 52836 46788 52892
rect 46508 52742 46564 52780
rect 46620 52780 46788 52836
rect 46172 52670 46174 52722
rect 46226 52670 46228 52722
rect 46172 52658 46228 52670
rect 46620 52162 46676 52780
rect 46732 52276 46788 52314
rect 46732 52210 46788 52220
rect 46620 52110 46622 52162
rect 46674 52110 46676 52162
rect 46620 52098 46676 52110
rect 46956 52164 47012 53116
rect 47516 53170 47572 53228
rect 47516 53118 47518 53170
rect 47570 53118 47572 53170
rect 47068 52946 47124 52958
rect 47068 52894 47070 52946
rect 47122 52894 47124 52946
rect 47068 52724 47124 52894
rect 47516 52948 47572 53118
rect 47292 52724 47348 52734
rect 47068 52722 47348 52724
rect 47068 52670 47294 52722
rect 47346 52670 47348 52722
rect 47068 52668 47348 52670
rect 47292 52658 47348 52668
rect 47180 52500 47236 52510
rect 46956 52108 47124 52164
rect 47068 52050 47124 52108
rect 47068 51998 47070 52050
rect 47122 51998 47124 52050
rect 47068 51986 47124 51998
rect 46844 51938 46900 51950
rect 46844 51886 46846 51938
rect 46898 51886 46900 51938
rect 46844 51380 46900 51886
rect 47180 51602 47236 52444
rect 47292 52052 47348 52062
rect 47292 52050 47460 52052
rect 47292 51998 47294 52050
rect 47346 51998 47460 52050
rect 47292 51996 47460 51998
rect 47292 51986 47348 51996
rect 47180 51550 47182 51602
rect 47234 51550 47236 51602
rect 47180 51538 47236 51550
rect 46956 51380 47012 51390
rect 46508 51378 47012 51380
rect 46508 51326 46958 51378
rect 47010 51326 47012 51378
rect 46508 51324 47012 51326
rect 46508 51266 46564 51324
rect 46956 51314 47012 51324
rect 47292 51380 47348 51390
rect 47292 51286 47348 51324
rect 46508 51214 46510 51266
rect 46562 51214 46564 51266
rect 46508 51202 46564 51214
rect 47404 50932 47460 51996
rect 47180 50876 47460 50932
rect 46060 50530 46116 50540
rect 46732 50596 46788 50606
rect 47180 50596 47236 50876
rect 46732 50502 46788 50540
rect 46844 50594 47236 50596
rect 46844 50542 47182 50594
rect 47234 50542 47236 50594
rect 46844 50540 47236 50542
rect 45052 50372 45108 50382
rect 44940 50370 45108 50372
rect 44940 50318 45054 50370
rect 45106 50318 45108 50370
rect 44940 50316 45108 50318
rect 43596 47954 43652 47964
rect 43932 48242 43988 48254
rect 43932 48190 43934 48242
rect 43986 48190 43988 48242
rect 43484 47170 43540 47180
rect 43596 47572 43652 47582
rect 43260 46722 43316 46732
rect 42140 45950 42142 46002
rect 42194 45950 42196 46002
rect 42140 44324 42196 45950
rect 43596 45108 43652 47516
rect 43932 47012 43988 48190
rect 44268 47572 44324 47582
rect 44268 47478 44324 47516
rect 44828 47572 44884 47582
rect 44828 47458 44884 47516
rect 44828 47406 44830 47458
rect 44882 47406 44884 47458
rect 44828 47394 44884 47406
rect 43932 46946 43988 46956
rect 44828 47236 44884 47246
rect 44492 46676 44548 46686
rect 44492 46582 44548 46620
rect 44828 46674 44884 47180
rect 44828 46622 44830 46674
rect 44882 46622 44884 46674
rect 44828 46610 44884 46622
rect 44940 46452 44996 50316
rect 45052 50306 45108 50316
rect 46732 49140 46788 49150
rect 46844 49140 46900 50540
rect 47180 50530 47236 50540
rect 47404 50596 47460 50606
rect 47516 50596 47572 52892
rect 47628 52722 47684 52734
rect 47628 52670 47630 52722
rect 47682 52670 47684 52722
rect 47628 52276 47684 52670
rect 47628 52274 47796 52276
rect 47628 52222 47630 52274
rect 47682 52222 47796 52274
rect 47628 52220 47796 52222
rect 47628 52210 47684 52220
rect 47404 50594 47572 50596
rect 47404 50542 47406 50594
rect 47458 50542 47572 50594
rect 47404 50540 47572 50542
rect 47404 50530 47460 50540
rect 47516 50428 47572 50540
rect 47628 51378 47684 51390
rect 47628 51326 47630 51378
rect 47682 51326 47684 51378
rect 47628 50596 47684 51326
rect 47740 51044 47796 52220
rect 47852 51266 47908 53788
rect 47964 53284 48020 56252
rect 48076 56082 48132 57372
rect 48188 57362 48244 57372
rect 48188 56306 48244 56318
rect 48188 56254 48190 56306
rect 48242 56254 48244 56306
rect 48188 56196 48244 56254
rect 48188 56130 48244 56140
rect 48076 56030 48078 56082
rect 48130 56030 48132 56082
rect 48076 56018 48132 56030
rect 47964 53170 48020 53228
rect 47964 53118 47966 53170
rect 48018 53118 48020 53170
rect 47964 53106 48020 53118
rect 48300 51604 48356 51614
rect 48300 51510 48356 51548
rect 47852 51214 47854 51266
rect 47906 51214 47908 51266
rect 47852 51202 47908 51214
rect 48188 51266 48244 51278
rect 48188 51214 48190 51266
rect 48242 51214 48244 51266
rect 48188 51044 48244 51214
rect 47740 50988 48244 51044
rect 47628 50530 47684 50540
rect 47852 50482 47908 50494
rect 47852 50430 47854 50482
rect 47906 50430 47908 50482
rect 47852 50428 47908 50430
rect 46732 49138 46900 49140
rect 46732 49086 46734 49138
rect 46786 49086 46900 49138
rect 46732 49084 46900 49086
rect 46956 50370 47012 50382
rect 46956 50318 46958 50370
rect 47010 50318 47012 50370
rect 46732 49074 46788 49084
rect 45612 47346 45668 47358
rect 45612 47294 45614 47346
rect 45666 47294 45668 47346
rect 45276 47012 45332 47022
rect 44156 46396 44996 46452
rect 45052 46564 45108 46574
rect 43820 45108 43876 45118
rect 43596 45106 43876 45108
rect 43596 45054 43822 45106
rect 43874 45054 43876 45106
rect 43596 45052 43876 45054
rect 43820 45042 43876 45052
rect 43596 44436 43652 44446
rect 43596 44434 44100 44436
rect 43596 44382 43598 44434
rect 43650 44382 44100 44434
rect 43596 44380 44100 44382
rect 43596 44370 43652 44380
rect 41468 44210 41524 44222
rect 41468 44158 41470 44210
rect 41522 44158 41524 44210
rect 41468 43708 41524 44158
rect 42140 43708 42196 44268
rect 43932 44210 43988 44222
rect 43932 44158 43934 44210
rect 43986 44158 43988 44210
rect 43932 43708 43988 44158
rect 41468 43652 41636 43708
rect 42140 43652 42532 43708
rect 41468 43540 41524 43550
rect 41356 43484 41468 43540
rect 41468 43446 41524 43484
rect 41580 42866 41636 43652
rect 41580 42814 41582 42866
rect 41634 42814 41636 42866
rect 41580 42802 41636 42814
rect 42252 43428 42308 43438
rect 42252 42980 42308 43372
rect 42476 43428 42532 43652
rect 43708 43652 43988 43708
rect 44044 44210 44100 44380
rect 44044 44158 44046 44210
rect 44098 44158 44100 44210
rect 42476 43334 42532 43372
rect 43036 43428 43092 43438
rect 41692 42644 41748 42654
rect 42028 42644 42084 42654
rect 41692 42642 42084 42644
rect 41692 42590 41694 42642
rect 41746 42590 42030 42642
rect 42082 42590 42084 42642
rect 41692 42588 42084 42590
rect 41692 42578 41748 42588
rect 42028 42578 42084 42588
rect 42252 42642 42308 42924
rect 42252 42590 42254 42642
rect 42306 42590 42308 42642
rect 42252 42578 42308 42590
rect 41468 42532 41524 42542
rect 41020 42530 41636 42532
rect 41020 42478 41022 42530
rect 41074 42478 41470 42530
rect 41522 42478 41636 42530
rect 41020 42476 41636 42478
rect 41020 42466 41076 42476
rect 41468 42466 41524 42476
rect 40348 41972 40404 41982
rect 41132 41972 41188 41982
rect 40348 41878 40404 41916
rect 41020 41970 41188 41972
rect 41020 41918 41134 41970
rect 41186 41918 41188 41970
rect 41020 41916 41188 41918
rect 40124 41300 40180 41310
rect 40124 41298 40292 41300
rect 40124 41246 40126 41298
rect 40178 41246 40292 41298
rect 40124 41244 40292 41246
rect 40124 41234 40180 41244
rect 40236 40514 40292 41244
rect 40236 40462 40238 40514
rect 40290 40462 40292 40514
rect 40236 40404 40292 40462
rect 40348 41188 40404 41198
rect 40348 40514 40404 41132
rect 40348 40462 40350 40514
rect 40402 40462 40404 40514
rect 40348 40404 40404 40462
rect 40796 40404 40852 40414
rect 41020 40404 41076 41916
rect 41132 41906 41188 41916
rect 41356 41972 41412 41982
rect 41356 41970 41524 41972
rect 41356 41918 41358 41970
rect 41410 41918 41524 41970
rect 41356 41916 41524 41918
rect 41356 41906 41412 41916
rect 41244 41858 41300 41870
rect 41244 41806 41246 41858
rect 41298 41806 41300 41858
rect 41132 41076 41188 41086
rect 41132 40626 41188 41020
rect 41132 40574 41134 40626
rect 41186 40574 41188 40626
rect 41132 40562 41188 40574
rect 41244 40628 41300 41806
rect 41244 40572 41412 40628
rect 40348 40402 41076 40404
rect 40348 40350 40798 40402
rect 40850 40350 41076 40402
rect 40348 40348 41076 40350
rect 41244 40404 41300 40414
rect 40236 40338 40292 40348
rect 40796 40338 40852 40348
rect 41244 40310 41300 40348
rect 41356 40402 41412 40572
rect 41356 40350 41358 40402
rect 41410 40350 41412 40402
rect 41356 40338 41412 40350
rect 41468 40404 41524 41916
rect 41468 40338 41524 40348
rect 40236 40178 40292 40190
rect 40236 40126 40238 40178
rect 40290 40126 40292 40178
rect 40012 38834 40068 38846
rect 40012 38782 40014 38834
rect 40066 38782 40068 38834
rect 39900 37492 39956 37502
rect 40012 37492 40068 38782
rect 40236 38612 40292 40126
rect 41580 39508 41636 42476
rect 41804 41972 41860 41982
rect 41804 40740 41860 41916
rect 43036 41300 43092 43372
rect 43596 42980 43652 42990
rect 43708 42980 43764 43652
rect 44044 43092 44100 44158
rect 44156 43652 44212 46396
rect 45052 45890 45108 46508
rect 45052 45838 45054 45890
rect 45106 45838 45108 45890
rect 45052 45826 45108 45838
rect 45276 45890 45332 46956
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45444 45332 45838
rect 45388 46676 45444 46686
rect 45388 45892 45444 46620
rect 45500 45892 45556 45902
rect 45388 45890 45556 45892
rect 45388 45838 45502 45890
rect 45554 45838 45556 45890
rect 45388 45836 45556 45838
rect 45500 45826 45556 45836
rect 45388 45668 45444 45678
rect 45612 45668 45668 47294
rect 45948 47012 46004 47022
rect 45948 46898 46004 46956
rect 45948 46846 45950 46898
rect 46002 46846 46004 46898
rect 45948 46834 46004 46846
rect 46172 46786 46228 46798
rect 46172 46734 46174 46786
rect 46226 46734 46228 46786
rect 45724 46676 45780 46686
rect 45724 46582 45780 46620
rect 45836 46564 45892 46574
rect 45836 46470 45892 46508
rect 45388 45666 45668 45668
rect 45388 45614 45390 45666
rect 45442 45614 45668 45666
rect 45388 45612 45668 45614
rect 45948 45668 46004 45678
rect 46172 45668 46228 46734
rect 45948 45666 46228 45668
rect 45948 45614 45950 45666
rect 46002 45614 46228 45666
rect 45948 45612 46228 45614
rect 45388 45602 45444 45612
rect 45276 45388 45444 45444
rect 45388 44546 45444 45388
rect 45388 44494 45390 44546
rect 45442 44494 45444 44546
rect 45388 44482 45444 44494
rect 45500 44434 45556 44446
rect 45500 44382 45502 44434
rect 45554 44382 45556 44434
rect 44268 44324 44324 44334
rect 44716 44324 44772 44334
rect 44268 44322 44772 44324
rect 44268 44270 44270 44322
rect 44322 44270 44718 44322
rect 44770 44270 44772 44322
rect 44268 44268 44772 44270
rect 44268 44258 44324 44268
rect 44716 44258 44772 44268
rect 44156 43586 44212 43596
rect 44268 43988 44324 43998
rect 43484 42924 43596 42980
rect 43652 42924 43764 42980
rect 43932 43036 44100 43092
rect 43484 42082 43540 42924
rect 43596 42914 43652 42924
rect 43932 42644 43988 43036
rect 44156 42980 44212 42990
rect 44156 42866 44212 42924
rect 44156 42814 44158 42866
rect 44210 42814 44212 42866
rect 44156 42802 44212 42814
rect 43820 42642 43988 42644
rect 43820 42590 43934 42642
rect 43986 42590 43988 42642
rect 43820 42588 43988 42590
rect 43484 42030 43486 42082
rect 43538 42030 43540 42082
rect 43484 42018 43540 42030
rect 43708 42532 43764 42542
rect 43484 41300 43540 41310
rect 43036 41298 43540 41300
rect 43036 41246 43486 41298
rect 43538 41246 43540 41298
rect 43036 41244 43540 41246
rect 43036 41186 43092 41244
rect 43484 41234 43540 41244
rect 43036 41134 43038 41186
rect 43090 41134 43092 41186
rect 43036 41122 43092 41134
rect 42252 41076 42308 41086
rect 42252 40982 42308 41020
rect 41692 39618 41748 39630
rect 41692 39566 41694 39618
rect 41746 39566 41748 39618
rect 41692 39508 41748 39566
rect 40684 39452 41748 39508
rect 40684 38668 40740 39452
rect 40236 38050 40292 38556
rect 40236 37998 40238 38050
rect 40290 37998 40292 38050
rect 40236 37986 40292 37998
rect 40460 38612 40740 38668
rect 39900 37490 40068 37492
rect 39900 37438 39902 37490
rect 39954 37438 40068 37490
rect 39900 37436 40068 37438
rect 39900 37426 39956 37436
rect 39732 33964 39844 34020
rect 40236 34468 40292 34478
rect 39676 33926 39732 33964
rect 39452 32722 39508 32732
rect 39788 33346 39844 33358
rect 39788 33294 39790 33346
rect 39842 33294 39844 33346
rect 38892 32450 38948 32462
rect 38892 32398 38894 32450
rect 38946 32398 38948 32450
rect 38892 32228 38948 32398
rect 38892 32162 38948 32172
rect 39564 32340 39620 32350
rect 39564 31890 39620 32284
rect 39564 31838 39566 31890
rect 39618 31838 39620 31890
rect 39564 31826 39620 31838
rect 38556 31602 38612 31612
rect 38892 31778 38948 31790
rect 38892 31726 38894 31778
rect 38946 31726 38948 31778
rect 38892 29988 38948 31726
rect 38668 29932 38892 29988
rect 38668 28644 38724 29932
rect 38892 29922 38948 29932
rect 39788 30324 39844 33294
rect 39900 33348 39956 33358
rect 39900 32562 39956 33292
rect 40236 33346 40292 34412
rect 40348 34132 40404 34142
rect 40348 34038 40404 34076
rect 40236 33294 40238 33346
rect 40290 33294 40292 33346
rect 40236 33282 40292 33294
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39900 32452 39956 32510
rect 39900 32386 39956 32396
rect 39900 30324 39956 30334
rect 39788 30322 39956 30324
rect 39788 30270 39902 30322
rect 39954 30270 39956 30322
rect 39788 30268 39956 30270
rect 39788 29876 39844 30268
rect 39900 30258 39956 30268
rect 40348 29988 40404 29998
rect 40348 29894 40404 29932
rect 39788 29810 39844 29820
rect 40236 29316 40292 29326
rect 40236 29222 40292 29260
rect 40124 29204 40180 29214
rect 38668 28550 38724 28588
rect 38892 29202 40180 29204
rect 38892 29150 40126 29202
rect 40178 29150 40180 29202
rect 38892 29148 40180 29150
rect 38892 28082 38948 29148
rect 40124 29138 40180 29148
rect 39340 28532 39396 28542
rect 39340 28530 39508 28532
rect 39340 28478 39342 28530
rect 39394 28478 39508 28530
rect 39340 28476 39508 28478
rect 39340 28466 39396 28476
rect 38892 28030 38894 28082
rect 38946 28030 38948 28082
rect 38892 28018 38948 28030
rect 38444 27972 38500 27982
rect 38444 27878 38500 27916
rect 39004 27972 39060 27982
rect 39004 27878 39060 27916
rect 39116 27970 39172 27982
rect 39116 27918 39118 27970
rect 39170 27918 39172 27970
rect 38668 27860 38724 27870
rect 38668 27766 38724 27804
rect 39116 27636 39172 27918
rect 39452 27746 39508 28476
rect 39452 27694 39454 27746
rect 39506 27694 39508 27746
rect 39452 27682 39508 27694
rect 40012 28084 40068 28094
rect 39116 27570 39172 27580
rect 40012 27076 40068 28028
rect 38668 26964 38724 27002
rect 40012 26982 40068 27020
rect 38668 26898 38724 26908
rect 39676 26964 39732 26974
rect 38332 26684 38612 26740
rect 37996 26450 38052 26460
rect 38444 26516 38500 26526
rect 37660 26180 37716 26190
rect 37436 26178 37716 26180
rect 37436 26126 37662 26178
rect 37714 26126 37716 26178
rect 37436 26124 37716 26126
rect 36988 25454 36990 25506
rect 37042 25454 37044 25506
rect 36988 25442 37044 25454
rect 37212 25620 37268 25630
rect 37212 25506 37268 25564
rect 37212 25454 37214 25506
rect 37266 25454 37268 25506
rect 37100 25284 37156 25294
rect 37100 25190 37156 25228
rect 37212 25060 37268 25454
rect 37436 25396 37492 26124
rect 37660 26114 37716 26124
rect 38332 25620 38388 25630
rect 37996 25618 38388 25620
rect 37996 25566 38334 25618
rect 38386 25566 38388 25618
rect 37996 25564 38388 25566
rect 37548 25508 37604 25518
rect 37996 25508 38052 25564
rect 38332 25554 38388 25564
rect 37548 25506 38052 25508
rect 37548 25454 37550 25506
rect 37602 25454 38052 25506
rect 37548 25452 38052 25454
rect 38444 25506 38500 26460
rect 38444 25454 38446 25506
rect 38498 25454 38500 25506
rect 37548 25442 37604 25452
rect 38444 25442 38500 25454
rect 37436 25330 37492 25340
rect 37996 25284 38052 25294
rect 37996 25190 38052 25228
rect 38220 25284 38276 25294
rect 38556 25284 38612 26684
rect 39228 26516 39284 26526
rect 39228 26422 39284 26460
rect 39452 26292 39508 26302
rect 39452 26198 39508 26236
rect 39340 26180 39396 26190
rect 39116 26068 39172 26078
rect 39116 25974 39172 26012
rect 39004 25620 39060 25630
rect 39340 25620 39396 26124
rect 39004 25618 39396 25620
rect 39004 25566 39006 25618
rect 39058 25566 39342 25618
rect 39394 25566 39396 25618
rect 39004 25564 39396 25566
rect 39004 25554 39060 25564
rect 39340 25554 39396 25564
rect 39676 25508 39732 26908
rect 39788 26404 39844 26414
rect 39844 26348 39956 26404
rect 39788 26310 39844 26348
rect 39788 26068 39844 26078
rect 39788 25730 39844 26012
rect 39788 25678 39790 25730
rect 39842 25678 39844 25730
rect 39788 25666 39844 25678
rect 39900 25730 39956 26348
rect 40124 26290 40180 26302
rect 40124 26238 40126 26290
rect 40178 26238 40180 26290
rect 40124 26180 40180 26238
rect 40124 26114 40180 26124
rect 39900 25678 39902 25730
rect 39954 25678 39956 25730
rect 39900 25666 39956 25678
rect 40012 25620 40068 25630
rect 39676 25452 39956 25508
rect 38220 25282 38612 25284
rect 38220 25230 38222 25282
rect 38274 25230 38612 25282
rect 38220 25228 38612 25230
rect 39228 25396 39284 25406
rect 36764 25004 37268 25060
rect 36876 24500 36932 25004
rect 36876 24434 36932 24444
rect 37884 24724 37940 24734
rect 37884 23380 37940 24668
rect 38220 24610 38276 25228
rect 39228 24946 39284 25340
rect 39228 24894 39230 24946
rect 39282 24894 39284 24946
rect 39228 24882 39284 24894
rect 38220 24558 38222 24610
rect 38274 24558 38276 24610
rect 38220 24546 38276 24558
rect 38444 24724 38500 24734
rect 38444 24050 38500 24668
rect 38444 23998 38446 24050
rect 38498 23998 38500 24050
rect 38444 23986 38500 23998
rect 38668 24610 38724 24622
rect 38668 24558 38670 24610
rect 38722 24558 38724 24610
rect 36428 23156 36484 23166
rect 36428 22484 36484 23100
rect 36428 22390 36484 22428
rect 37212 22372 37268 22382
rect 37212 22258 37268 22316
rect 37884 22370 37940 23324
rect 38108 23268 38164 23278
rect 38108 23156 38164 23212
rect 38444 23156 38500 23166
rect 38108 23154 38276 23156
rect 38108 23102 38110 23154
rect 38162 23102 38276 23154
rect 38108 23100 38276 23102
rect 38108 23090 38164 23100
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37884 22306 37940 22318
rect 37212 22206 37214 22258
rect 37266 22206 37268 22258
rect 36316 21812 36372 21822
rect 36316 21586 36372 21756
rect 36764 21812 36820 21822
rect 36764 21718 36820 21756
rect 36316 21534 36318 21586
rect 36370 21534 36372 21586
rect 36316 21522 36372 21534
rect 37100 21698 37156 21710
rect 37100 21646 37102 21698
rect 37154 21646 37156 21698
rect 35420 17666 36260 17668
rect 35420 17614 35534 17666
rect 35586 17614 36260 17666
rect 35420 17612 36260 17614
rect 36428 20244 36484 20254
rect 35420 17108 35476 17612
rect 35532 17602 35588 17612
rect 35420 17042 35476 17052
rect 35980 17444 36036 17454
rect 35084 16716 35364 16772
rect 35980 16772 36036 17388
rect 35980 16716 36260 16772
rect 34636 15428 34692 15438
rect 34636 15334 34692 15372
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 34300 13794 34356 13806
rect 34412 15092 34580 15148
rect 35084 15314 35140 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 36092 16322 36148 16334
rect 36092 16270 36094 16322
rect 36146 16270 36148 16322
rect 35532 16212 35588 16222
rect 35308 15986 35364 15998
rect 35308 15934 35310 15986
rect 35362 15934 35364 15986
rect 35308 15428 35364 15934
rect 35532 15986 35588 16156
rect 35644 16212 35700 16222
rect 36092 16212 36148 16270
rect 35644 16210 35812 16212
rect 35644 16158 35646 16210
rect 35698 16158 35812 16210
rect 35644 16156 35812 16158
rect 35644 16146 35700 16156
rect 35532 15934 35534 15986
rect 35586 15934 35588 15986
rect 35532 15764 35588 15934
rect 35532 15698 35588 15708
rect 35308 15362 35364 15372
rect 35756 15426 35812 16156
rect 36092 16118 36148 16156
rect 35756 15374 35758 15426
rect 35810 15374 35812 15426
rect 35756 15362 35812 15374
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 34412 13524 34468 15092
rect 35084 14084 35140 15262
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14028 35252 14084
rect 34524 13972 34580 13982
rect 34580 13916 34804 13972
rect 34524 13906 34580 13916
rect 34076 13346 34132 13356
rect 34188 13468 34468 13524
rect 34524 13746 34580 13758
rect 34524 13694 34526 13746
rect 34578 13694 34580 13746
rect 33964 13188 34020 13198
rect 33964 12738 34020 13132
rect 33964 12686 33966 12738
rect 34018 12686 34020 12738
rect 33964 12674 34020 12686
rect 34188 12292 34244 13468
rect 34524 13412 34580 13694
rect 34076 12236 34244 12292
rect 34412 13356 34580 13412
rect 33964 11284 34020 11294
rect 33964 11190 34020 11228
rect 33852 10108 34020 10164
rect 32172 9762 32228 9772
rect 32844 9714 32900 9996
rect 32956 9996 33796 10052
rect 32956 9826 33012 9996
rect 32956 9774 32958 9826
rect 33010 9774 33012 9826
rect 32956 9762 33012 9774
rect 33292 9828 33348 9838
rect 33516 9828 33572 9838
rect 33292 9734 33348 9772
rect 33404 9826 33572 9828
rect 33404 9774 33518 9826
rect 33570 9774 33572 9826
rect 33404 9772 33572 9774
rect 32844 9662 32846 9714
rect 32898 9662 32900 9714
rect 32620 9602 32676 9614
rect 32620 9550 32622 9602
rect 32674 9550 32676 9602
rect 31612 8204 32116 8260
rect 31612 8036 31668 8046
rect 31612 7942 31668 7980
rect 31724 8034 31780 8046
rect 31724 7982 31726 8034
rect 31778 7982 31780 8034
rect 30940 7634 30996 7644
rect 31276 7868 31556 7924
rect 30940 6692 30996 6702
rect 31276 6692 31332 7868
rect 31500 7700 31556 7710
rect 31500 7606 31556 7644
rect 31724 7364 31780 7982
rect 31724 7298 31780 7308
rect 31836 7362 31892 7374
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31836 6692 31892 7310
rect 30940 6690 31332 6692
rect 30940 6638 30942 6690
rect 30994 6638 31278 6690
rect 31330 6638 31332 6690
rect 30940 6636 31332 6638
rect 30940 6626 30996 6636
rect 31276 6626 31332 6636
rect 31724 6636 31836 6692
rect 31500 6580 31556 6590
rect 31500 6486 31556 6524
rect 30716 6468 30772 6478
rect 30716 6374 30772 6412
rect 30828 6466 30884 6478
rect 30828 6414 30830 6466
rect 30882 6414 30884 6466
rect 30828 6130 30884 6414
rect 31388 6466 31444 6478
rect 31388 6414 31390 6466
rect 31442 6414 31444 6466
rect 31388 6244 31444 6414
rect 31388 6188 31668 6244
rect 30828 6078 30830 6130
rect 30882 6078 30884 6130
rect 30828 6066 30884 6078
rect 31276 6132 31332 6142
rect 31276 6130 31556 6132
rect 31276 6078 31278 6130
rect 31330 6078 31556 6130
rect 31276 6076 31556 6078
rect 31276 6066 31332 6076
rect 30940 5906 30996 5918
rect 30940 5854 30942 5906
rect 30994 5854 30996 5906
rect 30604 5730 30660 5740
rect 30716 5794 30772 5806
rect 30716 5742 30718 5794
rect 30770 5742 30772 5794
rect 30716 5122 30772 5742
rect 30940 5796 30996 5854
rect 31388 5908 31444 5918
rect 31388 5814 31444 5852
rect 30996 5740 31220 5796
rect 30940 5702 30996 5740
rect 30940 5348 30996 5358
rect 30996 5292 31108 5348
rect 30940 5282 30996 5292
rect 31052 5234 31108 5292
rect 31052 5182 31054 5234
rect 31106 5182 31108 5234
rect 31052 5170 31108 5182
rect 30716 5070 30718 5122
rect 30770 5070 30772 5122
rect 30716 5058 30772 5070
rect 30940 5124 30996 5134
rect 30940 5030 30996 5068
rect 31164 5122 31220 5740
rect 31164 5070 31166 5122
rect 31218 5070 31220 5122
rect 31164 5058 31220 5070
rect 30380 4498 30436 4508
rect 31500 4450 31556 6076
rect 31612 6018 31668 6188
rect 31612 5966 31614 6018
rect 31666 5966 31668 6018
rect 31612 5954 31668 5966
rect 31612 5236 31668 5246
rect 31724 5236 31780 6636
rect 31836 6626 31892 6636
rect 31948 6802 32004 6814
rect 31948 6750 31950 6802
rect 32002 6750 32004 6802
rect 31948 6690 32004 6750
rect 31948 6638 31950 6690
rect 32002 6638 32004 6690
rect 31948 6244 32004 6638
rect 31948 6178 32004 6188
rect 31612 5234 31780 5236
rect 31612 5182 31614 5234
rect 31666 5182 31780 5234
rect 31612 5180 31780 5182
rect 32060 5684 32116 8204
rect 32172 8258 32228 8270
rect 32172 8206 32174 8258
rect 32226 8206 32228 8258
rect 32172 8036 32228 8206
rect 32508 8036 32564 8046
rect 32172 8034 32564 8036
rect 32172 7982 32510 8034
rect 32562 7982 32564 8034
rect 32172 7980 32564 7982
rect 32284 6914 32340 7980
rect 32508 7812 32564 7980
rect 32508 7746 32564 7756
rect 32620 7476 32676 9550
rect 32844 9604 32900 9662
rect 33404 9716 33460 9772
rect 33516 9762 33572 9772
rect 33404 9650 33460 9660
rect 32844 9548 33348 9604
rect 33292 9266 33348 9548
rect 33292 9214 33294 9266
rect 33346 9214 33348 9266
rect 33292 9202 33348 9214
rect 33516 9602 33572 9614
rect 33516 9550 33518 9602
rect 33570 9550 33572 9602
rect 33516 9154 33572 9550
rect 33740 9268 33796 9996
rect 33852 9940 33908 9950
rect 33852 9826 33908 9884
rect 33852 9774 33854 9826
rect 33906 9774 33908 9826
rect 33852 9762 33908 9774
rect 33964 9716 34020 10108
rect 33964 9650 34020 9660
rect 33852 9268 33908 9278
rect 33740 9266 33908 9268
rect 33740 9214 33854 9266
rect 33906 9214 33908 9266
rect 33740 9212 33908 9214
rect 33852 9202 33908 9212
rect 33516 9102 33518 9154
rect 33570 9102 33572 9154
rect 33516 8372 33572 9102
rect 33628 9156 33684 9166
rect 33628 9154 33796 9156
rect 33628 9102 33630 9154
rect 33682 9102 33796 9154
rect 33628 9100 33796 9102
rect 33628 9090 33684 9100
rect 33628 8372 33684 8382
rect 33516 8370 33684 8372
rect 33516 8318 33630 8370
rect 33682 8318 33684 8370
rect 33516 8316 33684 8318
rect 33628 8306 33684 8316
rect 33740 8260 33796 9100
rect 34076 8372 34132 12236
rect 34300 12178 34356 12190
rect 34300 12126 34302 12178
rect 34354 12126 34356 12178
rect 34300 12068 34356 12126
rect 34412 12180 34468 13356
rect 34636 13186 34692 13916
rect 34748 13746 34804 13916
rect 35084 13748 35140 13758
rect 34748 13694 34750 13746
rect 34802 13694 34804 13746
rect 34748 13682 34804 13694
rect 34860 13746 35140 13748
rect 34860 13694 35086 13746
rect 35138 13694 35140 13746
rect 34860 13692 35140 13694
rect 34636 13134 34638 13186
rect 34690 13134 34692 13186
rect 34636 13122 34692 13134
rect 34748 13188 34804 13198
rect 34860 13188 34916 13692
rect 35084 13682 35140 13692
rect 34972 13522 35028 13534
rect 35196 13524 35252 14028
rect 34972 13470 34974 13522
rect 35026 13470 35028 13522
rect 34972 13412 35028 13470
rect 34972 13346 35028 13356
rect 35084 13468 35252 13524
rect 35308 13860 35364 13870
rect 35756 13860 35812 13870
rect 35308 13858 35756 13860
rect 35308 13806 35310 13858
rect 35362 13806 35756 13858
rect 35308 13804 35756 13806
rect 35308 13524 35364 13804
rect 35756 13766 35812 13804
rect 34804 13132 34916 13188
rect 35084 13188 35140 13468
rect 35308 13458 35364 13468
rect 35532 13636 35588 13646
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13132 35364 13188
rect 34748 13094 34804 13132
rect 34972 13076 35028 13086
rect 34972 12982 35028 13020
rect 34524 12852 34580 12862
rect 34524 12402 34580 12796
rect 34636 12740 34692 12750
rect 34636 12738 34804 12740
rect 34636 12686 34638 12738
rect 34690 12686 34804 12738
rect 34636 12684 34804 12686
rect 34636 12674 34692 12684
rect 34524 12350 34526 12402
rect 34578 12350 34580 12402
rect 34524 12338 34580 12350
rect 34636 12180 34692 12190
rect 34412 12178 34692 12180
rect 34412 12126 34638 12178
rect 34690 12126 34692 12178
rect 34412 12124 34692 12126
rect 34300 12002 34356 12012
rect 34636 11956 34692 12124
rect 34748 12178 34804 12684
rect 34748 12126 34750 12178
rect 34802 12126 34804 12178
rect 34748 12114 34804 12126
rect 35308 12180 35364 13132
rect 35420 12852 35476 12862
rect 35420 12758 35476 12796
rect 35532 12292 35588 13580
rect 35644 13188 35700 13198
rect 35644 12962 35700 13132
rect 35644 12910 35646 12962
rect 35698 12910 35700 12962
rect 35644 12898 35700 12910
rect 35980 12852 36036 12862
rect 35980 12758 36036 12796
rect 35644 12738 35700 12750
rect 35644 12686 35646 12738
rect 35698 12686 35700 12738
rect 35644 12404 35700 12686
rect 35644 12348 36036 12404
rect 35532 12236 35812 12292
rect 35308 12178 35588 12180
rect 35308 12126 35310 12178
rect 35362 12126 35588 12178
rect 35308 12124 35588 12126
rect 35308 12114 35364 12124
rect 34636 11890 34692 11900
rect 35084 12068 35140 12078
rect 35084 11506 35140 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11454 35086 11506
rect 35138 11454 35140 11506
rect 35084 11442 35140 11454
rect 35532 11508 35588 12124
rect 35532 11442 35588 11452
rect 35532 11060 35588 11070
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 9940 35476 9950
rect 35532 9940 35588 11004
rect 35420 9938 35588 9940
rect 35420 9886 35422 9938
rect 35474 9886 35588 9938
rect 35420 9884 35588 9886
rect 35420 9874 35476 9884
rect 34636 9828 34692 9838
rect 34188 9716 34244 9726
rect 34188 9622 34244 9660
rect 34524 9714 34580 9726
rect 34524 9662 34526 9714
rect 34578 9662 34580 9714
rect 34524 9156 34580 9662
rect 34524 9090 34580 9100
rect 34076 8306 34132 8316
rect 33964 8260 34020 8270
rect 33740 8258 34020 8260
rect 33740 8206 33966 8258
rect 34018 8206 34020 8258
rect 33740 8204 34020 8206
rect 33740 8034 33796 8046
rect 33740 7982 33742 8034
rect 33794 7982 33796 8034
rect 32620 7410 32676 7420
rect 33628 7476 33684 7486
rect 33628 7382 33684 7420
rect 33740 7474 33796 7982
rect 33964 8036 34020 8204
rect 33964 7970 34020 7980
rect 33740 7422 33742 7474
rect 33794 7422 33796 7474
rect 33740 7410 33796 7422
rect 33964 7588 34020 7598
rect 33964 7252 34020 7532
rect 34300 7476 34356 7486
rect 34300 7382 34356 7420
rect 34412 7474 34468 7486
rect 34412 7422 34414 7474
rect 34466 7422 34468 7474
rect 32284 6862 32286 6914
rect 32338 6862 32340 6914
rect 32284 6802 32340 6862
rect 32284 6750 32286 6802
rect 32338 6750 32340 6802
rect 32284 6738 32340 6750
rect 33740 7196 34020 7252
rect 32508 6692 32564 6702
rect 32172 6468 32228 6478
rect 32172 6130 32228 6412
rect 32172 6078 32174 6130
rect 32226 6078 32228 6130
rect 32172 5908 32228 6078
rect 32508 6132 32564 6636
rect 33628 6356 33684 6366
rect 33740 6356 33796 7196
rect 34412 6580 34468 7422
rect 33684 6300 33796 6356
rect 33852 6524 34468 6580
rect 34636 7474 34692 9772
rect 35644 9828 35700 9838
rect 35644 9734 35700 9772
rect 35756 9604 35812 12236
rect 35980 12290 36036 12348
rect 35980 12238 35982 12290
rect 36034 12238 36036 12290
rect 35980 12226 36036 12238
rect 36204 11732 36260 16716
rect 36428 16322 36484 20188
rect 36988 19460 37044 19470
rect 36988 19234 37044 19404
rect 36988 19182 36990 19234
rect 37042 19182 37044 19234
rect 36988 19170 37044 19182
rect 37100 19236 37156 21646
rect 37212 21476 37268 22206
rect 37324 22260 37380 22270
rect 37324 22166 37380 22204
rect 37436 22258 37492 22270
rect 37436 22206 37438 22258
rect 37490 22206 37492 22258
rect 37436 21700 37492 22206
rect 38108 21700 38164 21710
rect 37436 21698 38164 21700
rect 37436 21646 38110 21698
rect 38162 21646 38164 21698
rect 37436 21644 38164 21646
rect 38108 21634 38164 21644
rect 37772 21476 37828 21486
rect 37212 21474 37828 21476
rect 37212 21422 37774 21474
rect 37826 21422 37828 21474
rect 37212 21420 37828 21422
rect 37772 21410 37828 21420
rect 37772 19908 37828 19918
rect 37436 19852 37772 19908
rect 37100 19170 37156 19180
rect 37212 19236 37268 19246
rect 37436 19236 37492 19852
rect 37772 19814 37828 19852
rect 37212 19234 37492 19236
rect 37212 19182 37214 19234
rect 37266 19182 37492 19234
rect 37212 19180 37492 19182
rect 37548 19236 37604 19246
rect 37996 19236 38052 19246
rect 37548 19234 38052 19236
rect 37548 19182 37550 19234
rect 37602 19182 37998 19234
rect 38050 19182 38052 19234
rect 37548 19180 38052 19182
rect 37100 19010 37156 19022
rect 37100 18958 37102 19010
rect 37154 18958 37156 19010
rect 37100 18564 37156 18958
rect 37100 18498 37156 18508
rect 37212 18340 37268 19180
rect 37548 19170 37604 19180
rect 37996 19170 38052 19180
rect 37884 19010 37940 19022
rect 37884 18958 37886 19010
rect 37938 18958 37940 19010
rect 37884 18900 37940 18958
rect 37884 18834 37940 18844
rect 38108 19010 38164 19022
rect 38108 18958 38110 19010
rect 38162 18958 38164 19010
rect 37212 18274 37268 18284
rect 38108 18338 38164 18958
rect 38108 18286 38110 18338
rect 38162 18286 38164 18338
rect 36428 16270 36430 16322
rect 36482 16270 36484 16322
rect 36428 16258 36484 16270
rect 37100 18116 37156 18126
rect 36428 13076 36484 13086
rect 36428 12982 36484 13020
rect 37100 13074 37156 18060
rect 37772 17892 37828 17902
rect 37772 17666 37828 17836
rect 37772 17614 37774 17666
rect 37826 17614 37828 17666
rect 37772 16322 37828 17614
rect 37772 16270 37774 16322
rect 37826 16270 37828 16322
rect 37772 16258 37828 16270
rect 37772 15988 37828 15998
rect 37548 15764 37604 15774
rect 37548 14532 37604 15708
rect 37772 15204 37828 15932
rect 37996 15874 38052 15886
rect 37996 15822 37998 15874
rect 38050 15822 38052 15874
rect 37884 15204 37940 15214
rect 37772 15202 37940 15204
rect 37772 15150 37886 15202
rect 37938 15150 37940 15202
rect 37772 15148 37940 15150
rect 37548 14530 37716 14532
rect 37548 14478 37550 14530
rect 37602 14478 37716 14530
rect 37548 14476 37716 14478
rect 37548 14466 37604 14476
rect 37212 14306 37268 14318
rect 37212 14254 37214 14306
rect 37266 14254 37268 14306
rect 37212 13860 37268 14254
rect 37212 13794 37268 13804
rect 37548 13860 37604 13870
rect 37548 13766 37604 13804
rect 37660 13522 37716 14476
rect 37660 13470 37662 13522
rect 37714 13470 37716 13522
rect 37660 13458 37716 13470
rect 37100 13022 37102 13074
rect 37154 13022 37156 13074
rect 37100 12852 37156 13022
rect 37100 12786 37156 12796
rect 36204 11666 36260 11676
rect 37660 11956 37716 11966
rect 35308 9548 35812 9604
rect 35868 9826 35924 9838
rect 35868 9774 35870 9826
rect 35922 9774 35924 9826
rect 35084 9044 35140 9054
rect 34636 7422 34638 7474
rect 34690 7422 34692 7474
rect 33628 6290 33684 6300
rect 32508 6130 32788 6132
rect 32508 6078 32510 6130
rect 32562 6078 32788 6130
rect 32508 6076 32788 6078
rect 32508 6066 32564 6076
rect 32172 5842 32228 5852
rect 32060 5234 32116 5628
rect 32060 5182 32062 5234
rect 32114 5182 32116 5234
rect 31612 5170 31668 5180
rect 32060 5124 32116 5182
rect 32732 5124 32788 6076
rect 33852 6018 33908 6524
rect 33852 5966 33854 6018
rect 33906 5966 33908 6018
rect 33852 5954 33908 5966
rect 33740 5684 33796 5694
rect 33516 5682 33796 5684
rect 33516 5630 33742 5682
rect 33794 5630 33796 5682
rect 33516 5628 33796 5630
rect 33516 5234 33572 5628
rect 33740 5618 33796 5628
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 34636 5236 34692 7422
rect 34972 8036 35028 8046
rect 34972 7252 35028 7980
rect 34972 7186 35028 7196
rect 35084 7474 35140 8988
rect 35308 9042 35364 9548
rect 35532 9156 35588 9166
rect 35532 9062 35588 9100
rect 35308 8990 35310 9042
rect 35362 8990 35364 9042
rect 35308 8978 35364 8990
rect 35868 9044 35924 9774
rect 36092 9828 36148 9838
rect 36092 9734 36148 9772
rect 37100 9828 37156 9838
rect 36540 9716 36596 9726
rect 36540 9622 36596 9660
rect 37100 9156 37156 9772
rect 37660 9826 37716 11900
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37660 9762 37716 9774
rect 37772 9714 37828 15148
rect 37884 15138 37940 15148
rect 37996 15148 38052 15822
rect 38108 15428 38164 18286
rect 38220 15538 38276 23100
rect 38444 23062 38500 23100
rect 38332 23042 38388 23054
rect 38332 22990 38334 23042
rect 38386 22990 38388 23042
rect 38332 21586 38388 22990
rect 38556 22370 38612 22382
rect 38556 22318 38558 22370
rect 38610 22318 38612 22370
rect 38444 22260 38500 22270
rect 38556 22260 38612 22318
rect 38500 22204 38612 22260
rect 38444 22194 38500 22204
rect 38332 21534 38334 21586
rect 38386 21534 38388 21586
rect 38332 21522 38388 21534
rect 38668 19908 38724 24558
rect 39228 23268 39284 23278
rect 39228 23174 39284 23212
rect 38780 23154 38836 23166
rect 38780 23102 38782 23154
rect 38834 23102 38836 23154
rect 38780 22484 38836 23102
rect 38780 22418 38836 22428
rect 38668 19842 38724 19852
rect 39004 21586 39060 21598
rect 39004 21534 39006 21586
rect 39058 21534 39060 21586
rect 38780 19796 38836 19806
rect 38780 19236 38836 19740
rect 38780 19142 38836 19180
rect 38332 19012 38388 19022
rect 38332 18918 38388 18956
rect 38892 19010 38948 19022
rect 38892 18958 38894 19010
rect 38946 18958 38948 19010
rect 38892 18900 38948 18958
rect 38668 18844 38948 18900
rect 38668 18676 38724 18844
rect 38444 18620 38724 18676
rect 38444 17668 38500 18620
rect 38556 18338 38612 18350
rect 38556 18286 38558 18338
rect 38610 18286 38612 18338
rect 38556 17892 38612 18286
rect 38556 17826 38612 17836
rect 38556 17668 38612 17678
rect 38444 17666 38612 17668
rect 38444 17614 38558 17666
rect 38610 17614 38612 17666
rect 38444 17612 38612 17614
rect 38556 17602 38612 17612
rect 38332 16324 38388 16334
rect 38332 16210 38388 16268
rect 38332 16158 38334 16210
rect 38386 16158 38388 16210
rect 38332 16146 38388 16158
rect 38220 15486 38222 15538
rect 38274 15486 38276 15538
rect 38220 15474 38276 15486
rect 38108 15362 38164 15372
rect 38556 15316 38612 15326
rect 38556 15222 38612 15260
rect 38780 15202 38836 15214
rect 38780 15150 38782 15202
rect 38834 15150 38836 15202
rect 38780 15148 38836 15150
rect 37996 15092 38612 15148
rect 38668 15092 38836 15148
rect 38556 15036 38724 15092
rect 38332 14756 38388 14766
rect 38332 14642 38388 14700
rect 38332 14590 38334 14642
rect 38386 14590 38388 14642
rect 38332 14578 38388 14590
rect 37884 14306 37940 14318
rect 37884 14254 37886 14306
rect 37938 14254 37940 14306
rect 37884 13860 37940 14254
rect 37884 13794 37940 13804
rect 38444 13860 38500 13870
rect 38444 13766 38500 13804
rect 38108 13634 38164 13646
rect 38108 13582 38110 13634
rect 38162 13582 38164 13634
rect 38108 13522 38164 13582
rect 38108 13470 38110 13522
rect 38162 13470 38164 13522
rect 38108 13458 38164 13470
rect 38108 12066 38164 12078
rect 38108 12014 38110 12066
rect 38162 12014 38164 12066
rect 38108 11956 38164 12014
rect 38108 11890 38164 11900
rect 37884 11620 37940 11630
rect 38556 11620 38612 15036
rect 39004 14306 39060 21534
rect 39116 19348 39172 19358
rect 39116 19234 39172 19292
rect 39788 19348 39844 19358
rect 39788 19254 39844 19292
rect 39116 19182 39118 19234
rect 39170 19182 39172 19234
rect 39116 19170 39172 19182
rect 39340 19124 39396 19134
rect 39340 19122 39732 19124
rect 39340 19070 39342 19122
rect 39394 19070 39732 19122
rect 39340 19068 39732 19070
rect 39340 19058 39396 19068
rect 39564 18788 39620 18798
rect 39564 18674 39620 18732
rect 39564 18622 39566 18674
rect 39618 18622 39620 18674
rect 39564 18610 39620 18622
rect 39676 18674 39732 19068
rect 39676 18622 39678 18674
rect 39730 18622 39732 18674
rect 39676 18610 39732 18622
rect 39788 18562 39844 18574
rect 39788 18510 39790 18562
rect 39842 18510 39844 18562
rect 39788 17780 39844 18510
rect 39900 18004 39956 25452
rect 40012 22260 40068 25564
rect 40124 25508 40180 25518
rect 40124 25414 40180 25452
rect 40236 25394 40292 25406
rect 40236 25342 40238 25394
rect 40290 25342 40292 25394
rect 40236 24052 40292 25342
rect 40236 23986 40292 23996
rect 40012 22204 40292 22260
rect 40236 21812 40292 22204
rect 40348 21812 40404 21822
rect 40236 21810 40404 21812
rect 40236 21758 40350 21810
rect 40402 21758 40404 21810
rect 40236 21756 40404 21758
rect 40348 21588 40404 21756
rect 40348 21522 40404 21532
rect 40460 20244 40516 38612
rect 41580 38050 41636 38062
rect 41580 37998 41582 38050
rect 41634 37998 41636 38050
rect 40796 37826 40852 37838
rect 40796 37774 40798 37826
rect 40850 37774 40852 37826
rect 40796 36708 40852 37774
rect 40908 37156 40964 37166
rect 40908 37062 40964 37100
rect 41244 37156 41300 37166
rect 40908 36708 40964 36718
rect 40796 36706 40964 36708
rect 40796 36654 40910 36706
rect 40962 36654 40964 36706
rect 40796 36652 40964 36654
rect 40908 36642 40964 36652
rect 41244 36706 41300 37100
rect 41244 36654 41246 36706
rect 41298 36654 41300 36706
rect 41244 36642 41300 36654
rect 41132 36260 41188 36270
rect 41580 36260 41636 37998
rect 41692 36260 41748 36270
rect 41132 36258 41748 36260
rect 41132 36206 41134 36258
rect 41186 36206 41694 36258
rect 41746 36206 41748 36258
rect 41132 36204 41748 36206
rect 41132 34356 41188 36204
rect 41692 36194 41748 36204
rect 40796 34300 41188 34356
rect 41468 34356 41524 34366
rect 40684 26292 40740 26302
rect 40684 25730 40740 26236
rect 40684 25678 40686 25730
rect 40738 25678 40740 25730
rect 40684 25666 40740 25678
rect 40684 25508 40740 25518
rect 40572 25396 40628 25406
rect 40572 25302 40628 25340
rect 40684 25394 40740 25452
rect 40684 25342 40686 25394
rect 40738 25342 40740 25394
rect 40684 25330 40740 25342
rect 40796 23548 40852 34300
rect 41468 34262 41524 34300
rect 41020 34132 41076 34142
rect 41020 34038 41076 34076
rect 41244 34132 41300 34142
rect 41244 33348 41300 34076
rect 41692 34130 41748 34142
rect 41692 34078 41694 34130
rect 41746 34078 41748 34130
rect 41580 34018 41636 34030
rect 41580 33966 41582 34018
rect 41634 33966 41636 34018
rect 41580 33348 41636 33966
rect 41692 33572 41748 34078
rect 41692 33506 41748 33516
rect 41692 33348 41748 33358
rect 41244 33346 41524 33348
rect 41244 33294 41246 33346
rect 41298 33294 41524 33346
rect 41244 33292 41524 33294
rect 41580 33346 41748 33348
rect 41580 33294 41694 33346
rect 41746 33294 41748 33346
rect 41580 33292 41748 33294
rect 41244 33282 41300 33292
rect 41468 33124 41524 33292
rect 41692 33282 41748 33292
rect 41468 33068 41748 33124
rect 41692 31890 41748 33068
rect 41692 31838 41694 31890
rect 41746 31838 41748 31890
rect 41692 31826 41748 31838
rect 41804 31668 41860 40684
rect 43372 40516 43428 40526
rect 43372 40292 43428 40460
rect 43596 40292 43652 40302
rect 43372 40290 43652 40292
rect 43372 40238 43598 40290
rect 43650 40238 43652 40290
rect 43372 40236 43652 40238
rect 43372 39730 43428 40236
rect 43596 40226 43652 40236
rect 43372 39678 43374 39730
rect 43426 39678 43428 39730
rect 43372 39666 43428 39678
rect 42252 39394 42308 39406
rect 42252 39342 42254 39394
rect 42306 39342 42308 39394
rect 42252 39284 42308 39342
rect 42140 39228 42252 39284
rect 42140 38050 42196 39228
rect 42252 39218 42308 39228
rect 42140 37998 42142 38050
rect 42194 37998 42196 38050
rect 42140 37986 42196 37998
rect 43036 37156 43092 37166
rect 43036 37062 43092 37100
rect 42476 35700 42532 35710
rect 42364 34804 42420 34814
rect 42364 34356 42420 34748
rect 42140 34300 42364 34356
rect 42028 34132 42084 34142
rect 42028 34038 42084 34076
rect 41244 31612 41860 31668
rect 41916 34020 41972 34030
rect 41132 27860 41188 27870
rect 41132 27766 41188 27804
rect 40908 27076 40964 27086
rect 40908 26982 40964 27020
rect 41132 26292 41188 26302
rect 40908 26236 41132 26292
rect 40908 24834 40964 26236
rect 41132 26198 41188 26236
rect 41020 26068 41076 26078
rect 41020 25974 41076 26012
rect 40908 24782 40910 24834
rect 40962 24782 40964 24834
rect 40908 24770 40964 24782
rect 41132 24836 41188 24846
rect 41132 24742 41188 24780
rect 41244 24724 41300 31612
rect 41916 31556 41972 33964
rect 42028 33348 42084 33358
rect 42140 33348 42196 34300
rect 42364 34262 42420 34300
rect 42028 33346 42196 33348
rect 42028 33294 42030 33346
rect 42082 33294 42196 33346
rect 42028 33292 42196 33294
rect 42364 33572 42420 33582
rect 42364 33346 42420 33516
rect 42364 33294 42366 33346
rect 42418 33294 42420 33346
rect 42028 33282 42084 33292
rect 42364 33236 42420 33294
rect 42364 33170 42420 33180
rect 42028 33122 42084 33134
rect 42028 33070 42030 33122
rect 42082 33070 42084 33122
rect 42028 32340 42084 33070
rect 42028 32274 42084 32284
rect 42476 31948 42532 35644
rect 42700 35586 42756 35598
rect 42700 35534 42702 35586
rect 42754 35534 42756 35586
rect 42700 34468 42756 35534
rect 43708 35028 43764 42476
rect 43820 41970 43876 42588
rect 43932 42578 43988 42588
rect 43820 41918 43822 41970
rect 43874 41918 43876 41970
rect 43820 41906 43876 41918
rect 43932 42420 43988 42430
rect 43820 41748 43876 41758
rect 43932 41748 43988 42364
rect 44268 41972 44324 43932
rect 45388 43538 45444 43550
rect 45388 43486 45390 43538
rect 45442 43486 45444 43538
rect 44940 43428 44996 43438
rect 45388 43428 45444 43486
rect 44996 43372 45108 43428
rect 44940 43334 44996 43372
rect 43820 41746 43988 41748
rect 43820 41694 43822 41746
rect 43874 41694 43988 41746
rect 43820 41692 43988 41694
rect 44044 41916 44324 41972
rect 43820 41682 43876 41692
rect 44044 40514 44100 41916
rect 44492 41858 44548 41870
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 44156 41410 44212 41422
rect 44156 41358 44158 41410
rect 44210 41358 44212 41410
rect 44156 41300 44212 41358
rect 44268 41300 44324 41310
rect 44156 41244 44268 41300
rect 44268 41234 44324 41244
rect 44268 41074 44324 41086
rect 44268 41022 44270 41074
rect 44322 41022 44324 41074
rect 44156 40964 44212 40974
rect 44156 40870 44212 40908
rect 44044 40462 44046 40514
rect 44098 40462 44100 40514
rect 44044 40450 44100 40462
rect 43820 40402 43876 40414
rect 43820 40350 43822 40402
rect 43874 40350 43876 40402
rect 43820 39620 43876 40350
rect 44268 40404 44324 41022
rect 44492 40964 44548 41806
rect 44492 40898 44548 40908
rect 44604 40404 44660 40414
rect 45052 40404 45108 43372
rect 45388 43362 45444 43372
rect 45164 42532 45220 42542
rect 45164 42438 45220 42476
rect 45500 42420 45556 44382
rect 45612 44322 45668 44334
rect 45612 44270 45614 44322
rect 45666 44270 45668 44322
rect 45612 42980 45668 44270
rect 45612 42886 45668 42924
rect 45612 42756 45668 42766
rect 45612 42642 45668 42700
rect 45612 42590 45614 42642
rect 45666 42590 45668 42642
rect 45612 42578 45668 42590
rect 45724 42642 45780 42654
rect 45724 42590 45726 42642
rect 45778 42590 45780 42642
rect 45500 42354 45556 42364
rect 45724 41972 45780 42590
rect 45948 42532 46004 45612
rect 46956 44548 47012 50318
rect 47068 50370 47124 50382
rect 47516 50372 47908 50428
rect 47068 50318 47070 50370
rect 47122 50318 47124 50370
rect 47068 50036 47124 50318
rect 47068 49980 47348 50036
rect 47292 49922 47348 49980
rect 47292 49870 47294 49922
rect 47346 49870 47348 49922
rect 47292 49858 47348 49870
rect 47404 49588 47460 49598
rect 47404 49494 47460 49532
rect 47740 47570 47796 47582
rect 47740 47518 47742 47570
rect 47794 47518 47796 47570
rect 47740 47236 47796 47518
rect 47740 47170 47796 47180
rect 48524 47234 48580 47246
rect 48524 47182 48526 47234
rect 48578 47182 48580 47234
rect 48076 46676 48132 46686
rect 48524 46676 48580 47182
rect 48076 46674 48580 46676
rect 48076 46622 48078 46674
rect 48130 46622 48580 46674
rect 48076 46620 48580 46622
rect 47628 46562 47684 46574
rect 47628 46510 47630 46562
rect 47682 46510 47684 46562
rect 47628 46452 47684 46510
rect 47628 46386 47684 46396
rect 48076 45668 48132 46620
rect 48412 45892 48468 45902
rect 48412 45798 48468 45836
rect 48132 45612 48356 45668
rect 48076 45574 48132 45612
rect 48300 45332 48356 45612
rect 48300 45238 48356 45276
rect 46508 44492 47124 44548
rect 46508 44322 46564 44492
rect 46508 44270 46510 44322
rect 46562 44270 46564 44322
rect 46508 44258 46564 44270
rect 46732 44380 47012 44436
rect 46620 44098 46676 44110
rect 46620 44046 46622 44098
rect 46674 44046 46676 44098
rect 46620 43708 46676 44046
rect 46060 43652 46676 43708
rect 46060 43650 46116 43652
rect 46060 43598 46062 43650
rect 46114 43598 46116 43650
rect 46060 43586 46116 43598
rect 46620 43428 46676 43438
rect 46620 42756 46676 43372
rect 46732 42866 46788 44380
rect 46956 44322 47012 44380
rect 46956 44270 46958 44322
rect 47010 44270 47012 44322
rect 46956 44258 47012 44270
rect 46844 44210 46900 44222
rect 46844 44158 46846 44210
rect 46898 44158 46900 44210
rect 46844 43428 46900 44158
rect 47068 44100 47124 44492
rect 46844 43362 46900 43372
rect 46956 44044 47124 44100
rect 46732 42814 46734 42866
rect 46786 42814 46788 42866
rect 46732 42802 46788 42814
rect 46620 42662 46676 42700
rect 45948 42466 46004 42476
rect 46396 42532 46452 42542
rect 46396 42438 46452 42476
rect 46844 42532 46900 42542
rect 46956 42532 47012 44044
rect 48188 43428 48244 43438
rect 48188 43334 48244 43372
rect 46844 42530 47012 42532
rect 46844 42478 46846 42530
rect 46898 42478 47012 42530
rect 46844 42476 47012 42478
rect 45724 41906 45780 41916
rect 46844 41972 46900 42476
rect 46844 41906 46900 41916
rect 45164 41300 45220 41310
rect 45164 41206 45220 41244
rect 45500 41300 45556 41310
rect 45500 41298 45892 41300
rect 45500 41246 45502 41298
rect 45554 41246 45892 41298
rect 45500 41244 45892 41246
rect 45500 41234 45556 41244
rect 44268 40402 44660 40404
rect 44268 40350 44606 40402
rect 44658 40350 44660 40402
rect 44268 40348 44660 40350
rect 44604 39844 44660 40348
rect 44604 39778 44660 39788
rect 44716 40402 45108 40404
rect 44716 40350 45054 40402
rect 45106 40350 45108 40402
rect 44716 40348 45108 40350
rect 43820 39526 43876 39564
rect 44268 39508 44324 39518
rect 44268 39414 44324 39452
rect 44716 39060 44772 40348
rect 45052 40338 45108 40348
rect 45164 40964 45220 40974
rect 45388 40964 45444 40974
rect 45164 40068 45220 40908
rect 44268 39058 44772 39060
rect 44268 39006 44718 39058
rect 44770 39006 44772 39058
rect 44268 39004 44772 39006
rect 44268 37492 44324 39004
rect 44716 38994 44772 39004
rect 44940 40012 45220 40068
rect 45276 40962 45444 40964
rect 45276 40910 45390 40962
rect 45442 40910 45444 40962
rect 45276 40908 45444 40910
rect 44940 38668 44996 40012
rect 45276 39730 45332 40908
rect 45388 40898 45444 40908
rect 45836 40514 45892 41244
rect 48636 41298 48692 59164
rect 48860 58772 48916 59390
rect 48972 59444 49028 59454
rect 49084 59444 49140 60956
rect 49644 61010 49700 61404
rect 49644 60958 49646 61010
rect 49698 60958 49700 61010
rect 49644 60946 49700 60958
rect 49756 61012 49812 61022
rect 48972 59442 49140 59444
rect 48972 59390 48974 59442
rect 49026 59390 49140 59442
rect 48972 59388 49140 59390
rect 49308 60786 49364 60798
rect 49308 60734 49310 60786
rect 49362 60734 49364 60786
rect 48972 59378 49028 59388
rect 48860 58706 48916 58716
rect 49308 59218 49364 60734
rect 49644 60786 49700 60798
rect 49644 60734 49646 60786
rect 49698 60734 49700 60786
rect 49532 60676 49588 60686
rect 49532 60004 49588 60620
rect 49644 60228 49700 60734
rect 49756 60676 49812 60956
rect 50092 60786 50148 62188
rect 50428 63810 50484 63822
rect 50428 63758 50430 63810
rect 50482 63758 50484 63810
rect 50428 61012 50484 63758
rect 50764 63810 50820 63980
rect 50876 63970 50932 63980
rect 50764 63758 50766 63810
rect 50818 63758 50820 63810
rect 50764 63746 50820 63758
rect 50652 63476 50708 63486
rect 50652 63138 50708 63420
rect 50652 63086 50654 63138
rect 50706 63086 50708 63138
rect 50652 63074 50708 63086
rect 50764 63140 50820 63150
rect 50764 63046 50820 63084
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50988 61908 51044 64204
rect 51324 64148 51380 65324
rect 51660 65314 51716 65324
rect 51772 65380 51828 65390
rect 51772 64930 51828 65324
rect 51772 64878 51774 64930
rect 51826 64878 51828 64930
rect 51772 64866 51828 64878
rect 51996 65378 52052 65390
rect 51996 65326 51998 65378
rect 52050 65326 52052 65378
rect 51212 64092 51380 64148
rect 51660 64594 51716 64606
rect 51660 64542 51662 64594
rect 51714 64542 51716 64594
rect 51212 64034 51268 64092
rect 51212 63982 51214 64034
rect 51266 63982 51268 64034
rect 50988 61842 51044 61852
rect 51100 63252 51156 63262
rect 51100 63138 51156 63196
rect 51100 63086 51102 63138
rect 51154 63086 51156 63138
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50428 60946 50484 60956
rect 50988 61012 51044 61022
rect 50988 60918 51044 60956
rect 50092 60734 50094 60786
rect 50146 60734 50148 60786
rect 50092 60722 50148 60734
rect 50204 60900 50260 60910
rect 49756 60582 49812 60620
rect 49644 60172 49924 60228
rect 49868 60114 49924 60172
rect 49868 60062 49870 60114
rect 49922 60062 49924 60114
rect 49532 59948 49700 60004
rect 49532 59442 49588 59454
rect 49532 59390 49534 59442
rect 49586 59390 49588 59442
rect 49532 59332 49588 59390
rect 49532 59266 49588 59276
rect 49308 59166 49310 59218
rect 49362 59166 49364 59218
rect 49196 56756 49252 56766
rect 48860 56754 49252 56756
rect 48860 56702 49198 56754
rect 49250 56702 49252 56754
rect 48860 56700 49252 56702
rect 48860 56306 48916 56700
rect 49196 56690 49252 56700
rect 48860 56254 48862 56306
rect 48914 56254 48916 56306
rect 48860 56242 48916 56254
rect 48748 56196 48804 56206
rect 48748 56102 48804 56140
rect 49308 55188 49364 59166
rect 49420 59218 49476 59230
rect 49420 59166 49422 59218
rect 49474 59166 49476 59218
rect 49420 57428 49476 59166
rect 49644 59106 49700 59948
rect 49868 59220 49924 60062
rect 50204 59890 50260 60844
rect 50988 60676 51044 60686
rect 50988 60002 51044 60620
rect 50988 59950 50990 60002
rect 51042 59950 51044 60002
rect 50988 59938 51044 59950
rect 51100 60004 51156 63086
rect 51212 63138 51268 63982
rect 51324 63924 51380 63934
rect 51324 63830 51380 63868
rect 51212 63086 51214 63138
rect 51266 63086 51268 63138
rect 51212 63074 51268 63086
rect 51436 63250 51492 63262
rect 51436 63198 51438 63250
rect 51490 63198 51492 63250
rect 51436 61012 51492 63198
rect 51660 63250 51716 64542
rect 51660 63198 51662 63250
rect 51714 63198 51716 63250
rect 51660 63186 51716 63198
rect 51772 63140 51828 63150
rect 51996 63140 52052 65326
rect 51772 63138 52052 63140
rect 51772 63086 51774 63138
rect 51826 63086 52052 63138
rect 51772 63084 52052 63086
rect 52108 64484 52164 64494
rect 51660 62244 51716 62254
rect 51660 62150 51716 62188
rect 51436 60946 51492 60956
rect 51212 60786 51268 60798
rect 51660 60788 51716 60798
rect 51212 60734 51214 60786
rect 51266 60734 51268 60786
rect 51212 60228 51268 60734
rect 51212 60162 51268 60172
rect 51548 60732 51660 60788
rect 51212 60004 51268 60014
rect 51100 60002 51268 60004
rect 51100 59950 51214 60002
rect 51266 59950 51268 60002
rect 51100 59948 51268 59950
rect 50204 59838 50206 59890
rect 50258 59838 50260 59890
rect 50204 59826 50260 59838
rect 50540 59780 50596 59790
rect 50540 59778 50932 59780
rect 50540 59726 50542 59778
rect 50594 59726 50932 59778
rect 50540 59724 50932 59726
rect 50540 59714 50596 59724
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50876 59556 50932 59724
rect 51100 59778 51156 59790
rect 51100 59726 51102 59778
rect 51154 59726 51156 59778
rect 51100 59556 51156 59726
rect 50876 59500 51156 59556
rect 50428 59444 50484 59454
rect 49980 59220 50036 59230
rect 49868 59218 50036 59220
rect 49868 59166 49982 59218
rect 50034 59166 50036 59218
rect 49868 59164 50036 59166
rect 49980 59154 50036 59164
rect 49644 59054 49646 59106
rect 49698 59054 49700 59106
rect 49644 59042 49700 59054
rect 49420 57362 49476 57372
rect 50428 56980 50484 59388
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50316 56978 50484 56980
rect 50316 56926 50430 56978
rect 50482 56926 50484 56978
rect 50316 56924 50484 56926
rect 49980 56868 50036 56878
rect 50316 56868 50372 56924
rect 50428 56914 50484 56924
rect 49980 56866 50372 56868
rect 49980 56814 49982 56866
rect 50034 56814 50372 56866
rect 49980 56812 50372 56814
rect 49980 56802 50036 56812
rect 49980 56308 50036 56318
rect 49980 56214 50036 56252
rect 50316 56308 50372 56812
rect 50988 56756 51044 59500
rect 50316 56242 50372 56252
rect 50428 56700 51044 56756
rect 51100 57540 51156 57550
rect 50316 56084 50372 56094
rect 50316 55990 50372 56028
rect 49308 55122 49364 55132
rect 49980 55188 50036 55198
rect 49980 55094 50036 55132
rect 49196 55074 49252 55086
rect 49196 55022 49198 55074
rect 49250 55022 49252 55074
rect 49196 54628 49252 55022
rect 49532 55076 49588 55086
rect 49532 54982 49588 55020
rect 50316 55074 50372 55086
rect 50316 55022 50318 55074
rect 50370 55022 50372 55074
rect 49196 54562 49252 54572
rect 50316 54516 50372 55022
rect 50316 54450 50372 54460
rect 50428 55076 50484 56700
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50876 56308 50932 56318
rect 50876 56082 50932 56252
rect 50876 56030 50878 56082
rect 50930 56030 50932 56082
rect 50876 55468 50932 56030
rect 50876 55412 51044 55468
rect 49756 52052 49812 52062
rect 48860 52050 49812 52052
rect 48860 51998 49758 52050
rect 49810 51998 49812 52050
rect 48860 51996 49812 51998
rect 48748 51604 48804 51614
rect 48748 51490 48804 51548
rect 48860 51602 48916 51996
rect 49756 51986 49812 51996
rect 50428 51940 50484 55020
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50876 54516 50932 54526
rect 50876 54422 50932 54460
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50988 53060 51044 55412
rect 50764 53004 50988 53060
rect 51100 53060 51156 57484
rect 51212 54626 51268 59948
rect 51436 59444 51492 59454
rect 51436 59218 51492 59388
rect 51436 59166 51438 59218
rect 51490 59166 51492 59218
rect 51436 59154 51492 59166
rect 51548 57876 51604 60732
rect 51660 60722 51716 60732
rect 51660 60004 51716 60014
rect 51772 60004 51828 63084
rect 52108 62580 52164 64428
rect 52332 64146 52388 65436
rect 54908 65490 54964 65502
rect 54908 65438 54910 65490
rect 54962 65438 54964 65490
rect 54124 65380 54180 65390
rect 54124 65286 54180 65324
rect 54908 65380 54964 65438
rect 54908 64818 54964 65324
rect 54908 64766 54910 64818
rect 54962 64766 54964 64818
rect 52780 64484 52836 64494
rect 52780 64390 52836 64428
rect 54908 64484 54964 64766
rect 52332 64094 52334 64146
rect 52386 64094 52388 64146
rect 52332 64082 52388 64094
rect 54236 64148 54292 64158
rect 54124 63924 54180 63934
rect 53564 63922 54180 63924
rect 53564 63870 54126 63922
rect 54178 63870 54180 63922
rect 53564 63868 54180 63870
rect 53564 63362 53620 63868
rect 54124 63858 54180 63868
rect 53564 63310 53566 63362
rect 53618 63310 53620 63362
rect 53564 63298 53620 63310
rect 53004 63252 53060 63262
rect 53900 63252 53956 63262
rect 53060 63196 53172 63252
rect 53004 63158 53060 63196
rect 52108 62486 52164 62524
rect 52444 62468 52500 62478
rect 52444 62374 52500 62412
rect 52892 62244 52948 62254
rect 52780 61684 52836 61694
rect 52892 61684 52948 62188
rect 52780 61682 52948 61684
rect 52780 61630 52782 61682
rect 52834 61630 52948 61682
rect 52780 61628 52948 61630
rect 52780 60676 52836 61628
rect 53116 61570 53172 63196
rect 53900 63158 53956 63196
rect 53228 63138 53284 63150
rect 53228 63086 53230 63138
rect 53282 63086 53284 63138
rect 53228 62468 53284 63086
rect 53228 62402 53284 62412
rect 54124 63138 54180 63150
rect 54124 63086 54126 63138
rect 54178 63086 54180 63138
rect 53116 61518 53118 61570
rect 53170 61518 53172 61570
rect 53116 61506 53172 61518
rect 53452 62354 53508 62366
rect 53452 62302 53454 62354
rect 53506 62302 53508 62354
rect 53004 60788 53060 60798
rect 53004 60694 53060 60732
rect 52780 60610 52836 60620
rect 53340 60676 53396 60686
rect 53452 60676 53508 62302
rect 54124 62244 54180 63086
rect 54124 62178 54180 62188
rect 54236 61570 54292 64092
rect 54572 64148 54628 64158
rect 54572 64054 54628 64092
rect 54796 63922 54852 63934
rect 54796 63870 54798 63922
rect 54850 63870 54852 63922
rect 54684 63810 54740 63822
rect 54684 63758 54686 63810
rect 54738 63758 54740 63810
rect 54684 63588 54740 63758
rect 54236 61518 54238 61570
rect 54290 61518 54292 61570
rect 54236 61506 54292 61518
rect 54348 63532 54740 63588
rect 54348 60900 54404 63532
rect 54460 63364 54516 63374
rect 54796 63364 54852 63870
rect 54460 63362 54852 63364
rect 54460 63310 54462 63362
rect 54514 63310 54852 63362
rect 54460 63308 54852 63310
rect 54460 63298 54516 63308
rect 54908 63250 54964 64428
rect 55020 63476 55076 66222
rect 55132 63812 55188 69200
rect 56028 66500 56084 66510
rect 56028 66406 56084 66444
rect 55468 65380 55524 65390
rect 55468 65286 55524 65324
rect 55356 65156 55412 65166
rect 55244 64932 55300 64942
rect 55244 64818 55300 64876
rect 55244 64766 55246 64818
rect 55298 64766 55300 64818
rect 55244 64754 55300 64766
rect 55244 64036 55300 64046
rect 55244 63942 55300 63980
rect 55132 63746 55188 63756
rect 55020 63410 55076 63420
rect 54908 63198 54910 63250
rect 54962 63198 54964 63250
rect 54348 60834 54404 60844
rect 54460 61012 54516 61022
rect 54460 60898 54516 60956
rect 54460 60846 54462 60898
rect 54514 60846 54516 60898
rect 54460 60834 54516 60846
rect 53340 60674 53508 60676
rect 53340 60622 53342 60674
rect 53394 60622 53508 60674
rect 53340 60620 53508 60622
rect 54684 60786 54740 60798
rect 54684 60734 54686 60786
rect 54738 60734 54740 60786
rect 53340 60564 53396 60620
rect 53340 60498 53396 60508
rect 54684 60564 54740 60734
rect 54684 60498 54740 60508
rect 51660 60002 51828 60004
rect 51660 59950 51662 60002
rect 51714 59950 51828 60002
rect 51660 59948 51828 59950
rect 51884 60228 51940 60238
rect 51884 60002 51940 60172
rect 54908 60114 54964 63198
rect 55244 63252 55300 63262
rect 55244 63158 55300 63196
rect 55020 62580 55076 62590
rect 55020 61682 55076 62524
rect 55356 62242 55412 65100
rect 57148 65156 57204 69200
rect 58156 66164 58212 66174
rect 57820 65602 57876 65614
rect 57820 65550 57822 65602
rect 57874 65550 57876 65602
rect 57596 65492 57652 65502
rect 57596 65398 57652 65436
rect 57148 65090 57204 65100
rect 57372 64596 57428 64606
rect 57260 64594 57428 64596
rect 57260 64542 57374 64594
rect 57426 64542 57428 64594
rect 57260 64540 57428 64542
rect 55804 64036 55860 64046
rect 55692 63980 55804 64036
rect 55580 63698 55636 63710
rect 55580 63646 55582 63698
rect 55634 63646 55636 63698
rect 55580 62580 55636 63646
rect 55580 62514 55636 62524
rect 55356 62190 55358 62242
rect 55410 62190 55412 62242
rect 55356 62178 55412 62190
rect 55020 61630 55022 61682
rect 55074 61630 55076 61682
rect 55020 61618 55076 61630
rect 55468 61572 55524 61582
rect 55468 61478 55524 61516
rect 54908 60062 54910 60114
rect 54962 60062 54964 60114
rect 51884 59950 51886 60002
rect 51938 59950 51940 60002
rect 51660 59938 51716 59948
rect 51660 57876 51716 57886
rect 51548 57874 51716 57876
rect 51548 57822 51662 57874
rect 51714 57822 51716 57874
rect 51548 57820 51716 57822
rect 51660 57810 51716 57820
rect 51436 57652 51492 57662
rect 51436 57558 51492 57596
rect 51548 57538 51604 57550
rect 51548 57486 51550 57538
rect 51602 57486 51604 57538
rect 51548 56196 51604 57486
rect 51660 56196 51716 56206
rect 51548 56194 51716 56196
rect 51548 56142 51662 56194
rect 51714 56142 51716 56194
rect 51548 56140 51716 56142
rect 51660 56130 51716 56140
rect 51436 56084 51492 56094
rect 51212 54574 51214 54626
rect 51266 54574 51268 54626
rect 51212 53396 51268 54574
rect 51324 54740 51380 54750
rect 51324 53508 51380 54684
rect 51436 53732 51492 56028
rect 51884 56084 51940 59950
rect 52108 60004 52164 60014
rect 52108 59910 52164 59948
rect 53340 60004 53396 60014
rect 51996 59778 52052 59790
rect 51996 59726 51998 59778
rect 52050 59726 52052 59778
rect 51996 58546 52052 59726
rect 52108 59106 52164 59118
rect 52108 59054 52110 59106
rect 52162 59054 52164 59106
rect 52108 58658 52164 59054
rect 52108 58606 52110 58658
rect 52162 58606 52164 58658
rect 52108 58594 52164 58606
rect 51996 58494 51998 58546
rect 52050 58494 52052 58546
rect 51996 58482 52052 58494
rect 53004 58434 53060 58446
rect 53004 58382 53006 58434
rect 53058 58382 53060 58434
rect 52556 58324 52612 58334
rect 52556 57874 52612 58268
rect 53004 58324 53060 58382
rect 53004 58258 53060 58268
rect 52556 57822 52558 57874
rect 52610 57822 52612 57874
rect 52556 57810 52612 57822
rect 51996 57650 52052 57662
rect 51996 57598 51998 57650
rect 52050 57598 52052 57650
rect 51996 56532 52052 57598
rect 51996 56466 52052 56476
rect 52780 56532 52836 56542
rect 51884 56018 51940 56028
rect 52780 55410 52836 56476
rect 52780 55358 52782 55410
rect 52834 55358 52836 55410
rect 52780 55346 52836 55358
rect 53340 55298 53396 59948
rect 54236 60004 54292 60014
rect 54908 60004 54964 60062
rect 55244 61012 55300 61022
rect 55244 60114 55300 60956
rect 55244 60062 55246 60114
rect 55298 60062 55300 60114
rect 55244 60050 55300 60062
rect 54236 59106 54292 59948
rect 54236 59054 54238 59106
rect 54290 59054 54292 59106
rect 54236 59042 54292 59054
rect 54684 59948 54908 60004
rect 54684 59444 54740 59948
rect 54908 59938 54964 59948
rect 54684 58548 54740 59388
rect 55692 59444 55748 63980
rect 55804 63942 55860 63980
rect 56364 63812 56420 63822
rect 57260 63812 57316 64540
rect 57372 64530 57428 64540
rect 55916 63700 55972 63710
rect 55916 63606 55972 63644
rect 56364 61794 56420 63756
rect 57036 63756 57316 63812
rect 56588 62636 56868 62692
rect 56588 62466 56644 62636
rect 56588 62414 56590 62466
rect 56642 62414 56644 62466
rect 56588 62402 56644 62414
rect 56700 62466 56756 62478
rect 56700 62414 56702 62466
rect 56754 62414 56756 62466
rect 56364 61742 56366 61794
rect 56418 61742 56420 61794
rect 56364 61730 56420 61742
rect 56700 61012 56756 62414
rect 56700 60946 56756 60956
rect 55804 60900 55860 60910
rect 55804 60806 55860 60844
rect 56588 60900 56644 60910
rect 56588 60806 56644 60844
rect 56028 60676 56084 60686
rect 56028 60674 56644 60676
rect 56028 60622 56030 60674
rect 56082 60622 56644 60674
rect 56028 60620 56644 60622
rect 56028 60610 56084 60620
rect 56028 59444 56084 59454
rect 55692 59442 56084 59444
rect 55692 59390 56030 59442
rect 56082 59390 56084 59442
rect 55692 59388 56084 59390
rect 55692 59220 55748 59388
rect 56028 59378 56084 59388
rect 56588 59330 56644 60620
rect 56700 60564 56756 60574
rect 56812 60564 56868 62636
rect 56924 62354 56980 62366
rect 56924 62302 56926 62354
rect 56978 62302 56980 62354
rect 56924 60786 56980 62302
rect 57036 61010 57092 63756
rect 57372 63700 57428 63710
rect 57372 63250 57428 63644
rect 57372 63198 57374 63250
rect 57426 63198 57428 63250
rect 57372 63186 57428 63198
rect 57036 60958 57038 61010
rect 57090 60958 57092 61010
rect 57036 60946 57092 60958
rect 57260 62242 57316 62254
rect 57260 62190 57262 62242
rect 57314 62190 57316 62242
rect 56924 60734 56926 60786
rect 56978 60734 56980 60786
rect 56924 60722 56980 60734
rect 57260 60786 57316 62190
rect 57820 61012 57876 65550
rect 58156 65492 58212 66108
rect 58156 65398 58212 65436
rect 58156 64706 58212 64718
rect 58156 64654 58158 64706
rect 58210 64654 58212 64706
rect 58156 63138 58212 64654
rect 58156 63086 58158 63138
rect 58210 63086 58212 63138
rect 57260 60734 57262 60786
rect 57314 60734 57316 60786
rect 56756 60508 56868 60564
rect 57148 60676 57204 60686
rect 57148 60562 57204 60620
rect 57148 60510 57150 60562
rect 57202 60510 57204 60562
rect 56700 60498 56756 60508
rect 57148 60498 57204 60510
rect 56700 59444 56756 59454
rect 56700 59350 56756 59388
rect 56588 59278 56590 59330
rect 56642 59278 56644 59330
rect 56588 59266 56644 59278
rect 56812 59330 56868 59342
rect 56812 59278 56814 59330
rect 56866 59278 56868 59330
rect 55692 59154 55748 59164
rect 56812 59220 56868 59278
rect 56812 59154 56868 59164
rect 54236 58546 54740 58548
rect 54236 58494 54686 58546
rect 54738 58494 54740 58546
rect 54236 58492 54740 58494
rect 54236 56308 54292 58492
rect 54684 58482 54740 58492
rect 55356 56980 55412 56990
rect 53900 56306 54292 56308
rect 53900 56254 54238 56306
rect 54290 56254 54292 56306
rect 53900 56252 54292 56254
rect 53340 55246 53342 55298
rect 53394 55246 53396 55298
rect 53340 55234 53396 55246
rect 53788 55970 53844 55982
rect 53788 55918 53790 55970
rect 53842 55918 53844 55970
rect 52780 55074 52836 55086
rect 52780 55022 52782 55074
rect 52834 55022 52836 55074
rect 51884 54740 51940 54750
rect 51884 54646 51940 54684
rect 51660 54516 51716 54526
rect 51660 53956 51716 54460
rect 51660 53890 51716 53900
rect 52668 53956 52724 53966
rect 52668 53862 52724 53900
rect 52780 53844 52836 55022
rect 52892 55076 52948 55086
rect 52892 54982 52948 55020
rect 53116 55074 53172 55086
rect 53116 55022 53118 55074
rect 53170 55022 53172 55074
rect 53116 54740 53172 55022
rect 53116 54674 53172 54684
rect 53788 55076 53844 55918
rect 53004 53844 53060 53854
rect 52780 53778 52836 53788
rect 52892 53788 53004 53844
rect 51436 53730 51940 53732
rect 51436 53678 51438 53730
rect 51490 53678 51940 53730
rect 51436 53676 51940 53678
rect 51436 53666 51492 53676
rect 51660 53508 51716 53518
rect 51324 53452 51604 53508
rect 51212 53340 51380 53396
rect 51100 53004 51268 53060
rect 50764 52948 50820 53004
rect 50988 52966 51044 53004
rect 50540 52946 50820 52948
rect 50540 52894 50766 52946
rect 50818 52894 50820 52946
rect 50540 52892 50820 52894
rect 50540 52162 50596 52892
rect 50764 52882 50820 52892
rect 51212 52274 51268 53004
rect 51324 52500 51380 53340
rect 51548 53172 51604 53452
rect 51660 53414 51716 53452
rect 51548 53058 51604 53116
rect 51548 53006 51550 53058
rect 51602 53006 51604 53058
rect 51548 52994 51604 53006
rect 51660 53060 51716 53070
rect 51716 53004 51828 53060
rect 51660 52994 51716 53004
rect 51324 52434 51380 52444
rect 51212 52222 51214 52274
rect 51266 52222 51268 52274
rect 50540 52110 50542 52162
rect 50594 52110 50596 52162
rect 50540 52098 50596 52110
rect 50988 52162 51044 52174
rect 50988 52110 50990 52162
rect 51042 52110 51044 52162
rect 50988 51940 51044 52110
rect 50428 51884 51044 51940
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 48860 51550 48862 51602
rect 48914 51550 48916 51602
rect 48860 51538 48916 51550
rect 48748 51438 48750 51490
rect 48802 51438 48804 51490
rect 48748 51426 48804 51438
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50876 49922 50932 49934
rect 50876 49870 50878 49922
rect 50930 49870 50932 49922
rect 50764 49812 50820 49822
rect 50764 49718 50820 49756
rect 49868 49700 49924 49710
rect 49644 49698 49924 49700
rect 49644 49646 49870 49698
rect 49922 49646 49924 49698
rect 49644 49644 49924 49646
rect 48860 49588 48916 49598
rect 48860 49138 48916 49532
rect 48860 49086 48862 49138
rect 48914 49086 48916 49138
rect 48860 49074 48916 49086
rect 49644 49026 49700 49644
rect 49644 48974 49646 49026
rect 49698 48974 49700 49026
rect 49644 48962 49700 48974
rect 49196 48356 49252 48366
rect 49196 48242 49252 48300
rect 49196 48190 49198 48242
rect 49250 48190 49252 48242
rect 48860 48132 48916 48142
rect 49196 48132 49252 48190
rect 48860 48130 49252 48132
rect 48860 48078 48862 48130
rect 48914 48078 49252 48130
rect 48860 48076 49252 48078
rect 49644 48130 49700 48142
rect 49644 48078 49646 48130
rect 49698 48078 49700 48130
rect 48860 48066 48916 48076
rect 48860 47236 48916 47246
rect 48748 46788 48804 46798
rect 48748 46694 48804 46732
rect 48748 45332 48804 45342
rect 48748 45238 48804 45276
rect 48636 41246 48638 41298
rect 48690 41246 48692 41298
rect 48636 41234 48692 41246
rect 45836 40462 45838 40514
rect 45890 40462 45892 40514
rect 45836 40450 45892 40462
rect 47964 40292 48020 40302
rect 47516 40290 48020 40292
rect 47516 40238 47966 40290
rect 48018 40238 48020 40290
rect 47516 40236 48020 40238
rect 45836 39844 45892 39854
rect 45836 39750 45892 39788
rect 45276 39678 45278 39730
rect 45330 39678 45332 39730
rect 45276 39666 45332 39678
rect 47516 39730 47572 40236
rect 47964 40226 48020 40236
rect 47516 39678 47518 39730
rect 47570 39678 47572 39730
rect 47516 39666 47572 39678
rect 48748 39844 48804 39854
rect 45388 39618 45444 39630
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 45052 39508 45108 39518
rect 45052 39414 45108 39452
rect 45388 39284 45444 39566
rect 47404 39620 47460 39630
rect 47404 39526 47460 39564
rect 45724 39508 45780 39518
rect 45724 39414 45780 39452
rect 45836 39394 45892 39406
rect 45836 39342 45838 39394
rect 45890 39342 45892 39394
rect 45836 39284 45892 39342
rect 45388 39228 45892 39284
rect 45836 38948 45892 39228
rect 48748 39284 48804 39788
rect 45836 38892 46340 38948
rect 45948 38724 46004 38734
rect 45724 38722 46004 38724
rect 45724 38670 45950 38722
rect 46002 38670 46004 38722
rect 45724 38668 46004 38670
rect 44940 38612 45108 38668
rect 43820 37490 44324 37492
rect 43820 37438 44270 37490
rect 44322 37438 44324 37490
rect 43820 37436 44324 37438
rect 43820 37266 43876 37436
rect 44268 37426 44324 37436
rect 43820 37214 43822 37266
rect 43874 37214 43876 37266
rect 43820 37202 43876 37214
rect 44044 36372 44100 36382
rect 44044 36370 44996 36372
rect 44044 36318 44046 36370
rect 44098 36318 44996 36370
rect 44044 36316 44996 36318
rect 44044 36306 44100 36316
rect 43820 36258 43876 36270
rect 43820 36206 43822 36258
rect 43874 36206 43876 36258
rect 43820 35476 43876 36206
rect 43932 36258 43988 36270
rect 43932 36206 43934 36258
rect 43986 36206 43988 36258
rect 43932 35924 43988 36206
rect 43932 35868 44884 35924
rect 44828 35810 44884 35868
rect 44828 35758 44830 35810
rect 44882 35758 44884 35810
rect 44828 35746 44884 35758
rect 43820 35420 44100 35476
rect 42700 34402 42756 34412
rect 43260 34972 43764 35028
rect 44044 35026 44100 35420
rect 44940 35138 44996 36316
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44940 35074 44996 35086
rect 44044 34974 44046 35026
rect 44098 34974 44100 35026
rect 43260 33348 43316 34972
rect 44044 34962 44100 34974
rect 45052 35028 45108 38612
rect 45724 38164 45780 38668
rect 45948 38658 46004 38668
rect 46172 38724 46228 38734
rect 46172 38630 46228 38668
rect 46284 38668 46340 38892
rect 48748 38836 48804 39228
rect 48860 39060 48916 47180
rect 48972 39620 49028 48076
rect 49644 48020 49700 48078
rect 49308 46676 49364 46686
rect 49364 46620 49588 46676
rect 49308 46582 49364 46620
rect 49308 45890 49364 45902
rect 49308 45838 49310 45890
rect 49362 45838 49364 45890
rect 49308 45780 49364 45838
rect 49084 45220 49140 45230
rect 49084 45126 49140 45164
rect 49196 41972 49252 41982
rect 49196 41878 49252 41916
rect 49084 40962 49140 40974
rect 49084 40910 49086 40962
rect 49138 40910 49140 40962
rect 49084 39844 49140 40910
rect 49084 39778 49140 39788
rect 48972 39564 49140 39620
rect 48972 39394 49028 39406
rect 48972 39342 48974 39394
rect 49026 39342 49028 39394
rect 48972 39284 49028 39342
rect 48972 39218 49028 39228
rect 48860 39004 49028 39060
rect 48860 38836 48916 38846
rect 48748 38834 48916 38836
rect 48748 38782 48862 38834
rect 48914 38782 48916 38834
rect 48748 38780 48916 38782
rect 48860 38770 48916 38780
rect 46284 38612 46564 38668
rect 46508 38610 46564 38612
rect 46508 38558 46510 38610
rect 46562 38558 46564 38610
rect 46508 38276 46564 38558
rect 46508 38220 46788 38276
rect 45388 38052 45444 38062
rect 45052 34916 45108 34972
rect 44940 34860 45108 34916
rect 45276 38050 45444 38052
rect 45276 37998 45390 38050
rect 45442 37998 45444 38050
rect 45276 37996 45444 37998
rect 45724 38052 45780 38108
rect 46396 38164 46452 38174
rect 46396 38070 46452 38108
rect 45836 38052 45892 38062
rect 45724 38050 45892 38052
rect 45724 37998 45838 38050
rect 45890 37998 45892 38050
rect 45724 37996 45892 37998
rect 45276 37826 45332 37996
rect 45388 37986 45444 37996
rect 45836 37986 45892 37996
rect 46060 38052 46116 38062
rect 46060 37938 46116 37996
rect 46060 37886 46062 37938
rect 46114 37886 46116 37938
rect 46060 37874 46116 37886
rect 46620 37940 46676 37950
rect 45276 37774 45278 37826
rect 45330 37774 45332 37826
rect 43596 34802 43652 34814
rect 43596 34750 43598 34802
rect 43650 34750 43652 34802
rect 43596 34468 43652 34750
rect 43820 34804 43876 34842
rect 44156 34804 44212 34814
rect 43820 34738 43876 34748
rect 44044 34802 44212 34804
rect 44044 34750 44158 34802
rect 44210 34750 44212 34802
rect 44044 34748 44212 34750
rect 43596 34402 43652 34412
rect 44044 34356 44100 34748
rect 44156 34738 44212 34748
rect 44268 34804 44324 34814
rect 43260 33282 43316 33292
rect 43708 34300 44100 34356
rect 44268 34354 44324 34748
rect 44940 34802 44996 34860
rect 44940 34750 44942 34802
rect 44994 34750 44996 34802
rect 44940 34738 44996 34750
rect 45052 34746 45108 34758
rect 45052 34694 45054 34746
rect 45106 34694 45108 34746
rect 44268 34302 44270 34354
rect 44322 34302 44324 34354
rect 43372 33236 43428 33246
rect 43708 33236 43764 34300
rect 44268 34290 44324 34302
rect 44492 34468 44548 34478
rect 44492 34354 44548 34412
rect 44492 34302 44494 34354
rect 44546 34302 44548 34354
rect 44492 34290 44548 34302
rect 43932 34130 43988 34142
rect 43932 34078 43934 34130
rect 43986 34078 43988 34130
rect 43932 33348 43988 34078
rect 44604 34132 44660 34142
rect 44604 34038 44660 34076
rect 45052 34132 45108 34694
rect 45052 34066 45108 34076
rect 43428 33234 43764 33236
rect 43428 33182 43710 33234
rect 43762 33182 43764 33234
rect 43428 33180 43764 33182
rect 43372 32786 43428 33180
rect 43708 33170 43764 33180
rect 43820 33346 43988 33348
rect 43820 33294 43934 33346
rect 43986 33294 43988 33346
rect 43820 33292 43988 33294
rect 43372 32734 43374 32786
rect 43426 32734 43428 32786
rect 43372 32722 43428 32734
rect 43596 32452 43652 32462
rect 43596 32358 43652 32396
rect 43260 32340 43316 32350
rect 42140 31892 42532 31948
rect 43036 32338 43316 32340
rect 43036 32286 43262 32338
rect 43314 32286 43316 32338
rect 43036 32284 43316 32286
rect 42140 31890 42196 31892
rect 42140 31838 42142 31890
rect 42194 31838 42196 31890
rect 42140 31826 42196 31838
rect 41692 31500 41972 31556
rect 41468 29316 41524 29326
rect 41468 28754 41524 29260
rect 41468 28702 41470 28754
rect 41522 28702 41524 28754
rect 41468 28690 41524 28702
rect 41692 26908 41748 31500
rect 42364 30994 42420 31892
rect 43036 31106 43092 32284
rect 43260 32274 43316 32284
rect 43708 32004 43764 32014
rect 43820 32004 43876 33292
rect 43932 33282 43988 33292
rect 43708 32002 43876 32004
rect 43708 31950 43710 32002
rect 43762 31950 43876 32002
rect 43708 31948 43876 31950
rect 43932 32562 43988 32574
rect 43932 32510 43934 32562
rect 43986 32510 43988 32562
rect 43932 32004 43988 32510
rect 44156 32562 44212 32574
rect 44156 32510 44158 32562
rect 44210 32510 44212 32562
rect 44044 32452 44100 32462
rect 44044 32358 44100 32396
rect 44044 32004 44100 32014
rect 43932 32002 44100 32004
rect 43932 31950 44046 32002
rect 44098 31950 44100 32002
rect 43932 31948 44100 31950
rect 43708 31938 43764 31948
rect 43036 31054 43038 31106
rect 43090 31054 43092 31106
rect 43036 31042 43092 31054
rect 42364 30942 42366 30994
rect 42418 30942 42420 30994
rect 42364 30212 42420 30942
rect 43932 30772 43988 31948
rect 44044 31938 44100 31948
rect 44156 31780 44212 32510
rect 44492 32564 44548 32574
rect 44940 32564 44996 32574
rect 45276 32564 45332 37774
rect 45948 37826 46004 37838
rect 45948 37774 45950 37826
rect 46002 37774 46004 37826
rect 45948 37492 46004 37774
rect 45948 37436 46564 37492
rect 46508 37378 46564 37436
rect 46620 37490 46676 37884
rect 46620 37438 46622 37490
rect 46674 37438 46676 37490
rect 46620 37426 46676 37438
rect 46732 37490 46788 38220
rect 48524 37940 48580 37950
rect 48524 37846 48580 37884
rect 46732 37438 46734 37490
rect 46786 37438 46788 37490
rect 46732 37426 46788 37438
rect 46508 37326 46510 37378
rect 46562 37326 46564 37378
rect 46508 37314 46564 37326
rect 45500 35700 45556 35710
rect 45500 35606 45556 35644
rect 45500 35028 45556 35038
rect 45500 34934 45556 34972
rect 46060 35026 46116 35038
rect 46060 34974 46062 35026
rect 46114 34974 46116 35026
rect 45724 34132 45780 34142
rect 45724 34038 45780 34076
rect 45948 34132 46004 34142
rect 46060 34132 46116 34974
rect 48860 35028 48916 35038
rect 48860 34914 48916 34972
rect 48860 34862 48862 34914
rect 48914 34862 48916 34914
rect 48188 34804 48244 34814
rect 47292 34802 48244 34804
rect 47292 34750 48190 34802
rect 48242 34750 48244 34802
rect 47292 34748 48244 34750
rect 45948 34130 46116 34132
rect 45948 34078 45950 34130
rect 46002 34078 46116 34130
rect 45948 34076 46116 34078
rect 47180 34242 47236 34254
rect 47180 34190 47182 34242
rect 47234 34190 47236 34242
rect 45948 33124 46004 34076
rect 46620 34020 46676 34030
rect 46956 34020 47012 34030
rect 46620 34018 47012 34020
rect 46620 33966 46622 34018
rect 46674 33966 46958 34018
rect 47010 33966 47012 34018
rect 46620 33964 47012 33966
rect 46620 33954 46676 33964
rect 46956 33954 47012 33964
rect 47180 33796 47236 34190
rect 47292 34018 47348 34748
rect 48188 34738 48244 34748
rect 47740 34356 47796 34366
rect 47740 34020 47796 34300
rect 47292 33966 47294 34018
rect 47346 33966 47348 34018
rect 47292 33954 47348 33966
rect 47628 34018 47796 34020
rect 47628 33966 47742 34018
rect 47794 33966 47796 34018
rect 47628 33964 47796 33966
rect 47628 33796 47684 33964
rect 47740 33954 47796 33964
rect 47180 33740 47684 33796
rect 45948 33058 46004 33068
rect 44492 32562 45332 32564
rect 44492 32510 44494 32562
rect 44546 32510 44942 32562
rect 44994 32510 45332 32562
rect 44492 32508 45332 32510
rect 46732 32564 46788 32574
rect 44268 31780 44324 31790
rect 44156 31724 44268 31780
rect 44268 31686 44324 31724
rect 41916 30156 42364 30212
rect 41916 29988 41972 30156
rect 42364 30146 42420 30156
rect 43484 30716 43988 30772
rect 41804 29204 41860 29214
rect 41804 27970 41860 29148
rect 41804 27918 41806 27970
rect 41858 27918 41860 27970
rect 41804 27906 41860 27918
rect 41916 28754 41972 29932
rect 42924 29652 42980 29662
rect 43484 29652 43540 30716
rect 42924 29650 43540 29652
rect 42924 29598 42926 29650
rect 42978 29598 43486 29650
rect 43538 29598 43540 29650
rect 42924 29596 43540 29598
rect 42924 29586 42980 29596
rect 43484 29586 43540 29596
rect 44044 29314 44100 29326
rect 44044 29262 44046 29314
rect 44098 29262 44100 29314
rect 42812 29204 42868 29214
rect 42812 29110 42868 29148
rect 43148 29204 43204 29214
rect 43148 29202 43428 29204
rect 43148 29150 43150 29202
rect 43202 29150 43428 29202
rect 43148 29148 43428 29150
rect 43148 29138 43204 29148
rect 41916 28702 41918 28754
rect 41970 28702 41972 28754
rect 41916 27860 41972 28702
rect 43372 28756 43428 29148
rect 43820 29202 43876 29214
rect 43820 29150 43822 29202
rect 43874 29150 43876 29202
rect 43484 28756 43540 28766
rect 43372 28754 43540 28756
rect 43372 28702 43486 28754
rect 43538 28702 43540 28754
rect 43372 28700 43540 28702
rect 43484 28690 43540 28700
rect 42700 28644 42756 28654
rect 42924 28644 42980 28654
rect 42700 28642 42980 28644
rect 42700 28590 42702 28642
rect 42754 28590 42926 28642
rect 42978 28590 42980 28642
rect 42700 28588 42980 28590
rect 42700 27972 42756 28588
rect 42924 28578 42980 28588
rect 43372 28420 43428 28430
rect 43372 28326 43428 28364
rect 43596 28420 43652 28430
rect 43820 28420 43876 29150
rect 44044 28420 44100 29262
rect 43596 28418 43876 28420
rect 43596 28366 43598 28418
rect 43650 28366 43876 28418
rect 43596 28364 43876 28366
rect 43932 28364 44044 28420
rect 41916 27186 41972 27804
rect 41916 27134 41918 27186
rect 41970 27134 41972 27186
rect 41916 26964 41972 27134
rect 42364 27916 42756 27972
rect 42364 26908 42420 27916
rect 43596 27524 43652 28364
rect 43932 27746 43988 28364
rect 44044 28354 44100 28364
rect 44380 28756 44436 28766
rect 44380 28082 44436 28700
rect 44380 28030 44382 28082
rect 44434 28030 44436 28082
rect 44380 28018 44436 28030
rect 43932 27694 43934 27746
rect 43986 27694 43988 27746
rect 43932 27682 43988 27694
rect 43596 27468 44100 27524
rect 41692 26852 41860 26908
rect 41916 26898 41972 26908
rect 41468 26404 41524 26414
rect 41468 26310 41524 26348
rect 41356 26066 41412 26078
rect 41356 26014 41358 26066
rect 41410 26014 41412 26066
rect 41356 25284 41412 26014
rect 41468 25396 41524 25406
rect 41468 25302 41524 25340
rect 41356 25218 41412 25228
rect 41692 25282 41748 25294
rect 41692 25230 41694 25282
rect 41746 25230 41748 25282
rect 41244 24658 41300 24668
rect 41020 24612 41076 24622
rect 40460 20178 40516 20188
rect 40572 23492 40852 23548
rect 40908 24610 41076 24612
rect 40908 24558 41022 24610
rect 41074 24558 41076 24610
rect 40908 24556 41076 24558
rect 40348 20132 40404 20142
rect 40348 20038 40404 20076
rect 40236 18900 40292 18910
rect 40236 18450 40292 18844
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 40236 18340 40292 18398
rect 40236 18274 40292 18284
rect 40572 18116 40628 23492
rect 40684 22484 40740 22494
rect 40684 22390 40740 22428
rect 40908 21812 40964 24556
rect 41020 24546 41076 24556
rect 41020 23380 41076 23390
rect 41076 23324 41300 23380
rect 41020 23286 41076 23324
rect 41244 22370 41300 23324
rect 41244 22318 41246 22370
rect 41298 22318 41300 22370
rect 41244 22306 41300 22318
rect 40908 21746 40964 21756
rect 41468 22260 41524 22270
rect 41468 21810 41524 22204
rect 41468 21758 41470 21810
rect 41522 21758 41524 21810
rect 41468 21746 41524 21758
rect 41132 21588 41188 21598
rect 40908 21586 41188 21588
rect 40908 21534 41134 21586
rect 41186 21534 41188 21586
rect 40908 21532 41188 21534
rect 40908 20018 40964 21532
rect 41132 21522 41188 21532
rect 41468 21588 41524 21598
rect 41468 21494 41524 21532
rect 41692 20804 41748 25230
rect 41804 24836 41860 26852
rect 42140 26852 42420 26908
rect 42588 26908 42644 26918
rect 43932 26852 43988 26862
rect 41916 26180 41972 26190
rect 41916 26086 41972 26124
rect 41916 25506 41972 25518
rect 41916 25454 41918 25506
rect 41970 25454 41972 25506
rect 41916 25396 41972 25454
rect 41916 25330 41972 25340
rect 42140 25172 42196 26852
rect 42588 26290 42644 26852
rect 42588 26238 42590 26290
rect 42642 26238 42644 26290
rect 42476 25284 42532 25294
rect 42588 25284 42644 26238
rect 43820 26796 43932 26852
rect 43260 26178 43316 26190
rect 43260 26126 43262 26178
rect 43314 26126 43316 26178
rect 43260 25732 43316 26126
rect 43596 25732 43652 25742
rect 43260 25730 43652 25732
rect 43260 25678 43598 25730
rect 43650 25678 43652 25730
rect 43260 25676 43652 25678
rect 43596 25666 43652 25676
rect 43708 25506 43764 25518
rect 43708 25454 43710 25506
rect 43762 25454 43764 25506
rect 42924 25284 42980 25294
rect 42588 25282 42980 25284
rect 42588 25230 42926 25282
rect 42978 25230 42980 25282
rect 42588 25228 42980 25230
rect 42476 25190 42532 25228
rect 41804 24780 41972 24836
rect 41804 24612 41860 24622
rect 41804 24518 41860 24556
rect 41916 23492 41972 24780
rect 42140 24834 42196 25116
rect 42140 24782 42142 24834
rect 42194 24782 42196 24834
rect 42140 24770 42196 24782
rect 42700 24722 42756 24734
rect 42700 24670 42702 24722
rect 42754 24670 42756 24722
rect 42700 24612 42756 24670
rect 42700 23604 42756 24556
rect 42700 23538 42756 23548
rect 41804 23380 41860 23390
rect 41916 23380 41972 23436
rect 42476 23492 42532 23502
rect 41804 23378 41972 23380
rect 41804 23326 41806 23378
rect 41858 23326 41972 23378
rect 41804 23324 41972 23326
rect 42028 23380 42084 23390
rect 42028 23378 42420 23380
rect 42028 23326 42030 23378
rect 42082 23326 42420 23378
rect 42028 23324 42420 23326
rect 41804 23314 41860 23324
rect 42028 23314 42084 23324
rect 42252 23154 42308 23166
rect 42252 23102 42254 23154
rect 42306 23102 42308 23154
rect 42140 23042 42196 23054
rect 42140 22990 42142 23042
rect 42194 22990 42196 23042
rect 42140 22484 42196 22990
rect 41804 22428 42196 22484
rect 42252 22484 42308 23102
rect 41804 21698 41860 22428
rect 42252 22418 42308 22428
rect 42028 22260 42084 22270
rect 42028 22166 42084 22204
rect 41804 21646 41806 21698
rect 41858 21646 41860 21698
rect 41804 21634 41860 21646
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40908 19796 40964 19966
rect 41132 20748 41748 20804
rect 41020 19908 41076 19918
rect 41020 19814 41076 19852
rect 40908 19730 40964 19740
rect 40572 18050 40628 18060
rect 40012 18004 40068 18014
rect 39900 17948 40012 18004
rect 40012 17938 40068 17948
rect 39788 17714 39844 17724
rect 40684 17780 40740 17790
rect 40572 17668 40628 17678
rect 39676 15876 39732 15886
rect 39228 15428 39284 15438
rect 39228 15334 39284 15372
rect 39676 15316 39732 15820
rect 39676 15222 39732 15260
rect 40236 15314 40292 15326
rect 40236 15262 40238 15314
rect 40290 15262 40292 15314
rect 39788 15202 39844 15214
rect 39788 15150 39790 15202
rect 39842 15150 39844 15202
rect 39788 14532 39844 15150
rect 39676 14530 39844 14532
rect 39676 14478 39790 14530
rect 39842 14478 39844 14530
rect 39676 14476 39844 14478
rect 39004 14254 39006 14306
rect 39058 14254 39060 14306
rect 39004 13748 39060 14254
rect 39116 14418 39172 14430
rect 39564 14420 39620 14430
rect 39116 14366 39118 14418
rect 39170 14366 39172 14418
rect 39116 13972 39172 14366
rect 39116 13906 39172 13916
rect 39340 14364 39564 14420
rect 39004 13692 39284 13748
rect 39004 13524 39060 13534
rect 38892 13522 39060 13524
rect 38892 13470 39006 13522
rect 39058 13470 39060 13522
rect 38892 13468 39060 13470
rect 38780 12964 38836 12974
rect 38780 12870 38836 12908
rect 38780 12178 38836 12190
rect 38780 12126 38782 12178
rect 38834 12126 38836 12178
rect 38780 11956 38836 12126
rect 38892 11956 38948 13468
rect 39004 13458 39060 13468
rect 39116 13524 39172 13534
rect 39116 13430 39172 13468
rect 39228 12516 39284 13692
rect 39340 13746 39396 14364
rect 39564 14326 39620 14364
rect 39340 13694 39342 13746
rect 39394 13694 39396 13746
rect 39340 13682 39396 13694
rect 39564 13748 39620 13758
rect 39676 13748 39732 14476
rect 39788 14466 39844 14476
rect 40012 14756 40068 14766
rect 39564 13746 39732 13748
rect 39564 13694 39566 13746
rect 39618 13694 39732 13746
rect 39564 13692 39732 13694
rect 40012 13970 40068 14700
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 39564 13682 39620 13692
rect 40012 13524 40068 13918
rect 40012 13458 40068 13468
rect 39676 12964 39732 12974
rect 39676 12870 39732 12908
rect 39228 12460 39844 12516
rect 39004 12404 39060 12414
rect 39004 12402 39620 12404
rect 39004 12350 39006 12402
rect 39058 12350 39620 12402
rect 39004 12348 39620 12350
rect 39004 12338 39060 12348
rect 39116 12180 39172 12190
rect 39116 12086 39172 12124
rect 39228 12178 39284 12190
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 11956 39284 12126
rect 39564 12178 39620 12348
rect 39564 12126 39566 12178
rect 39618 12126 39620 12178
rect 39564 12114 39620 12126
rect 39788 12180 39844 12460
rect 39900 12404 39956 12414
rect 40236 12404 40292 15262
rect 39900 12402 40180 12404
rect 39900 12350 39902 12402
rect 39954 12350 40180 12402
rect 39900 12348 40180 12350
rect 39900 12338 39956 12348
rect 39900 12180 39956 12190
rect 39788 12178 39956 12180
rect 39788 12126 39902 12178
rect 39954 12126 39956 12178
rect 39788 12124 39956 12126
rect 39900 12114 39956 12124
rect 38892 11900 39284 11956
rect 38780 11890 38836 11900
rect 38668 11620 38724 11630
rect 38556 11564 38668 11620
rect 37884 11506 37940 11564
rect 37884 11454 37886 11506
rect 37938 11454 37940 11506
rect 37884 11442 37940 11454
rect 38332 11508 38388 11518
rect 38332 11414 38388 11452
rect 38668 11394 38724 11564
rect 38668 11342 38670 11394
rect 38722 11342 38724 11394
rect 38668 11330 38724 11342
rect 39452 11508 39508 11518
rect 40124 11508 40180 12348
rect 40236 12338 40292 12348
rect 40236 12178 40292 12190
rect 40236 12126 40238 12178
rect 40290 12126 40292 12178
rect 40236 12068 40292 12126
rect 40236 12002 40292 12012
rect 40236 11508 40292 11518
rect 40124 11506 40292 11508
rect 40124 11454 40238 11506
rect 40290 11454 40292 11506
rect 40124 11452 40292 11454
rect 39452 11394 39508 11452
rect 40236 11442 40292 11452
rect 39452 11342 39454 11394
rect 39506 11342 39508 11394
rect 39004 11170 39060 11182
rect 39004 11118 39006 11170
rect 39058 11118 39060 11170
rect 39004 10836 39060 11118
rect 39004 10770 39060 10780
rect 37772 9662 37774 9714
rect 37826 9662 37828 9714
rect 37772 9650 37828 9662
rect 37324 9492 37380 9502
rect 37100 9154 37268 9156
rect 37100 9102 37102 9154
rect 37154 9102 37268 9154
rect 37100 9100 37268 9102
rect 37100 9090 37156 9100
rect 35868 8978 35924 8988
rect 35420 8930 35476 8942
rect 35420 8878 35422 8930
rect 35474 8878 35476 8930
rect 35420 8820 35476 8878
rect 35420 8764 35588 8820
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35308 8484 35364 8494
rect 35532 8484 35588 8764
rect 35308 8482 35924 8484
rect 35308 8430 35310 8482
rect 35362 8430 35924 8482
rect 35308 8428 35924 8430
rect 35308 8418 35364 8428
rect 35532 8258 35588 8270
rect 35532 8206 35534 8258
rect 35586 8206 35588 8258
rect 35532 8036 35588 8206
rect 35868 8258 35924 8428
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 8194 35924 8206
rect 36316 8260 36372 8270
rect 36316 8146 36372 8204
rect 36316 8094 36318 8146
rect 36370 8094 36372 8146
rect 35532 7970 35588 7980
rect 35980 8034 36036 8046
rect 35980 7982 35982 8034
rect 36034 7982 36036 8034
rect 35644 7588 35700 7598
rect 35644 7494 35700 7532
rect 35084 7422 35086 7474
rect 35138 7422 35140 7474
rect 34636 5170 34692 5180
rect 32060 5058 32116 5068
rect 32284 5122 33236 5124
rect 32284 5070 32734 5122
rect 32786 5070 33236 5122
rect 32284 5068 33236 5070
rect 31500 4398 31502 4450
rect 31554 4398 31556 4450
rect 31500 4386 31556 4398
rect 32284 4338 32340 5068
rect 32732 5058 32788 5068
rect 33180 4562 33236 5068
rect 33180 4510 33182 4562
rect 33234 4510 33236 4562
rect 33180 4498 33236 4510
rect 32284 4286 32286 4338
rect 32338 4286 32340 4338
rect 32284 4274 32340 4286
rect 29372 4174 29374 4226
rect 29426 4174 29428 4226
rect 29372 4162 29428 4174
rect 34300 4228 34356 4238
rect 35084 4228 35140 7422
rect 35308 7474 35364 7486
rect 35308 7422 35310 7474
rect 35362 7422 35364 7474
rect 35308 7252 35364 7422
rect 35420 7476 35476 7486
rect 35980 7476 36036 7982
rect 36092 8036 36148 8046
rect 36092 7700 36148 7980
rect 36316 7924 36372 8094
rect 36316 7858 36372 7868
rect 36092 7644 36372 7700
rect 36092 7476 36148 7486
rect 35980 7474 36148 7476
rect 35980 7422 36094 7474
rect 36146 7422 36148 7474
rect 35980 7420 36148 7422
rect 35420 7382 35476 7420
rect 36092 7410 36148 7420
rect 35980 7252 36036 7262
rect 35308 7196 35588 7252
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35420 6020 35476 6030
rect 35532 6020 35588 7196
rect 35980 7158 36036 7196
rect 36204 7252 36260 7262
rect 36204 6802 36260 7196
rect 36316 7140 36372 7644
rect 36428 7588 36484 7598
rect 36428 7494 36484 7532
rect 36764 7474 36820 7486
rect 36764 7422 36766 7474
rect 36818 7422 36820 7474
rect 36764 7252 36820 7422
rect 36764 7186 36820 7196
rect 36428 7140 36484 7150
rect 36316 7084 36428 7140
rect 36428 7074 36484 7084
rect 37212 6916 37268 9100
rect 37324 9154 37380 9436
rect 39228 9268 39284 9278
rect 39228 9174 39284 9212
rect 37324 9102 37326 9154
rect 37378 9102 37380 9154
rect 37324 9090 37380 9102
rect 37660 9156 37716 9166
rect 37660 9062 37716 9100
rect 37548 8930 37604 8942
rect 37548 8878 37550 8930
rect 37602 8878 37604 8930
rect 37548 7476 37604 8878
rect 39452 8428 39508 11342
rect 40236 10836 40292 10846
rect 39564 9714 39620 9726
rect 39564 9662 39566 9714
rect 39618 9662 39620 9714
rect 39564 9380 39620 9662
rect 39564 9324 40068 9380
rect 39564 9154 39620 9324
rect 39564 9102 39566 9154
rect 39618 9102 39620 9154
rect 39564 9090 39620 9102
rect 39788 9156 39844 9166
rect 39452 8372 39620 8428
rect 39004 8148 39060 8158
rect 39004 8054 39060 8092
rect 39340 8034 39396 8046
rect 39340 7982 39342 8034
rect 39394 7982 39396 8034
rect 38892 7924 38948 7934
rect 38444 7700 38500 7710
rect 37884 7698 38500 7700
rect 37884 7646 38446 7698
rect 38498 7646 38500 7698
rect 37884 7644 38500 7646
rect 37884 7476 37940 7644
rect 38444 7634 38500 7644
rect 38892 7698 38948 7868
rect 38892 7646 38894 7698
rect 38946 7646 38948 7698
rect 38892 7634 38948 7646
rect 37548 7474 37940 7476
rect 37548 7422 37886 7474
rect 37938 7422 37940 7474
rect 37548 7420 37940 7422
rect 37884 7410 37940 7420
rect 38108 7476 38164 7486
rect 38108 7382 38164 7420
rect 38668 7476 38724 7486
rect 38668 7382 38724 7420
rect 38220 7364 38276 7374
rect 37548 7250 37604 7262
rect 37548 7198 37550 7250
rect 37602 7198 37604 7250
rect 37548 7140 37604 7198
rect 37548 7074 37604 7084
rect 36204 6750 36206 6802
rect 36258 6750 36260 6802
rect 36204 6738 36260 6750
rect 36988 6860 37940 6916
rect 35420 6018 35588 6020
rect 35420 5966 35422 6018
rect 35474 5966 35588 6018
rect 35420 5964 35588 5966
rect 35420 5954 35476 5964
rect 35532 5684 35588 5694
rect 35532 5682 36484 5684
rect 35532 5630 35534 5682
rect 35586 5630 36484 5682
rect 35532 5628 36484 5630
rect 35532 5618 35588 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 5236 35700 5246
rect 35644 5142 35700 5180
rect 36428 4450 36484 5628
rect 36988 5234 37044 6860
rect 37884 6690 37940 6860
rect 37884 6638 37886 6690
rect 37938 6638 37940 6690
rect 37884 6626 37940 6638
rect 38220 6690 38276 7308
rect 38556 7362 38612 7374
rect 38556 7310 38558 7362
rect 38610 7310 38612 7362
rect 38556 7252 38612 7310
rect 39340 7364 39396 7982
rect 38556 7196 38948 7252
rect 38780 7028 38836 7038
rect 38780 6914 38836 6972
rect 38780 6862 38782 6914
rect 38834 6862 38836 6914
rect 38780 6850 38836 6862
rect 38892 6914 38948 7196
rect 38892 6862 38894 6914
rect 38946 6862 38948 6914
rect 38892 6850 38948 6862
rect 38220 6638 38222 6690
rect 38274 6638 38276 6690
rect 38220 6626 38276 6638
rect 38556 6692 38612 6702
rect 38556 6578 38612 6636
rect 38556 6526 38558 6578
rect 38610 6526 38612 6578
rect 38556 6514 38612 6526
rect 39340 6580 39396 7308
rect 39340 6514 39396 6524
rect 38108 6466 38164 6478
rect 38108 6414 38110 6466
rect 38162 6414 38164 6466
rect 36988 5182 36990 5234
rect 37042 5182 37044 5234
rect 36988 5170 37044 5182
rect 37660 5348 37716 5358
rect 37660 4564 37716 5292
rect 36428 4398 36430 4450
rect 36482 4398 36484 4450
rect 36428 4386 36484 4398
rect 37212 4562 37716 4564
rect 37212 4510 37662 4562
rect 37714 4510 37716 4562
rect 37212 4508 37716 4510
rect 37212 4338 37268 4508
rect 37660 4498 37716 4508
rect 38108 4450 38164 6414
rect 39564 5348 39620 8372
rect 39676 8148 39732 8158
rect 39676 8054 39732 8092
rect 39788 7586 39844 9100
rect 39900 9154 39956 9166
rect 39900 9102 39902 9154
rect 39954 9102 39956 9154
rect 39900 7924 39956 9102
rect 40012 8148 40068 9324
rect 40236 9266 40292 10780
rect 40460 10388 40516 10398
rect 40348 9716 40404 9726
rect 40348 9622 40404 9660
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 40236 9202 40292 9214
rect 40460 8260 40516 10332
rect 40572 9268 40628 17612
rect 40684 15316 40740 17724
rect 41132 16996 41188 20748
rect 41580 20578 41636 20590
rect 41580 20526 41582 20578
rect 41634 20526 41636 20578
rect 41580 20468 41636 20526
rect 41580 20412 41860 20468
rect 41244 20132 41300 20142
rect 41244 20038 41300 20076
rect 41468 20020 41524 20030
rect 41468 19926 41524 19964
rect 41804 20018 41860 20412
rect 41804 19966 41806 20018
rect 41858 19966 41860 20018
rect 41804 19236 41860 19966
rect 42140 20020 42196 20030
rect 41692 19180 41860 19236
rect 41916 19796 41972 19806
rect 41244 18788 41300 18798
rect 41244 18674 41300 18732
rect 41244 18622 41246 18674
rect 41298 18622 41300 18674
rect 41244 18610 41300 18622
rect 41356 18452 41412 18462
rect 41356 18358 41412 18396
rect 41468 18450 41524 18462
rect 41468 18398 41470 18450
rect 41522 18398 41524 18450
rect 41468 17892 41524 18398
rect 41468 17826 41524 17836
rect 40908 16940 41188 16996
rect 41468 17668 41524 17678
rect 41692 17668 41748 19180
rect 41804 19010 41860 19022
rect 41804 18958 41806 19010
rect 41858 18958 41860 19010
rect 41804 18450 41860 18958
rect 41916 18788 41972 19740
rect 42140 19346 42196 19964
rect 42140 19294 42142 19346
rect 42194 19294 42196 19346
rect 42140 19282 42196 19294
rect 42364 19460 42420 23324
rect 42476 23378 42532 23436
rect 42476 23326 42478 23378
rect 42530 23326 42532 23378
rect 42476 23314 42532 23326
rect 42924 23380 42980 25228
rect 43260 25284 43316 25294
rect 42924 23314 42980 23324
rect 43036 24722 43092 24734
rect 43036 24670 43038 24722
rect 43090 24670 43092 24722
rect 43036 24500 43092 24670
rect 43036 22484 43092 24444
rect 42924 22428 43092 22484
rect 43148 24612 43204 24622
rect 42588 19908 42644 19918
rect 42588 19814 42644 19852
rect 42252 19236 42308 19246
rect 42364 19236 42420 19404
rect 42252 19234 42420 19236
rect 42252 19182 42254 19234
rect 42306 19182 42420 19234
rect 42252 19180 42420 19182
rect 42252 19170 42308 19180
rect 42028 19012 42084 19022
rect 42028 18918 42084 18956
rect 41916 18732 42084 18788
rect 41804 18398 41806 18450
rect 41858 18398 41860 18450
rect 41804 18340 41860 18398
rect 42028 18450 42084 18732
rect 42028 18398 42030 18450
rect 42082 18398 42084 18450
rect 42028 18386 42084 18398
rect 42364 18676 42420 18686
rect 42364 18450 42420 18620
rect 42364 18398 42366 18450
rect 42418 18398 42420 18450
rect 42364 18386 42420 18398
rect 42588 18452 42644 18462
rect 42588 18358 42644 18396
rect 41804 18274 41860 18284
rect 42252 18338 42308 18350
rect 42252 18286 42254 18338
rect 42306 18286 42308 18338
rect 42140 17780 42196 17790
rect 42252 17780 42308 18286
rect 42140 17778 42308 17780
rect 42140 17726 42142 17778
rect 42194 17726 42308 17778
rect 42140 17724 42308 17726
rect 42364 18228 42420 18238
rect 42140 17714 42196 17724
rect 41468 17666 41692 17668
rect 41468 17614 41470 17666
rect 41522 17614 41692 17666
rect 41468 17612 41692 17614
rect 40908 15764 40964 16940
rect 40908 15698 40964 15708
rect 41020 16772 41076 16782
rect 41468 16772 41524 17612
rect 41692 17574 41748 17612
rect 41020 16770 41524 16772
rect 41020 16718 41022 16770
rect 41074 16718 41470 16770
rect 41522 16718 41524 16770
rect 41020 16716 41524 16718
rect 41020 16324 41076 16716
rect 40908 15316 40964 15326
rect 40684 15314 40964 15316
rect 40684 15262 40910 15314
rect 40962 15262 40964 15314
rect 40684 15260 40964 15262
rect 40908 15250 40964 15260
rect 41020 15316 41076 16268
rect 41468 16210 41524 16716
rect 41468 16158 41470 16210
rect 41522 16158 41524 16210
rect 41468 16146 41524 16158
rect 40908 14420 40964 14430
rect 40908 12290 40964 14364
rect 40908 12238 40910 12290
rect 40962 12238 40964 12290
rect 40908 12226 40964 12238
rect 41020 13074 41076 15260
rect 41132 15876 41188 15886
rect 41132 15314 41188 15820
rect 41132 15262 41134 15314
rect 41186 15262 41188 15314
rect 41132 15250 41188 15262
rect 41916 15316 41972 15326
rect 41916 15222 41972 15260
rect 41468 15090 41524 15102
rect 41468 15038 41470 15090
rect 41522 15038 41524 15090
rect 41468 14644 41524 15038
rect 41468 14550 41524 14588
rect 41692 15092 41748 15102
rect 41692 14530 41748 15036
rect 41692 14478 41694 14530
rect 41746 14478 41748 14530
rect 41692 14466 41748 14478
rect 41916 14532 41972 14542
rect 41916 14438 41972 14476
rect 41020 13022 41022 13074
rect 41074 13022 41076 13074
rect 41020 11508 41076 13022
rect 41132 14308 41188 14318
rect 41132 12852 41188 14252
rect 41468 14308 41524 14318
rect 41468 13858 41524 14252
rect 41468 13806 41470 13858
rect 41522 13806 41524 13858
rect 41468 13794 41524 13806
rect 41916 13972 41972 13982
rect 42364 13972 42420 18172
rect 42588 15202 42644 15214
rect 42588 15150 42590 15202
rect 42642 15150 42644 15202
rect 42588 15148 42644 15150
rect 41692 13748 41748 13758
rect 41580 13746 41748 13748
rect 41580 13694 41694 13746
rect 41746 13694 41748 13746
rect 41580 13692 41748 13694
rect 41580 12852 41636 13692
rect 41692 13682 41748 13692
rect 41916 13746 41972 13916
rect 41916 13694 41918 13746
rect 41970 13694 41972 13746
rect 41916 13682 41972 13694
rect 42252 13916 42420 13972
rect 42476 15092 42644 15148
rect 42812 15092 42868 15102
rect 42476 13970 42532 15092
rect 42588 14644 42644 14654
rect 42588 14530 42644 14588
rect 42588 14478 42590 14530
rect 42642 14478 42644 14530
rect 42588 14466 42644 14478
rect 42812 14530 42868 15036
rect 42812 14478 42814 14530
rect 42866 14478 42868 14530
rect 42700 14308 42756 14318
rect 42700 14214 42756 14252
rect 42476 13918 42478 13970
rect 42530 13918 42532 13970
rect 42140 13636 42196 13646
rect 41132 12402 41188 12796
rect 41132 12350 41134 12402
rect 41186 12350 41188 12402
rect 41132 12338 41188 12350
rect 41244 12796 41636 12852
rect 42028 12852 42084 12862
rect 41244 12066 41300 12796
rect 42028 12758 42084 12796
rect 42140 12292 42196 13580
rect 42252 12516 42308 13916
rect 42476 13906 42532 13918
rect 42812 13858 42868 14478
rect 42812 13806 42814 13858
rect 42866 13806 42868 13858
rect 42812 13794 42868 13806
rect 42364 13748 42420 13758
rect 42700 13748 42756 13758
rect 42364 13746 42756 13748
rect 42364 13694 42366 13746
rect 42418 13694 42702 13746
rect 42754 13694 42756 13746
rect 42364 13692 42756 13694
rect 42364 13682 42420 13692
rect 42700 13682 42756 13692
rect 42812 13076 42868 13086
rect 42924 13076 42980 22428
rect 43148 22372 43204 24556
rect 43036 22316 43204 22372
rect 43036 14756 43092 22316
rect 43148 18676 43204 18686
rect 43148 18450 43204 18620
rect 43148 18398 43150 18450
rect 43202 18398 43204 18450
rect 43148 18386 43204 18398
rect 43036 14690 43092 14700
rect 43036 14532 43092 14542
rect 43036 14418 43092 14476
rect 43036 14366 43038 14418
rect 43090 14366 43092 14418
rect 43036 14354 43092 14366
rect 43260 13972 43316 25228
rect 43708 25284 43764 25454
rect 43708 25218 43764 25228
rect 43484 24612 43540 24622
rect 43484 24518 43540 24556
rect 43596 23604 43652 23614
rect 43372 23492 43428 23502
rect 43372 23378 43428 23436
rect 43372 23326 43374 23378
rect 43426 23326 43428 23378
rect 43372 22596 43428 23326
rect 43372 22530 43428 22540
rect 43596 22260 43652 23548
rect 43260 13878 43316 13916
rect 43484 22204 43652 22260
rect 43708 23042 43764 23054
rect 43708 22990 43710 23042
rect 43762 22990 43764 23042
rect 43708 22260 43764 22990
rect 43372 13076 43428 13086
rect 43484 13076 43540 22204
rect 43708 22194 43764 22204
rect 43596 18338 43652 18350
rect 43596 18286 43598 18338
rect 43650 18286 43652 18338
rect 43596 18228 43652 18286
rect 43596 18162 43652 18172
rect 43820 15148 43876 26796
rect 43932 26758 43988 26796
rect 44044 26852 44100 27468
rect 44268 26964 44324 27002
rect 44268 26898 44324 26908
rect 44156 26852 44212 26862
rect 44044 26850 44212 26852
rect 44044 26798 44158 26850
rect 44210 26798 44212 26850
rect 44044 26796 44212 26798
rect 43932 26068 43988 26078
rect 43932 25730 43988 26012
rect 43932 25678 43934 25730
rect 43986 25678 43988 25730
rect 43932 25666 43988 25678
rect 44044 25730 44100 26796
rect 44156 26786 44212 26796
rect 44044 25678 44046 25730
rect 44098 25678 44100 25730
rect 44044 25666 44100 25678
rect 44380 25844 44436 25854
rect 44380 25284 44436 25788
rect 44380 24946 44436 25228
rect 44380 24894 44382 24946
rect 44434 24894 44436 24946
rect 44380 24882 44436 24894
rect 44156 23492 44212 23502
rect 44156 23378 44212 23436
rect 44156 23326 44158 23378
rect 44210 23326 44212 23378
rect 44156 23314 44212 23326
rect 44156 22484 44212 22494
rect 43932 18450 43988 18462
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43932 18228 43988 18398
rect 43932 18162 43988 18172
rect 44156 16772 44212 22428
rect 44380 19908 44436 19918
rect 44380 19348 44436 19852
rect 44268 17892 44324 17902
rect 44268 17778 44324 17836
rect 44268 17726 44270 17778
rect 44322 17726 44324 17778
rect 44268 17714 44324 17726
rect 44156 16706 44212 16716
rect 44380 15148 44436 19292
rect 44492 18452 44548 32508
rect 44940 32498 44996 32508
rect 46732 32470 46788 32508
rect 47404 32564 47460 32574
rect 47404 32470 47460 32508
rect 46508 32450 46564 32462
rect 46508 32398 46510 32450
rect 46562 32398 46564 32450
rect 45388 31892 45444 31902
rect 45388 31798 45444 31836
rect 45164 31780 45220 31790
rect 45164 30882 45220 31724
rect 45164 30830 45166 30882
rect 45218 30830 45220 30882
rect 45164 30818 45220 30830
rect 45612 30882 45668 30894
rect 45612 30830 45614 30882
rect 45666 30830 45668 30882
rect 45276 30212 45332 30222
rect 45276 28756 45332 30156
rect 45612 30212 45668 30830
rect 46508 30434 46564 32398
rect 47516 31668 47572 31678
rect 47516 31574 47572 31612
rect 46508 30382 46510 30434
rect 46562 30382 46564 30434
rect 46508 30370 46564 30382
rect 46956 30324 47012 30334
rect 45612 30146 45668 30156
rect 46620 30268 46956 30324
rect 46620 30210 46676 30268
rect 46956 30230 47012 30268
rect 46620 30158 46622 30210
rect 46674 30158 46676 30210
rect 46620 30146 46676 30158
rect 46508 29986 46564 29998
rect 46508 29934 46510 29986
rect 46562 29934 46564 29986
rect 46508 29316 46564 29934
rect 46508 29250 46564 29260
rect 45332 28700 45668 28756
rect 45276 28662 45332 28700
rect 45612 28642 45668 28700
rect 45612 28590 45614 28642
rect 45666 28590 45668 28642
rect 45612 28578 45668 28590
rect 46396 28530 46452 28542
rect 46396 28478 46398 28530
rect 46450 28478 46452 28530
rect 44828 26962 44884 26974
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44828 26852 44884 26910
rect 45052 26964 45108 26974
rect 44828 26786 44884 26796
rect 44940 26850 44996 26862
rect 44940 26798 44942 26850
rect 44994 26798 44996 26850
rect 44940 26068 44996 26798
rect 44940 26002 44996 26012
rect 45052 25618 45108 26908
rect 45052 25566 45054 25618
rect 45106 25566 45108 25618
rect 45052 25554 45108 25566
rect 45164 26962 45220 26974
rect 45164 26910 45166 26962
rect 45218 26910 45220 26962
rect 45164 25508 45220 26910
rect 45388 26962 45444 26974
rect 45388 26910 45390 26962
rect 45442 26910 45444 26962
rect 45388 26180 45444 26910
rect 46396 26404 46452 28478
rect 46396 26338 46452 26348
rect 44828 25396 44884 25406
rect 44828 25302 44884 25340
rect 45052 25396 45108 25406
rect 45164 25396 45220 25452
rect 45052 25394 45220 25396
rect 45052 25342 45054 25394
rect 45106 25342 45220 25394
rect 45052 25340 45220 25342
rect 45276 26178 45444 26180
rect 45276 26126 45390 26178
rect 45442 26126 45444 26178
rect 45276 26124 45444 26126
rect 45276 25394 45332 26124
rect 45388 26114 45444 26124
rect 45836 26292 45892 26302
rect 45276 25342 45278 25394
rect 45330 25342 45332 25394
rect 45052 25330 45108 25340
rect 45276 25330 45332 25342
rect 45724 25506 45780 25518
rect 45724 25454 45726 25506
rect 45778 25454 45780 25506
rect 45164 24724 45220 24734
rect 44828 24610 44884 24622
rect 44828 24558 44830 24610
rect 44882 24558 44884 24610
rect 44828 24500 44884 24558
rect 44828 24434 44884 24444
rect 44604 24052 44660 24062
rect 44604 23378 44660 23996
rect 45164 24050 45220 24668
rect 45276 24612 45332 24622
rect 45276 24518 45332 24556
rect 45724 24612 45780 25454
rect 45836 25396 45892 26236
rect 47628 26292 47684 33740
rect 48860 33684 48916 34862
rect 48524 33628 48916 33684
rect 48972 33684 49028 39004
rect 48300 33348 48356 33358
rect 48524 33348 48580 33628
rect 48972 33618 49028 33628
rect 49084 33572 49140 39564
rect 49308 39506 49364 45724
rect 49532 45892 49588 46620
rect 49532 45778 49588 45836
rect 49532 45726 49534 45778
rect 49586 45726 49588 45778
rect 49532 45714 49588 45726
rect 49644 42530 49700 47964
rect 49868 47460 49924 49644
rect 50428 49698 50484 49710
rect 50428 49646 50430 49698
rect 50482 49646 50484 49698
rect 50428 49588 50484 49646
rect 50876 49588 50932 49870
rect 50428 49532 50932 49588
rect 50428 48916 50484 49532
rect 50204 48860 50484 48916
rect 50876 49028 50932 49038
rect 50092 48244 50148 48254
rect 50204 48244 50260 48860
rect 50876 48804 50932 48972
rect 49756 47236 49812 47246
rect 49756 47142 49812 47180
rect 49756 46676 49812 46686
rect 49756 46582 49812 46620
rect 49868 45108 49924 47404
rect 49980 48242 50260 48244
rect 49980 48190 50094 48242
rect 50146 48190 50260 48242
rect 49980 48188 50260 48190
rect 50316 48748 50932 48804
rect 50988 48802 51044 51884
rect 51100 51156 51156 51166
rect 51100 50034 51156 51100
rect 51212 50708 51268 52222
rect 51772 52274 51828 53004
rect 51772 52222 51774 52274
rect 51826 52222 51828 52274
rect 51772 52210 51828 52222
rect 51884 51602 51940 53676
rect 52780 53508 52836 53518
rect 52780 53414 52836 53452
rect 51884 51550 51886 51602
rect 51938 51550 51940 51602
rect 51884 51538 51940 51550
rect 52780 51604 52836 51614
rect 52892 51604 52948 53788
rect 53004 53750 53060 53788
rect 53676 53508 53732 53518
rect 53676 52834 53732 53452
rect 53788 52948 53844 55020
rect 53900 55524 53956 56252
rect 54236 56242 54292 56252
rect 55244 56978 55412 56980
rect 55244 56926 55358 56978
rect 55410 56926 55412 56978
rect 55244 56924 55412 56926
rect 54908 56084 54964 56094
rect 53900 53842 53956 55468
rect 54796 56082 54964 56084
rect 54796 56030 54910 56082
rect 54962 56030 54964 56082
rect 54796 56028 54964 56030
rect 54572 54292 54628 54302
rect 53900 53790 53902 53842
rect 53954 53790 53956 53842
rect 53900 53778 53956 53790
rect 54460 54290 54628 54292
rect 54460 54238 54574 54290
rect 54626 54238 54628 54290
rect 54460 54236 54628 54238
rect 54236 53618 54292 53630
rect 54236 53566 54238 53618
rect 54290 53566 54292 53618
rect 54124 52948 54180 52958
rect 53788 52946 54180 52948
rect 53788 52894 54126 52946
rect 54178 52894 54180 52946
rect 53788 52892 54180 52894
rect 54124 52882 54180 52892
rect 53676 52782 53678 52834
rect 53730 52782 53732 52834
rect 53340 52276 53396 52286
rect 52780 51602 52948 51604
rect 52780 51550 52782 51602
rect 52834 51550 52948 51602
rect 52780 51548 52948 51550
rect 53228 52164 53284 52174
rect 52780 51538 52836 51548
rect 53228 51490 53284 52108
rect 53228 51438 53230 51490
rect 53282 51438 53284 51490
rect 53228 51426 53284 51438
rect 52108 51380 52164 51390
rect 52444 51380 52500 51390
rect 52108 51378 52276 51380
rect 52108 51326 52110 51378
rect 52162 51326 52276 51378
rect 52108 51324 52276 51326
rect 52108 51314 52164 51324
rect 51772 51156 51828 51166
rect 51772 51062 51828 51100
rect 52220 51156 52276 51324
rect 52444 51286 52500 51324
rect 53116 51156 53172 51166
rect 52220 51154 53172 51156
rect 52220 51102 53118 51154
rect 53170 51102 53172 51154
rect 52220 51100 53172 51102
rect 51212 50642 51268 50652
rect 51100 49982 51102 50034
rect 51154 49982 51156 50034
rect 51100 49970 51156 49982
rect 51212 49924 51268 49934
rect 51100 49812 51156 49822
rect 51100 49026 51156 49756
rect 51100 48974 51102 49026
rect 51154 48974 51156 49026
rect 51100 48962 51156 48974
rect 50988 48750 50990 48802
rect 51042 48750 51044 48802
rect 49980 47236 50036 48188
rect 50092 48178 50148 48188
rect 50204 48020 50260 48030
rect 50316 48020 50372 48748
rect 50988 48738 51044 48750
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 51212 48580 51268 49868
rect 51660 49924 51716 49934
rect 51996 49924 52052 49934
rect 51716 49922 52052 49924
rect 51716 49870 51998 49922
rect 52050 49870 52052 49922
rect 51716 49868 52052 49870
rect 51660 49830 51716 49868
rect 51996 49858 52052 49868
rect 52220 49922 52276 51100
rect 53116 51090 53172 51100
rect 52220 49870 52222 49922
rect 52274 49870 52276 49922
rect 52220 49858 52276 49870
rect 53228 50820 53284 50830
rect 52668 49812 52724 49822
rect 52668 49718 52724 49756
rect 52444 49698 52500 49710
rect 52444 49646 52446 49698
rect 52498 49646 52500 49698
rect 52444 49364 52500 49646
rect 52444 49308 53060 49364
rect 53004 49250 53060 49308
rect 53004 49198 53006 49250
rect 53058 49198 53060 49250
rect 53004 49186 53060 49198
rect 51548 49028 51604 49038
rect 51548 48934 51604 48972
rect 52780 49026 52836 49038
rect 52780 48974 52782 49026
rect 52834 48974 52836 49026
rect 50556 48570 50820 48580
rect 50876 48524 51268 48580
rect 52108 48804 52164 48814
rect 52780 48804 52836 48974
rect 53228 49026 53284 50764
rect 53228 48974 53230 49026
rect 53282 48974 53284 49026
rect 53228 48962 53284 48974
rect 53116 48804 53172 48814
rect 52108 48802 52836 48804
rect 52108 48750 52110 48802
rect 52162 48750 52836 48802
rect 52108 48748 52836 48750
rect 53004 48802 53172 48804
rect 53004 48750 53118 48802
rect 53170 48750 53172 48802
rect 53004 48748 53172 48750
rect 50876 48130 50932 48524
rect 50876 48078 50878 48130
rect 50930 48078 50932 48130
rect 50876 48066 50932 48078
rect 49980 47170 50036 47180
rect 50092 48018 50372 48020
rect 50092 47966 50206 48018
rect 50258 47966 50372 48018
rect 50092 47964 50372 47966
rect 49980 45780 50036 45790
rect 50092 45780 50148 47964
rect 50204 47954 50260 47964
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50540 46676 50596 46686
rect 50540 46582 50596 46620
rect 50204 46564 50260 46574
rect 50316 46564 50372 46574
rect 50204 46562 50316 46564
rect 50204 46510 50206 46562
rect 50258 46510 50316 46562
rect 50204 46508 50316 46510
rect 50204 46498 50260 46508
rect 50036 45724 50148 45780
rect 49980 45686 50036 45724
rect 49980 45108 50036 45118
rect 49868 45052 49980 45108
rect 49980 45014 50036 45052
rect 50316 43092 50372 46508
rect 51100 46562 51156 46574
rect 51100 46510 51102 46562
rect 51154 46510 51156 46562
rect 50876 46002 50932 46014
rect 50876 45950 50878 46002
rect 50930 45950 50932 46002
rect 50652 45668 50708 45678
rect 50428 45666 50708 45668
rect 50428 45614 50654 45666
rect 50706 45614 50708 45666
rect 50428 45612 50708 45614
rect 50428 45220 50484 45612
rect 50652 45602 50708 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50428 45154 50484 45164
rect 50764 45220 50820 45230
rect 50876 45220 50932 45950
rect 50764 45218 50932 45220
rect 50764 45166 50766 45218
rect 50818 45166 50932 45218
rect 50764 45164 50932 45166
rect 50988 45666 51044 45678
rect 50988 45614 50990 45666
rect 51042 45614 51044 45666
rect 50988 45220 51044 45614
rect 50764 45154 50820 45164
rect 50988 45108 51044 45164
rect 50876 45052 51044 45108
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50316 43036 50484 43092
rect 50092 42980 50148 42990
rect 50092 42978 50372 42980
rect 50092 42926 50094 42978
rect 50146 42926 50372 42978
rect 50092 42924 50372 42926
rect 50092 42914 50148 42924
rect 50204 42644 50260 42654
rect 50204 42550 50260 42588
rect 49644 42478 49646 42530
rect 49698 42478 49700 42530
rect 49644 42420 49700 42478
rect 50092 42530 50148 42542
rect 50092 42478 50094 42530
rect 50146 42478 50148 42530
rect 50092 42420 50148 42478
rect 49644 42364 50148 42420
rect 49644 40964 49700 42364
rect 50204 41972 50260 41982
rect 49868 41858 49924 41870
rect 49868 41806 49870 41858
rect 49922 41806 49924 41858
rect 49868 41412 49924 41806
rect 49868 41346 49924 41356
rect 49644 40898 49700 40908
rect 49308 39454 49310 39506
rect 49362 39454 49364 39506
rect 49308 39396 49364 39454
rect 49756 39396 49812 39406
rect 49308 39394 49812 39396
rect 49308 39342 49758 39394
rect 49810 39342 49812 39394
rect 49308 39340 49812 39342
rect 49420 38724 49476 38734
rect 49644 38668 49700 39340
rect 49756 39330 49812 39340
rect 50204 38834 50260 41916
rect 50316 41410 50372 42924
rect 50316 41358 50318 41410
rect 50370 41358 50372 41410
rect 50316 41346 50372 41358
rect 50428 41188 50484 43036
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50540 41300 50596 41310
rect 50540 41206 50596 41244
rect 50204 38782 50206 38834
rect 50258 38782 50260 38834
rect 50204 38724 50260 38782
rect 49420 38630 49476 38668
rect 49532 38612 49700 38668
rect 49756 38668 50260 38724
rect 50316 41132 50484 41188
rect 50652 41188 50708 41198
rect 49532 38276 49588 38612
rect 49084 33506 49140 33516
rect 49196 38220 49588 38276
rect 48300 33346 48580 33348
rect 48300 33294 48302 33346
rect 48354 33294 48580 33346
rect 48300 33292 48580 33294
rect 48300 31892 48356 33292
rect 49084 33234 49140 33246
rect 49084 33182 49086 33234
rect 49138 33182 49140 33234
rect 49084 32786 49140 33182
rect 49084 32734 49086 32786
rect 49138 32734 49140 32786
rect 49084 32722 49140 32734
rect 49196 32788 49252 38220
rect 49308 38050 49364 38062
rect 49308 37998 49310 38050
rect 49362 37998 49364 38050
rect 49308 37828 49364 37998
rect 49756 37828 49812 38668
rect 49308 37826 49812 37828
rect 49308 37774 49758 37826
rect 49810 37774 49812 37826
rect 49308 37772 49812 37774
rect 49308 36482 49364 37772
rect 49756 37762 49812 37772
rect 50316 36596 50372 41132
rect 50652 41094 50708 41132
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50652 39396 50708 39406
rect 50876 39396 50932 45052
rect 51100 44884 51156 46510
rect 52108 46564 52164 48748
rect 53004 48354 53060 48748
rect 53116 48738 53172 48748
rect 53004 48302 53006 48354
rect 53058 48302 53060 48354
rect 53004 48290 53060 48302
rect 52668 47460 52724 47470
rect 52668 47366 52724 47404
rect 53340 46900 53396 52220
rect 53676 52164 53732 52782
rect 53676 52098 53732 52108
rect 54012 52722 54068 52734
rect 54012 52670 54014 52722
rect 54066 52670 54068 52722
rect 54012 50820 54068 52670
rect 54124 52164 54180 52174
rect 54124 52070 54180 52108
rect 54012 50754 54068 50764
rect 54236 50428 54292 53566
rect 54460 52946 54516 54236
rect 54572 54226 54628 54236
rect 54796 54180 54852 56028
rect 54908 56018 54964 56028
rect 55132 55970 55188 55982
rect 55132 55918 55134 55970
rect 55186 55918 55188 55970
rect 54908 55524 54964 55534
rect 54908 55300 54964 55468
rect 55132 55524 55188 55918
rect 55132 55458 55188 55468
rect 55244 55468 55300 56924
rect 55356 56914 55412 56924
rect 55580 56754 55636 56766
rect 55580 56702 55582 56754
rect 55634 56702 55636 56754
rect 55356 56642 55412 56654
rect 55356 56590 55358 56642
rect 55410 56590 55412 56642
rect 55356 55748 55412 56590
rect 55580 55858 55636 56702
rect 55580 55806 55582 55858
rect 55634 55806 55636 55858
rect 55580 55794 55636 55806
rect 55356 55692 55524 55748
rect 55468 55636 55524 55692
rect 55468 55580 55748 55636
rect 55692 55468 55748 55580
rect 55244 55412 55412 55468
rect 55580 55412 55636 55422
rect 55692 55412 55860 55468
rect 55356 55410 55636 55412
rect 55356 55358 55582 55410
rect 55634 55358 55636 55410
rect 55356 55356 55636 55358
rect 55580 55346 55636 55356
rect 55020 55300 55076 55310
rect 54908 55298 55020 55300
rect 54908 55246 54910 55298
rect 54962 55246 55020 55298
rect 54908 55244 55020 55246
rect 54908 55206 54964 55244
rect 54796 53618 54852 54124
rect 54908 54292 54964 54302
rect 54908 53730 54964 54236
rect 54908 53678 54910 53730
rect 54962 53678 54964 53730
rect 54908 53666 54964 53678
rect 54796 53566 54798 53618
rect 54850 53566 54852 53618
rect 54796 53554 54852 53566
rect 55020 53172 55076 55244
rect 55132 54628 55188 54638
rect 55132 54402 55188 54572
rect 55132 54350 55134 54402
rect 55186 54350 55188 54402
rect 55132 54180 55188 54350
rect 55132 54114 55188 54124
rect 55804 54626 55860 55412
rect 55804 54574 55806 54626
rect 55858 54574 55860 54626
rect 55804 53844 55860 54574
rect 56476 55412 56532 55422
rect 56476 54516 56532 55356
rect 56364 54514 56532 54516
rect 56364 54462 56478 54514
rect 56530 54462 56532 54514
rect 56364 54460 56532 54462
rect 55916 54402 55972 54414
rect 56140 54404 56196 54414
rect 55916 54350 55918 54402
rect 55970 54350 55972 54402
rect 55916 53844 55972 54350
rect 56028 54348 56140 54404
rect 56028 54290 56084 54348
rect 56140 54338 56196 54348
rect 56028 54238 56030 54290
rect 56082 54238 56084 54290
rect 56028 54226 56084 54238
rect 56028 53844 56084 53854
rect 55916 53842 56084 53844
rect 55916 53790 56030 53842
rect 56082 53790 56084 53842
rect 55916 53788 56084 53790
rect 55244 53730 55300 53742
rect 55244 53678 55246 53730
rect 55298 53678 55300 53730
rect 55244 53172 55300 53678
rect 55020 53170 55300 53172
rect 55020 53118 55022 53170
rect 55074 53118 55300 53170
rect 55020 53116 55300 53118
rect 55020 53106 55076 53116
rect 54460 52894 54462 52946
rect 54514 52894 54516 52946
rect 54460 52882 54516 52894
rect 54348 52722 54404 52734
rect 54348 52670 54350 52722
rect 54402 52670 54404 52722
rect 54348 51940 54404 52670
rect 55804 52388 55860 53788
rect 56028 53778 56084 53788
rect 56364 53284 56420 54460
rect 56476 54450 56532 54460
rect 56812 54628 56868 54638
rect 56812 54514 56868 54572
rect 56812 54462 56814 54514
rect 56866 54462 56868 54514
rect 56812 54450 56868 54462
rect 57148 54514 57204 54526
rect 57148 54462 57150 54514
rect 57202 54462 57204 54514
rect 56700 54404 56756 54414
rect 56700 54310 56756 54348
rect 57148 54292 57204 54462
rect 57148 54226 57204 54236
rect 56252 53228 56420 53284
rect 55916 52388 55972 52398
rect 55804 52386 55972 52388
rect 55804 52334 55918 52386
rect 55970 52334 55972 52386
rect 55804 52332 55972 52334
rect 55916 52322 55972 52332
rect 56140 52388 56196 52398
rect 56140 52294 56196 52332
rect 56252 52386 56308 53228
rect 56252 52334 56254 52386
rect 56306 52334 56308 52386
rect 55132 52164 55188 52174
rect 56252 52164 56308 52334
rect 56588 52388 56644 52398
rect 56644 52332 56756 52388
rect 56588 52322 56644 52332
rect 54460 51940 54516 51950
rect 54348 51938 54516 51940
rect 54348 51886 54462 51938
rect 54514 51886 54516 51938
rect 54348 51884 54516 51886
rect 54460 51492 54516 51884
rect 54684 51492 54740 51502
rect 54460 51436 54684 51492
rect 54236 50372 54516 50428
rect 54460 49812 54516 50372
rect 54124 49026 54180 49038
rect 54124 48974 54126 49026
rect 54178 48974 54180 49026
rect 53900 48804 53956 48814
rect 54124 48804 54180 48974
rect 54460 49026 54516 49756
rect 54460 48974 54462 49026
rect 54514 48974 54516 49026
rect 54460 48962 54516 48974
rect 53900 48802 54180 48804
rect 53900 48750 53902 48802
rect 53954 48750 54180 48802
rect 53900 48748 54180 48750
rect 54684 48914 54740 51436
rect 55132 51378 55188 52108
rect 55916 52108 56308 52164
rect 55468 51604 55524 51614
rect 55468 51490 55524 51548
rect 55916 51602 55972 52108
rect 56252 51940 56308 51950
rect 55916 51550 55918 51602
rect 55970 51550 55972 51602
rect 55916 51538 55972 51550
rect 56028 51938 56308 51940
rect 56028 51886 56254 51938
rect 56306 51886 56308 51938
rect 56028 51884 56308 51886
rect 55468 51438 55470 51490
rect 55522 51438 55524 51490
rect 55468 51426 55524 51438
rect 55132 51326 55134 51378
rect 55186 51326 55188 51378
rect 55132 51314 55188 51326
rect 55356 51378 55412 51390
rect 55356 51326 55358 51378
rect 55410 51326 55412 51378
rect 55356 51268 55412 51326
rect 55244 50594 55300 50606
rect 55244 50542 55246 50594
rect 55298 50542 55300 50594
rect 55244 50428 55300 50542
rect 54908 50372 54964 50382
rect 55020 50372 55300 50428
rect 55356 50428 55412 51212
rect 56028 50706 56084 51884
rect 56252 51874 56308 51884
rect 56700 51602 56756 52332
rect 56700 51550 56702 51602
rect 56754 51550 56756 51602
rect 56700 51538 56756 51550
rect 57036 51604 57092 51614
rect 56812 51492 56868 51502
rect 56476 51380 56532 51390
rect 56476 51286 56532 51324
rect 56812 51378 56868 51436
rect 56812 51326 56814 51378
rect 56866 51326 56868 51378
rect 56812 51314 56868 51326
rect 57036 51378 57092 51548
rect 57036 51326 57038 51378
rect 57090 51326 57092 51378
rect 57036 51314 57092 51326
rect 56028 50654 56030 50706
rect 56082 50654 56084 50706
rect 56028 50642 56084 50654
rect 57260 50428 57316 60734
rect 57484 60956 57876 61012
rect 57932 61012 57988 61022
rect 57372 59890 57428 59902
rect 57372 59838 57374 59890
rect 57426 59838 57428 59890
rect 57372 59444 57428 59838
rect 57372 59378 57428 59388
rect 57372 52836 57428 52846
rect 57372 52742 57428 52780
rect 55356 50372 55524 50428
rect 54908 50370 55076 50372
rect 54908 50318 54910 50370
rect 54962 50318 55076 50370
rect 54908 50316 55076 50318
rect 54908 50306 54964 50316
rect 54908 49252 54964 49262
rect 54908 49026 54964 49196
rect 54908 48974 54910 49026
rect 54962 48974 54964 49026
rect 54908 48962 54964 48974
rect 55020 49028 55076 50316
rect 55468 49252 55524 50372
rect 57148 50372 57316 50428
rect 55468 49186 55524 49196
rect 56028 49252 56084 49262
rect 56084 49196 56196 49252
rect 56028 49186 56084 49196
rect 55244 49028 55300 49038
rect 55020 49026 55300 49028
rect 55020 48974 55246 49026
rect 55298 48974 55300 49026
rect 55020 48972 55300 48974
rect 54684 48862 54686 48914
rect 54738 48862 54740 48914
rect 53900 48468 53956 48748
rect 54684 48692 54740 48862
rect 54684 48626 54740 48636
rect 54796 48802 54852 48814
rect 54796 48750 54798 48802
rect 54850 48750 54852 48802
rect 53900 48402 53956 48412
rect 54796 48356 54852 48750
rect 54796 48290 54852 48300
rect 53676 48244 53732 48254
rect 54236 48244 54292 48254
rect 53676 48242 54236 48244
rect 53676 48190 53678 48242
rect 53730 48190 54236 48242
rect 53676 48188 54236 48190
rect 53676 47460 53732 48188
rect 54236 48150 54292 48188
rect 54908 48244 54964 48254
rect 55244 48244 55300 48972
rect 56028 48916 56084 48926
rect 55916 48914 56084 48916
rect 55916 48862 56030 48914
rect 56082 48862 56084 48914
rect 55916 48860 56084 48862
rect 55692 48692 55748 48702
rect 55468 48356 55524 48366
rect 55468 48262 55524 48300
rect 55692 48354 55748 48636
rect 55916 48466 55972 48860
rect 56028 48850 56084 48860
rect 55916 48414 55918 48466
rect 55970 48414 55972 48466
rect 55916 48402 55972 48414
rect 55692 48302 55694 48354
rect 55746 48302 55748 48354
rect 55692 48290 55748 48302
rect 54964 48188 55300 48244
rect 56140 48242 56196 49196
rect 56140 48190 56142 48242
rect 56194 48190 56196 48242
rect 54908 48150 54964 48188
rect 56140 48178 56196 48190
rect 56252 48244 56308 48254
rect 56252 47570 56308 48188
rect 56252 47518 56254 47570
rect 56306 47518 56308 47570
rect 56252 47506 56308 47518
rect 53676 47394 53732 47404
rect 53452 47348 53508 47358
rect 53452 47346 53620 47348
rect 53452 47294 53454 47346
rect 53506 47294 53620 47346
rect 53452 47292 53620 47294
rect 53452 47282 53508 47292
rect 52108 46498 52164 46508
rect 52332 46844 53396 46900
rect 53564 46898 53620 47292
rect 53564 46846 53566 46898
rect 53618 46846 53620 46898
rect 51100 44818 51156 44828
rect 51212 45778 51268 45790
rect 51212 45726 51214 45778
rect 51266 45726 51268 45778
rect 51212 44546 51268 45726
rect 51884 44996 51940 45006
rect 51212 44494 51214 44546
rect 51266 44494 51268 44546
rect 51212 44482 51268 44494
rect 51436 44884 51492 44894
rect 50988 40292 51044 40302
rect 50988 40290 51380 40292
rect 50988 40238 50990 40290
rect 51042 40238 51380 40290
rect 50988 40236 51380 40238
rect 50988 40226 51044 40236
rect 51324 39842 51380 40236
rect 51324 39790 51326 39842
rect 51378 39790 51380 39842
rect 51324 39778 51380 39790
rect 50652 39394 50932 39396
rect 50652 39342 50654 39394
rect 50706 39342 50932 39394
rect 50652 39340 50932 39342
rect 50652 39330 50708 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50876 38724 50932 39340
rect 50988 39730 51044 39742
rect 50988 39678 50990 39730
rect 51042 39678 51044 39730
rect 50988 38946 51044 39678
rect 50988 38894 50990 38946
rect 51042 38894 51044 38946
rect 50988 38882 51044 38894
rect 51100 39394 51156 39406
rect 51100 39342 51102 39394
rect 51154 39342 51156 39394
rect 51100 38724 51156 39342
rect 50876 38668 51156 38724
rect 51436 38668 51492 44828
rect 51772 44434 51828 44446
rect 51772 44382 51774 44434
rect 51826 44382 51828 44434
rect 51772 43764 51828 44382
rect 51548 43708 51772 43764
rect 51548 42754 51604 43708
rect 51772 43698 51828 43708
rect 51884 44322 51940 44940
rect 51884 44270 51886 44322
rect 51938 44270 51940 44322
rect 51548 42702 51550 42754
rect 51602 42702 51604 42754
rect 51548 41074 51604 42702
rect 51660 42866 51716 42878
rect 51660 42814 51662 42866
rect 51714 42814 51716 42866
rect 51660 42644 51716 42814
rect 51772 42756 51828 42766
rect 51884 42756 51940 44270
rect 51772 42754 51940 42756
rect 51772 42702 51774 42754
rect 51826 42702 51940 42754
rect 51772 42700 51940 42702
rect 51772 42690 51828 42700
rect 51660 41860 51716 42588
rect 51660 41804 51828 41860
rect 51660 41188 51716 41198
rect 51660 41094 51716 41132
rect 51548 41022 51550 41074
rect 51602 41022 51604 41074
rect 51548 41010 51604 41022
rect 51660 40404 51716 40414
rect 51660 40310 51716 40348
rect 51772 40290 51828 41804
rect 51884 41412 51940 42700
rect 51884 41186 51940 41356
rect 51884 41134 51886 41186
rect 51938 41134 51940 41186
rect 51884 41122 51940 41134
rect 51996 42530 52052 42542
rect 51996 42478 51998 42530
rect 52050 42478 52052 42530
rect 51996 41858 52052 42478
rect 51996 41806 51998 41858
rect 52050 41806 52052 41858
rect 51996 41300 52052 41806
rect 51996 41186 52052 41244
rect 51996 41134 51998 41186
rect 52050 41134 52052 41186
rect 51996 41122 52052 41134
rect 51772 40238 51774 40290
rect 51826 40238 51828 40290
rect 51772 40226 51828 40238
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 49308 36430 49310 36482
rect 49362 36430 49364 36482
rect 49308 36418 49364 36430
rect 50204 36540 50372 36596
rect 49980 36372 50036 36382
rect 49980 36278 50036 36316
rect 50092 35476 50148 35486
rect 49980 35028 50036 35038
rect 49980 34934 50036 34972
rect 49420 34802 49476 34814
rect 49420 34750 49422 34802
rect 49474 34750 49476 34802
rect 49420 33460 49476 34750
rect 49532 34804 49588 34814
rect 50092 34804 50148 35420
rect 49532 34802 50148 34804
rect 49532 34750 49534 34802
rect 49586 34750 50148 34802
rect 49532 34748 50148 34750
rect 49532 34738 49588 34748
rect 49420 33394 49476 33404
rect 49196 32732 49812 32788
rect 48972 32564 49028 32574
rect 48972 32470 49028 32508
rect 49196 32562 49252 32574
rect 49196 32510 49198 32562
rect 49250 32510 49252 32562
rect 49084 32228 49140 32238
rect 48748 31892 48804 31902
rect 48300 31890 48804 31892
rect 48300 31838 48750 31890
rect 48802 31838 48804 31890
rect 48300 31836 48804 31838
rect 48300 31778 48356 31836
rect 48748 31826 48804 31836
rect 48300 31726 48302 31778
rect 48354 31726 48356 31778
rect 48300 30660 48356 31726
rect 49084 31218 49140 32172
rect 49196 31780 49252 32510
rect 49644 32564 49700 32574
rect 49644 32470 49700 32508
rect 49532 32228 49588 32238
rect 49308 31780 49364 31790
rect 49196 31724 49308 31780
rect 49308 31686 49364 31724
rect 49532 31778 49588 32172
rect 49532 31726 49534 31778
rect 49586 31726 49588 31778
rect 49532 31714 49588 31726
rect 49420 31668 49476 31678
rect 49420 31574 49476 31612
rect 49756 31556 49812 32732
rect 49084 31166 49086 31218
rect 49138 31166 49140 31218
rect 49084 31154 49140 31166
rect 49532 31500 49812 31556
rect 49868 32002 49924 32014
rect 49868 31950 49870 32002
rect 49922 31950 49924 32002
rect 48412 30660 48468 30670
rect 48300 30604 48412 30660
rect 48412 30594 48468 30604
rect 49084 30098 49140 30110
rect 49084 30046 49086 30098
rect 49138 30046 49140 30098
rect 49084 29652 49140 30046
rect 49084 29586 49140 29596
rect 49532 28868 49588 31500
rect 49868 30882 49924 31950
rect 50092 31892 50148 31902
rect 50092 31778 50148 31836
rect 50092 31726 50094 31778
rect 50146 31726 50148 31778
rect 50092 31714 50148 31726
rect 49868 30830 49870 30882
rect 49922 30830 49924 30882
rect 49868 30818 49924 30830
rect 49980 31106 50036 31118
rect 50204 31108 50260 36540
rect 50316 36372 50372 36382
rect 50372 36316 50484 36372
rect 50316 36306 50372 36316
rect 50428 35922 50484 36316
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50428 35870 50430 35922
rect 50482 35870 50484 35922
rect 50428 35858 50484 35870
rect 50652 35698 50708 35710
rect 50652 35646 50654 35698
rect 50706 35646 50708 35698
rect 50316 35476 50372 35486
rect 50652 35476 50708 35646
rect 50876 35476 50932 35486
rect 50652 35474 50932 35476
rect 50652 35422 50878 35474
rect 50930 35422 50932 35474
rect 50652 35420 50932 35422
rect 50316 35382 50372 35420
rect 50876 35410 50932 35420
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 51100 34356 51156 38668
rect 51212 38612 51492 38668
rect 51212 35922 51268 38612
rect 51212 35870 51214 35922
rect 51266 35870 51268 35922
rect 51212 35474 51268 35870
rect 52108 36594 52164 36606
rect 52108 36542 52110 36594
rect 52162 36542 52164 36594
rect 51996 35812 52052 35822
rect 52108 35812 52164 36542
rect 51996 35810 52164 35812
rect 51996 35758 51998 35810
rect 52050 35758 52164 35810
rect 51996 35756 52164 35758
rect 51996 35746 52052 35756
rect 52108 35700 52164 35756
rect 52220 35700 52276 35710
rect 52108 35644 52220 35700
rect 52220 35634 52276 35644
rect 51996 35586 52052 35598
rect 51996 35534 51998 35586
rect 52050 35534 52052 35586
rect 51212 35422 51214 35474
rect 51266 35422 51268 35474
rect 51212 35410 51268 35422
rect 51772 35476 51828 35486
rect 51772 35382 51828 35420
rect 51100 34290 51156 34300
rect 51212 33460 51268 33470
rect 51996 33460 52052 35534
rect 51212 33458 51716 33460
rect 51212 33406 51214 33458
rect 51266 33406 51716 33458
rect 51212 33404 51716 33406
rect 51996 33404 52276 33460
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51212 32788 51268 33404
rect 50652 32732 51268 32788
rect 51548 33234 51604 33246
rect 51548 33182 51550 33234
rect 51602 33182 51604 33234
rect 50652 32674 50708 32732
rect 50652 32622 50654 32674
rect 50706 32622 50708 32674
rect 50652 32610 50708 32622
rect 50316 32562 50372 32574
rect 50316 32510 50318 32562
rect 50370 32510 50372 32562
rect 50316 31948 50372 32510
rect 50428 32564 50484 32574
rect 50428 32470 50484 32508
rect 50876 32562 50932 32574
rect 50876 32510 50878 32562
rect 50930 32510 50932 32562
rect 50316 31892 50484 31948
rect 49980 31054 49982 31106
rect 50034 31054 50036 31106
rect 49868 30660 49924 30670
rect 49868 30212 49924 30604
rect 49980 30324 50036 31054
rect 49980 30258 50036 30268
rect 50092 31052 50260 31108
rect 50428 31780 50484 31892
rect 50876 31892 50932 32510
rect 51436 32450 51492 32462
rect 51436 32398 51438 32450
rect 51490 32398 51492 32450
rect 51436 32116 51492 32398
rect 51436 32050 51492 32060
rect 51548 31892 51604 33182
rect 51660 32564 51716 33404
rect 51884 33348 51940 33358
rect 51884 33254 51940 33292
rect 51996 33236 52052 33246
rect 51996 33142 52052 33180
rect 52108 33234 52164 33246
rect 52108 33182 52110 33234
rect 52162 33182 52164 33234
rect 52108 32900 52164 33182
rect 51772 32844 52164 32900
rect 51772 32786 51828 32844
rect 51772 32734 51774 32786
rect 51826 32734 51828 32786
rect 51772 32722 51828 32734
rect 51996 32674 52052 32686
rect 51996 32622 51998 32674
rect 52050 32622 52052 32674
rect 51996 32564 52052 32622
rect 52108 32676 52164 32686
rect 52220 32676 52276 33404
rect 52108 32674 52220 32676
rect 52108 32622 52110 32674
rect 52162 32622 52220 32674
rect 52108 32620 52220 32622
rect 52108 32610 52164 32620
rect 52220 32582 52276 32620
rect 51660 32508 52052 32564
rect 51772 31892 51828 31902
rect 51548 31836 51772 31892
rect 50876 31826 50932 31836
rect 50428 31554 50484 31724
rect 50428 31502 50430 31554
rect 50482 31502 50484 31554
rect 49868 30118 49924 30156
rect 50092 30100 50148 31052
rect 50204 30884 50260 30894
rect 50204 30790 50260 30828
rect 50428 30660 50484 31502
rect 50764 31556 50820 31594
rect 50820 31500 50932 31556
rect 50764 31490 50820 31500
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50876 30884 50932 31500
rect 50876 30818 50932 30828
rect 50204 30604 50484 30660
rect 50204 30210 50260 30604
rect 51548 30436 51604 30446
rect 50204 30158 50206 30210
rect 50258 30158 50260 30210
rect 50204 30146 50260 30158
rect 50316 30324 50372 30334
rect 48524 28756 48580 28766
rect 48524 28662 48580 28700
rect 49532 28754 49588 28812
rect 49980 30044 50148 30100
rect 50316 30098 50372 30268
rect 50316 30046 50318 30098
rect 50370 30046 50372 30098
rect 49532 28702 49534 28754
rect 49586 28702 49588 28754
rect 49532 28690 49588 28702
rect 49756 28756 49812 28766
rect 49756 28662 49812 28700
rect 48188 26292 48244 26302
rect 47628 26290 48244 26292
rect 47628 26238 47630 26290
rect 47682 26238 48190 26290
rect 48242 26238 48244 26290
rect 47628 26236 48244 26238
rect 47628 26226 47684 26236
rect 48188 26226 48244 26236
rect 47292 26066 47348 26078
rect 47292 26014 47294 26066
rect 47346 26014 47348 26066
rect 46620 25620 46676 25630
rect 46620 25526 46676 25564
rect 46956 25618 47012 25630
rect 46956 25566 46958 25618
rect 47010 25566 47012 25618
rect 45948 25508 46004 25518
rect 45948 25414 46004 25452
rect 46956 25508 47012 25566
rect 47292 25620 47348 26014
rect 47628 26068 47684 26078
rect 47628 25974 47684 26012
rect 49084 26068 49140 26078
rect 47292 25554 47348 25564
rect 49084 25618 49140 26012
rect 49980 25844 50036 30044
rect 50316 30034 50372 30046
rect 50876 30212 50932 30222
rect 50876 30100 50932 30156
rect 51548 30212 51604 30380
rect 51772 30324 51828 31836
rect 52332 31220 52388 46844
rect 53564 46834 53620 46846
rect 55692 47234 55748 47246
rect 55692 47182 55694 47234
rect 55746 47182 55748 47234
rect 53340 46674 53396 46686
rect 53340 46622 53342 46674
rect 53394 46622 53396 46674
rect 53004 46564 53060 46574
rect 53340 46564 53396 46622
rect 53676 46676 53732 46686
rect 54124 46676 54180 46686
rect 53676 46674 54180 46676
rect 53676 46622 53678 46674
rect 53730 46622 54126 46674
rect 54178 46622 54180 46674
rect 53676 46620 54180 46622
rect 53676 46610 53732 46620
rect 54124 46610 54180 46620
rect 55020 46674 55076 46686
rect 55020 46622 55022 46674
rect 55074 46622 55076 46674
rect 53004 46562 53396 46564
rect 53004 46510 53006 46562
rect 53058 46510 53396 46562
rect 53004 46508 53396 46510
rect 54796 46564 54852 46574
rect 53004 46452 53060 46508
rect 54796 46470 54852 46508
rect 53004 46386 53060 46396
rect 54908 45892 54964 45902
rect 53340 45332 53396 45342
rect 54908 45332 54964 45836
rect 53340 45238 53396 45276
rect 54796 45276 54908 45332
rect 52892 44996 52948 45006
rect 52892 44902 52948 44940
rect 54572 44548 54628 44558
rect 54572 44454 54628 44492
rect 54236 44436 54292 44446
rect 53676 44434 54292 44436
rect 53676 44382 54238 44434
rect 54290 44382 54292 44434
rect 53676 44380 54292 44382
rect 53564 43652 53620 43662
rect 52780 43540 52836 43550
rect 52780 43446 52836 43484
rect 53228 43540 53284 43550
rect 53228 43446 53284 43484
rect 53116 42980 53172 42990
rect 53116 42866 53172 42924
rect 53564 42978 53620 43596
rect 53564 42926 53566 42978
rect 53618 42926 53620 42978
rect 53564 42914 53620 42926
rect 53676 42978 53732 44380
rect 54236 44370 54292 44380
rect 54348 44100 54404 44110
rect 54348 44006 54404 44044
rect 54796 43426 54852 45276
rect 54908 45266 54964 45276
rect 55020 45108 55076 46622
rect 55692 46564 55748 47182
rect 55804 46564 55860 46574
rect 55692 46508 55804 46564
rect 55244 46004 55300 46014
rect 55244 46002 55412 46004
rect 55244 45950 55246 46002
rect 55298 45950 55412 46002
rect 55244 45948 55412 45950
rect 55244 45938 55300 45948
rect 55020 45042 55076 45052
rect 55132 45220 55188 45230
rect 55132 44884 55188 45164
rect 54908 44098 54964 44110
rect 54908 44046 54910 44098
rect 54962 44046 54964 44098
rect 54908 43764 54964 44046
rect 54908 43698 54964 43708
rect 54796 43374 54798 43426
rect 54850 43374 54852 43426
rect 53676 42926 53678 42978
rect 53730 42926 53732 42978
rect 53676 42914 53732 42926
rect 53900 42980 53956 42990
rect 53900 42886 53956 42924
rect 53116 42814 53118 42866
rect 53170 42814 53172 42866
rect 53116 42802 53172 42814
rect 54012 42642 54068 42654
rect 54012 42590 54014 42642
rect 54066 42590 54068 42642
rect 54012 42196 54068 42590
rect 53788 42140 54068 42196
rect 53788 42082 53844 42140
rect 53788 42030 53790 42082
rect 53842 42030 53844 42082
rect 53788 42018 53844 42030
rect 52444 41972 52500 41982
rect 52444 41878 52500 41916
rect 53116 41972 53172 41982
rect 53116 41878 53172 41916
rect 53676 41972 53732 41982
rect 52892 41412 52948 41422
rect 52892 41318 52948 41356
rect 52668 41300 52724 41310
rect 52668 41206 52724 41244
rect 53116 41186 53172 41198
rect 53116 41134 53118 41186
rect 53170 41134 53172 41186
rect 53116 40404 53172 41134
rect 53564 40964 53620 40974
rect 53564 40870 53620 40908
rect 53116 38722 53172 40348
rect 53676 39620 53732 41916
rect 54796 41972 54852 43374
rect 55132 42980 55188 44828
rect 55356 45108 55412 45948
rect 55468 45108 55524 45118
rect 55356 45106 55524 45108
rect 55356 45054 55470 45106
rect 55522 45054 55524 45106
rect 55356 45052 55524 45054
rect 55244 44548 55300 44558
rect 55244 44454 55300 44492
rect 55132 42914 55188 42924
rect 55356 44324 55412 45052
rect 55468 45042 55524 45052
rect 55692 45108 55748 45118
rect 55804 45108 55860 46508
rect 57148 45892 57204 50372
rect 57036 45836 57204 45892
rect 55916 45332 55972 45342
rect 55916 45330 56868 45332
rect 55916 45278 55918 45330
rect 55970 45278 56868 45330
rect 55916 45276 56868 45278
rect 55916 45266 55972 45276
rect 56028 45108 56084 45118
rect 56588 45108 56644 45118
rect 55804 45106 56084 45108
rect 55804 45054 56030 45106
rect 56082 45054 56084 45106
rect 55804 45052 56084 45054
rect 55356 42644 55412 44268
rect 55468 44322 55524 44334
rect 55468 44270 55470 44322
rect 55522 44270 55524 44322
rect 55468 44100 55524 44270
rect 55468 43764 55524 44044
rect 55692 43988 55748 45052
rect 56028 44100 56084 45052
rect 56140 45106 56644 45108
rect 56140 45054 56590 45106
rect 56642 45054 56644 45106
rect 56140 45052 56644 45054
rect 56140 44548 56196 45052
rect 56588 45042 56644 45052
rect 56812 45106 56868 45276
rect 56812 45054 56814 45106
rect 56866 45054 56868 45106
rect 56812 45042 56868 45054
rect 57036 45220 57092 45836
rect 57372 45780 57428 45790
rect 57036 45106 57092 45164
rect 57148 45778 57428 45780
rect 57148 45726 57374 45778
rect 57426 45726 57428 45778
rect 57148 45724 57428 45726
rect 57148 45218 57204 45724
rect 57372 45714 57428 45724
rect 57148 45166 57150 45218
rect 57202 45166 57204 45218
rect 57148 45154 57204 45166
rect 57036 45054 57038 45106
rect 57090 45054 57092 45106
rect 57036 45042 57092 45054
rect 56140 44454 56196 44492
rect 57484 44436 57540 60956
rect 57932 60918 57988 60956
rect 57820 60676 57876 60686
rect 57820 60582 57876 60620
rect 57708 60564 57764 60574
rect 57708 60470 57764 60508
rect 58044 60004 58100 60014
rect 58156 60004 58212 63086
rect 58100 59948 58212 60004
rect 58044 59910 58100 59948
rect 58156 59220 58212 59230
rect 57708 59108 57764 59118
rect 57708 59106 57876 59108
rect 57708 59054 57710 59106
rect 57762 59054 57876 59106
rect 57708 59052 57876 59054
rect 57708 59042 57764 59052
rect 57708 55410 57764 55422
rect 57708 55358 57710 55410
rect 57762 55358 57764 55410
rect 57708 54628 57764 55358
rect 57708 54562 57764 54572
rect 57596 52834 57652 52846
rect 57596 52782 57598 52834
rect 57650 52782 57652 52834
rect 57596 52276 57652 52782
rect 57596 52210 57652 52220
rect 57708 44994 57764 45006
rect 57708 44942 57710 44994
rect 57762 44942 57764 44994
rect 57596 44436 57652 44446
rect 57372 44434 57652 44436
rect 57372 44382 57598 44434
rect 57650 44382 57652 44434
rect 57372 44380 57652 44382
rect 56588 44324 56644 44334
rect 56588 44230 56644 44268
rect 56700 44210 56756 44222
rect 56700 44158 56702 44210
rect 56754 44158 56756 44210
rect 56700 44100 56756 44158
rect 56028 44044 56756 44100
rect 55692 43922 55748 43932
rect 56364 43764 56420 43774
rect 55468 43708 55972 43764
rect 55916 42754 55972 43708
rect 55916 42702 55918 42754
rect 55970 42702 55972 42754
rect 55468 42644 55524 42654
rect 55356 42642 55524 42644
rect 55356 42590 55470 42642
rect 55522 42590 55524 42642
rect 55356 42588 55524 42590
rect 55468 42578 55524 42588
rect 54796 41906 54852 41916
rect 55356 41860 55412 41870
rect 55356 41074 55412 41804
rect 55916 41858 55972 42702
rect 55916 41806 55918 41858
rect 55970 41806 55972 41858
rect 55916 41794 55972 41806
rect 56252 41972 56308 41982
rect 55356 41022 55358 41074
rect 55410 41022 55412 41074
rect 55356 41010 55412 41022
rect 55692 41186 55748 41198
rect 55692 41134 55694 41186
rect 55746 41134 55748 41186
rect 55692 40626 55748 41134
rect 55692 40574 55694 40626
rect 55746 40574 55748 40626
rect 55692 40562 55748 40574
rect 55804 41132 56084 41188
rect 53564 39618 53732 39620
rect 53564 39566 53678 39618
rect 53730 39566 53732 39618
rect 53564 39564 53732 39566
rect 53564 39060 53620 39564
rect 53676 39554 53732 39564
rect 54348 39508 54404 39518
rect 54236 39506 54404 39508
rect 54236 39454 54350 39506
rect 54402 39454 54404 39506
rect 54236 39452 54404 39454
rect 53116 38670 53118 38722
rect 53170 38670 53172 38722
rect 53116 38658 53172 38670
rect 53340 39058 53620 39060
rect 53340 39006 53566 39058
rect 53618 39006 53620 39058
rect 53340 39004 53620 39006
rect 52892 36596 52948 36606
rect 53340 36596 53396 39004
rect 53564 38994 53620 39004
rect 54124 39060 54180 39070
rect 54124 38966 54180 39004
rect 53676 38724 53732 38734
rect 53900 38724 53956 38734
rect 53732 38722 53956 38724
rect 53732 38670 53902 38722
rect 53954 38670 53956 38722
rect 53732 38668 53956 38670
rect 53564 37828 53620 37838
rect 53676 37828 53732 38668
rect 53900 38658 53956 38668
rect 54236 38722 54292 39452
rect 54348 39442 54404 39452
rect 54236 38670 54238 38722
rect 54290 38670 54292 38722
rect 54236 38658 54292 38670
rect 55804 38668 55860 41132
rect 55916 40964 55972 40974
rect 55916 40626 55972 40908
rect 56028 40962 56084 41132
rect 56028 40910 56030 40962
rect 56082 40910 56084 40962
rect 56028 40898 56084 40910
rect 55916 40574 55918 40626
rect 55970 40574 55972 40626
rect 55916 40562 55972 40574
rect 56028 40402 56084 40414
rect 56028 40350 56030 40402
rect 56082 40350 56084 40402
rect 56028 40292 56084 40350
rect 56028 40226 56084 40236
rect 56252 38668 56308 41916
rect 56364 39060 56420 43708
rect 56476 42756 56532 42766
rect 56700 42756 56756 44044
rect 56812 44210 56868 44222
rect 56812 44158 56814 44210
rect 56866 44158 56868 44210
rect 56812 43764 56868 44158
rect 56812 43698 56868 43708
rect 57372 43650 57428 44380
rect 57596 44370 57652 44380
rect 57372 43598 57374 43650
rect 57426 43598 57428 43650
rect 57372 43586 57428 43598
rect 57148 43426 57204 43438
rect 57148 43374 57150 43426
rect 57202 43374 57204 43426
rect 56476 42754 56756 42756
rect 56476 42702 56478 42754
rect 56530 42702 56756 42754
rect 56476 42700 56756 42702
rect 57036 42866 57092 42878
rect 57036 42814 57038 42866
rect 57090 42814 57092 42866
rect 56476 42690 56532 42700
rect 56924 42642 56980 42654
rect 56924 42590 56926 42642
rect 56978 42590 56980 42642
rect 56700 41972 56756 41982
rect 56700 41878 56756 41916
rect 56924 41188 56980 42590
rect 57036 42082 57092 42814
rect 57036 42030 57038 42082
rect 57090 42030 57092 42082
rect 57036 41860 57092 42030
rect 57148 41972 57204 43374
rect 57596 43314 57652 43326
rect 57596 43262 57598 43314
rect 57650 43262 57652 43314
rect 57596 42082 57652 43262
rect 57596 42030 57598 42082
rect 57650 42030 57652 42082
rect 57372 41972 57428 41982
rect 57148 41970 57428 41972
rect 57148 41918 57374 41970
rect 57426 41918 57428 41970
rect 57148 41916 57428 41918
rect 57036 41794 57092 41804
rect 56812 41132 56980 41188
rect 57260 41748 57316 41758
rect 56812 39844 56868 41132
rect 57260 41074 57316 41692
rect 57372 41524 57428 41916
rect 57484 41860 57540 41870
rect 57484 41766 57540 41804
rect 57596 41748 57652 42030
rect 57596 41682 57652 41692
rect 57372 41458 57428 41468
rect 57260 41022 57262 41074
rect 57314 41022 57316 41074
rect 57260 41010 57316 41022
rect 57596 41300 57652 41310
rect 57596 41186 57652 41244
rect 57596 41134 57598 41186
rect 57650 41134 57652 41186
rect 56924 40964 56980 40974
rect 56924 40514 56980 40908
rect 56924 40462 56926 40514
rect 56978 40462 56980 40514
rect 56924 40450 56980 40462
rect 57036 40402 57092 40414
rect 57036 40350 57038 40402
rect 57090 40350 57092 40402
rect 57036 40292 57092 40350
rect 57484 40404 57540 40414
rect 57484 40310 57540 40348
rect 57036 39844 57092 40236
rect 57260 40290 57316 40302
rect 57260 40238 57262 40290
rect 57314 40238 57316 40290
rect 57260 40068 57316 40238
rect 57484 40068 57540 40078
rect 57260 40012 57484 40068
rect 57484 40002 57540 40012
rect 57484 39844 57540 39854
rect 56476 39788 56980 39844
rect 57036 39842 57540 39844
rect 57036 39790 57486 39842
rect 57538 39790 57540 39842
rect 57036 39788 57540 39790
rect 56476 39730 56532 39788
rect 56476 39678 56478 39730
rect 56530 39678 56532 39730
rect 56476 39666 56532 39678
rect 56924 39620 56980 39788
rect 57484 39778 57540 39788
rect 57036 39620 57092 39630
rect 56924 39618 57092 39620
rect 56924 39566 57038 39618
rect 57090 39566 57092 39618
rect 56924 39564 57092 39566
rect 57036 39554 57092 39564
rect 57596 39506 57652 41134
rect 57596 39454 57598 39506
rect 57650 39454 57652 39506
rect 57596 39442 57652 39454
rect 56364 38994 56420 39004
rect 56812 39394 56868 39406
rect 56812 39342 56814 39394
rect 56866 39342 56868 39394
rect 56812 39060 56868 39342
rect 56812 38994 56868 39004
rect 57596 38836 57652 38846
rect 57596 38742 57652 38780
rect 56700 38722 56756 38734
rect 56700 38670 56702 38722
rect 56754 38670 56756 38722
rect 56700 38668 56756 38670
rect 55804 38612 55972 38668
rect 56252 38612 56756 38668
rect 54908 38052 54964 38062
rect 54908 37958 54964 37996
rect 55356 38052 55412 38062
rect 55356 37958 55412 37996
rect 53564 37826 53732 37828
rect 53564 37774 53566 37826
rect 53618 37774 53732 37826
rect 53564 37772 53732 37774
rect 53564 37762 53620 37772
rect 52892 36594 53396 36596
rect 52892 36542 52894 36594
rect 52946 36542 53396 36594
rect 52892 36540 53396 36542
rect 52892 36530 52948 36540
rect 53340 36482 53396 36540
rect 53340 36430 53342 36482
rect 53394 36430 53396 36482
rect 53340 36418 53396 36430
rect 52892 35700 52948 35710
rect 52892 35606 52948 35644
rect 53116 35476 53172 35486
rect 53452 35476 53508 35486
rect 53116 35382 53172 35420
rect 53228 35474 53508 35476
rect 53228 35422 53454 35474
rect 53506 35422 53508 35474
rect 53228 35420 53508 35422
rect 53228 34914 53284 35420
rect 53452 35410 53508 35420
rect 53228 34862 53230 34914
rect 53282 34862 53284 34914
rect 52780 33346 52836 33358
rect 52780 33294 52782 33346
rect 52834 33294 52836 33346
rect 52668 32676 52724 32686
rect 52332 31154 52388 31164
rect 52556 32620 52668 32676
rect 51548 30210 51716 30212
rect 51548 30158 51550 30210
rect 51602 30158 51716 30210
rect 51548 30156 51716 30158
rect 51548 30146 51604 30156
rect 50876 30044 51380 30100
rect 50540 29988 50596 29998
rect 50540 29986 51268 29988
rect 50540 29934 50542 29986
rect 50594 29934 51268 29986
rect 50540 29932 51268 29934
rect 50540 29922 50596 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 51100 29652 51156 29662
rect 51100 29558 51156 29596
rect 50988 29428 51044 29438
rect 50988 29334 51044 29372
rect 51212 29426 51268 29932
rect 51212 29374 51214 29426
rect 51266 29374 51268 29426
rect 51212 29362 51268 29374
rect 50652 28868 50708 28878
rect 50652 28754 50708 28812
rect 50652 28702 50654 28754
rect 50706 28702 50708 28754
rect 50652 28690 50708 28702
rect 51324 28756 51380 30044
rect 51548 29540 51604 29550
rect 51548 29446 51604 29484
rect 51436 28756 51492 28766
rect 51324 28700 51436 28756
rect 50092 28418 50148 28430
rect 50092 28366 50094 28418
rect 50146 28366 50148 28418
rect 50092 28084 50148 28366
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50092 28018 50148 28028
rect 49980 25778 50036 25788
rect 50316 27860 50372 27870
rect 50316 25620 50372 27804
rect 51436 27860 51492 28700
rect 51660 28084 51716 30156
rect 51772 30098 51828 30268
rect 51772 30046 51774 30098
rect 51826 30046 51828 30098
rect 51772 30034 51828 30046
rect 52556 28644 52612 32620
rect 52668 32610 52724 32620
rect 52780 32116 52836 33294
rect 52892 32676 52948 32686
rect 52892 32674 53172 32676
rect 52892 32622 52894 32674
rect 52946 32622 53172 32674
rect 52892 32620 53172 32622
rect 52892 32610 52948 32620
rect 52780 32050 52836 32060
rect 53116 31556 53172 32620
rect 53228 32674 53284 34862
rect 53452 34692 53508 34702
rect 53452 34598 53508 34636
rect 53452 33236 53508 33246
rect 53452 33142 53508 33180
rect 53228 32622 53230 32674
rect 53282 32622 53284 32674
rect 53228 32610 53284 32622
rect 52668 30324 52724 30334
rect 52668 30210 52724 30268
rect 52668 30158 52670 30210
rect 52722 30158 52724 30210
rect 52668 30146 52724 30158
rect 53004 29986 53060 29998
rect 53004 29934 53006 29986
rect 53058 29934 53060 29986
rect 53004 29540 53060 29934
rect 53116 29652 53172 31500
rect 53228 29988 53284 29998
rect 53228 29652 53284 29932
rect 53116 29650 53284 29652
rect 53116 29598 53118 29650
rect 53170 29598 53284 29650
rect 53116 29596 53284 29598
rect 53116 29586 53172 29596
rect 53452 29540 53508 29550
rect 53004 28756 53060 29484
rect 53340 29538 53508 29540
rect 53340 29486 53454 29538
rect 53506 29486 53508 29538
rect 53340 29484 53508 29486
rect 53228 29428 53284 29438
rect 53004 28700 53172 28756
rect 52668 28644 52724 28654
rect 52556 28642 52724 28644
rect 52556 28590 52670 28642
rect 52722 28590 52724 28642
rect 52556 28588 52724 28590
rect 51660 28018 51716 28028
rect 52668 27972 52724 28588
rect 52668 27906 52724 27916
rect 52780 28532 52836 28542
rect 52780 27860 52836 28476
rect 53004 28532 53060 28542
rect 53004 28438 53060 28476
rect 53116 28420 53172 28700
rect 53228 28642 53284 29372
rect 53228 28590 53230 28642
rect 53282 28590 53284 28642
rect 53228 28578 53284 28590
rect 53116 28364 53284 28420
rect 52780 27804 52948 27860
rect 51436 27766 51492 27804
rect 52108 27748 52164 27758
rect 52108 27746 52836 27748
rect 52108 27694 52110 27746
rect 52162 27694 52836 27746
rect 52108 27692 52836 27694
rect 52108 27682 52164 27692
rect 52780 27186 52836 27692
rect 52780 27134 52782 27186
rect 52834 27134 52836 27186
rect 52780 27122 52836 27134
rect 52556 27074 52612 27086
rect 52556 27022 52558 27074
rect 52610 27022 52612 27074
rect 52556 26908 52612 27022
rect 52892 26908 52948 27804
rect 53228 27074 53284 28364
rect 53340 27860 53396 29484
rect 53452 29474 53508 29484
rect 53564 28532 53620 28542
rect 53564 28438 53620 28476
rect 53340 27794 53396 27804
rect 53452 28418 53508 28430
rect 53452 28366 53454 28418
rect 53506 28366 53508 28418
rect 53452 27748 53508 28366
rect 53676 28308 53732 37772
rect 54012 36372 54068 36382
rect 55580 36372 55636 36382
rect 54012 36370 55188 36372
rect 54012 36318 54014 36370
rect 54066 36318 55188 36370
rect 54012 36316 55188 36318
rect 54012 36306 54068 36316
rect 55132 35922 55188 36316
rect 55132 35870 55134 35922
rect 55186 35870 55188 35922
rect 55132 35858 55188 35870
rect 54908 35700 54964 35710
rect 54684 35698 54964 35700
rect 54684 35646 54910 35698
rect 54962 35646 54964 35698
rect 54684 35644 54964 35646
rect 54012 35364 54068 35374
rect 54012 34692 54068 35308
rect 53788 33348 53844 33358
rect 53788 32340 53844 33292
rect 54012 33236 54068 34636
rect 54684 34354 54740 35644
rect 54908 35634 54964 35644
rect 55356 35700 55412 35710
rect 55356 35606 55412 35644
rect 55580 35698 55636 36316
rect 55580 35646 55582 35698
rect 55634 35646 55636 35698
rect 54684 34302 54686 34354
rect 54738 34302 54740 34354
rect 54684 34290 54740 34302
rect 53900 32788 53956 32798
rect 53900 32694 53956 32732
rect 54012 32674 54068 33180
rect 54908 34242 54964 34254
rect 54908 34190 54910 34242
rect 54962 34190 54964 34242
rect 54908 32788 54964 34190
rect 55020 34130 55076 34142
rect 55020 34078 55022 34130
rect 55074 34078 55076 34130
rect 55020 33348 55076 34078
rect 55580 34132 55636 35646
rect 55580 34066 55636 34076
rect 55020 32788 55076 33292
rect 55580 33458 55636 33470
rect 55580 33406 55582 33458
rect 55634 33406 55636 33458
rect 55132 32788 55188 32798
rect 55020 32786 55188 32788
rect 55020 32734 55134 32786
rect 55186 32734 55188 32786
rect 55020 32732 55188 32734
rect 54908 32722 54964 32732
rect 55132 32722 55188 32732
rect 55580 32788 55636 33406
rect 55580 32722 55636 32732
rect 54012 32622 54014 32674
rect 54066 32622 54068 32674
rect 54012 32610 54068 32622
rect 54796 32676 54852 32686
rect 54796 32582 54852 32620
rect 53900 32340 53956 32350
rect 53788 32338 53956 32340
rect 53788 32286 53902 32338
rect 53954 32286 53956 32338
rect 53788 32284 53956 32286
rect 53900 32274 53956 32284
rect 55244 32116 55300 32126
rect 55244 31778 55300 32060
rect 55244 31726 55246 31778
rect 55298 31726 55300 31778
rect 55132 30994 55188 31006
rect 55132 30942 55134 30994
rect 55186 30942 55188 30994
rect 55132 30436 55188 30942
rect 54572 29988 54628 29998
rect 54572 29894 54628 29932
rect 54908 29988 54964 29998
rect 54908 29894 54964 29932
rect 53900 29314 53956 29326
rect 53900 29262 53902 29314
rect 53954 29262 53956 29314
rect 53900 28644 53956 29262
rect 54460 28644 54516 28654
rect 53900 28642 54516 28644
rect 53900 28590 54462 28642
rect 54514 28590 54516 28642
rect 53900 28588 54516 28590
rect 53452 27682 53508 27692
rect 53564 28252 53732 28308
rect 53228 27022 53230 27074
rect 53282 27022 53284 27074
rect 52332 26852 52612 26908
rect 52668 26852 52948 26908
rect 53004 26964 53060 27002
rect 53228 26908 53284 27022
rect 53004 26898 53060 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 52332 26514 52388 26852
rect 52332 26462 52334 26514
rect 52386 26462 52388 26514
rect 52332 26450 52388 26462
rect 52556 26404 52612 26414
rect 52444 26402 52612 26404
rect 52444 26350 52558 26402
rect 52610 26350 52612 26402
rect 52444 26348 52612 26350
rect 52332 25620 52388 25630
rect 49084 25566 49086 25618
rect 49138 25566 49140 25618
rect 49084 25554 49140 25566
rect 49868 25618 50372 25620
rect 49868 25566 50318 25618
rect 50370 25566 50372 25618
rect 49868 25564 50372 25566
rect 49868 25508 49924 25564
rect 46956 25442 47012 25452
rect 49532 25506 49924 25508
rect 49532 25454 49870 25506
rect 49922 25454 49924 25506
rect 49532 25452 49924 25454
rect 45836 24946 45892 25340
rect 45836 24894 45838 24946
rect 45890 24894 45892 24946
rect 45836 24882 45892 24894
rect 49532 24722 49588 25452
rect 49868 25442 49924 25452
rect 50204 25284 50260 25294
rect 50204 24834 50260 25228
rect 50204 24782 50206 24834
rect 50258 24782 50260 24834
rect 50204 24770 50260 24782
rect 49532 24670 49534 24722
rect 49586 24670 49588 24722
rect 49532 24658 49588 24670
rect 45724 24546 45780 24556
rect 45164 23998 45166 24050
rect 45218 23998 45220 24050
rect 45164 23940 45220 23998
rect 45164 23874 45220 23884
rect 45500 24052 45556 24062
rect 45500 23938 45556 23996
rect 45500 23886 45502 23938
rect 45554 23886 45556 23938
rect 45500 23874 45556 23886
rect 46060 23940 46116 23950
rect 46060 23846 46116 23884
rect 45836 23714 45892 23726
rect 45836 23662 45838 23714
rect 45890 23662 45892 23714
rect 44604 23326 44606 23378
rect 44658 23326 44660 23378
rect 44604 23314 44660 23326
rect 45052 23380 45108 23390
rect 44940 23268 44996 23278
rect 44940 23174 44996 23212
rect 45052 23156 45108 23324
rect 45836 23380 45892 23662
rect 45836 23314 45892 23324
rect 46508 23714 46564 23726
rect 46508 23662 46510 23714
rect 46562 23662 46564 23714
rect 45612 23268 45668 23278
rect 45276 23156 45332 23166
rect 45052 23154 45556 23156
rect 45052 23102 45278 23154
rect 45330 23102 45556 23154
rect 45052 23100 45556 23102
rect 45052 22482 45108 23100
rect 45276 23090 45332 23100
rect 45052 22430 45054 22482
rect 45106 22430 45108 22482
rect 45052 22418 45108 22430
rect 45500 22482 45556 23100
rect 45500 22430 45502 22482
rect 45554 22430 45556 22482
rect 45500 22418 45556 22430
rect 45612 22372 45668 23212
rect 46060 23044 46116 23054
rect 45836 23042 46116 23044
rect 45836 22990 46062 23042
rect 46114 22990 46116 23042
rect 45836 22988 46116 22990
rect 45836 22482 45892 22988
rect 46060 22978 46116 22988
rect 46508 23044 46564 23662
rect 46508 22978 46564 22988
rect 46620 23714 46676 23726
rect 46620 23662 46622 23714
rect 46674 23662 46676 23714
rect 45836 22430 45838 22482
rect 45890 22430 45892 22482
rect 45836 22418 45892 22430
rect 46172 22708 46228 22718
rect 45388 22260 45444 22270
rect 45388 21476 45444 22204
rect 45276 21474 45444 21476
rect 45276 21422 45390 21474
rect 45442 21422 45444 21474
rect 45276 21420 45444 21422
rect 44716 19906 44772 19918
rect 44716 19854 44718 19906
rect 44770 19854 44772 19906
rect 44716 19012 44772 19854
rect 45164 19908 45220 19918
rect 45276 19908 45332 21420
rect 45388 21410 45444 21420
rect 45220 19852 45332 19908
rect 45164 19842 45220 19852
rect 45612 19234 45668 22316
rect 45948 22370 46004 22382
rect 45948 22318 45950 22370
rect 46002 22318 46004 22370
rect 45948 22260 46004 22318
rect 45948 22194 46004 22204
rect 46172 21924 46228 22652
rect 46284 22372 46340 22382
rect 46620 22372 46676 23662
rect 46732 23716 46788 23726
rect 46732 23714 46900 23716
rect 46732 23662 46734 23714
rect 46786 23662 46900 23714
rect 46732 23660 46900 23662
rect 46732 23650 46788 23660
rect 46844 23380 46900 23660
rect 50316 23604 50372 25564
rect 52220 25564 52332 25620
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 51436 23716 51492 23726
rect 50316 23548 50484 23604
rect 46284 22370 46676 22372
rect 46284 22318 46286 22370
rect 46338 22318 46676 22370
rect 46284 22316 46676 22318
rect 46732 22372 46788 22382
rect 46284 22306 46340 22316
rect 46172 21868 46452 21924
rect 46396 21810 46452 21868
rect 46396 21758 46398 21810
rect 46450 21758 46452 21810
rect 46284 20020 46340 20030
rect 46284 19906 46340 19964
rect 46284 19854 46286 19906
rect 46338 19854 46340 19906
rect 45612 19182 45614 19234
rect 45666 19182 45668 19234
rect 45612 19170 45668 19182
rect 46172 19460 46228 19470
rect 46172 19234 46228 19404
rect 46172 19182 46174 19234
rect 46226 19182 46228 19234
rect 46172 19170 46228 19182
rect 45948 19122 46004 19134
rect 45948 19070 45950 19122
rect 46002 19070 46004 19122
rect 44716 18564 44772 18956
rect 45276 19010 45332 19022
rect 45276 18958 45278 19010
rect 45330 18958 45332 19010
rect 45276 18676 45332 18958
rect 45276 18610 45332 18620
rect 45836 19010 45892 19022
rect 45836 18958 45838 19010
rect 45890 18958 45892 19010
rect 44716 18498 44772 18508
rect 45836 18562 45892 18958
rect 45948 18676 46004 19070
rect 45948 18610 46004 18620
rect 45836 18510 45838 18562
rect 45890 18510 45892 18562
rect 45836 18498 45892 18510
rect 45052 18452 45108 18462
rect 44492 18358 44548 18396
rect 44940 18450 45108 18452
rect 44940 18398 45054 18450
rect 45106 18398 45108 18450
rect 44940 18396 45108 18398
rect 44940 17668 44996 18396
rect 45052 18386 45108 18396
rect 44940 17574 44996 17612
rect 45276 17892 45332 17902
rect 43708 15092 43876 15148
rect 44268 15092 44436 15148
rect 44492 17444 44548 17454
rect 43708 14644 43764 15092
rect 43708 14642 44212 14644
rect 43708 14590 43710 14642
rect 43762 14590 44212 14642
rect 43708 14588 44212 14590
rect 43708 14578 43764 14588
rect 43708 13636 43764 13646
rect 43708 13542 43764 13580
rect 42364 13074 42924 13076
rect 42364 13022 42814 13074
rect 42866 13022 42924 13074
rect 42364 13020 42924 13022
rect 42364 12962 42420 13020
rect 42812 13010 42868 13020
rect 42924 12982 42980 13020
rect 43036 13074 43764 13076
rect 43036 13022 43374 13074
rect 43426 13022 43764 13074
rect 43036 13020 43764 13022
rect 42364 12910 42366 12962
rect 42418 12910 42420 12962
rect 42364 12898 42420 12910
rect 42588 12852 42644 12862
rect 43036 12852 43092 13020
rect 43372 13010 43428 13020
rect 43708 12962 43764 13020
rect 43708 12910 43710 12962
rect 43762 12910 43764 12962
rect 43708 12898 43764 12910
rect 42252 12460 42532 12516
rect 42028 12236 42196 12292
rect 42364 12292 42420 12302
rect 41244 12014 41246 12066
rect 41298 12014 41300 12066
rect 41244 12002 41300 12014
rect 41692 12066 41748 12078
rect 41692 12014 41694 12066
rect 41746 12014 41748 12066
rect 41692 11956 41748 12014
rect 41692 11890 41748 11900
rect 41020 11442 41076 11452
rect 42028 11396 42084 12236
rect 42028 11330 42084 11340
rect 42140 12068 42196 12078
rect 41692 10836 41748 10846
rect 41692 10742 41748 10780
rect 42140 10836 42196 12012
rect 42364 11506 42420 12236
rect 42364 11454 42366 11506
rect 42418 11454 42420 11506
rect 42364 11442 42420 11454
rect 42140 10770 42196 10780
rect 42252 11172 42308 11182
rect 42252 10612 42308 11116
rect 42252 10518 42308 10556
rect 42476 9940 42532 12460
rect 42588 12402 42644 12796
rect 42588 12350 42590 12402
rect 42642 12350 42644 12402
rect 42588 12338 42644 12350
rect 42700 12796 43092 12852
rect 42588 9940 42644 9950
rect 42476 9938 42644 9940
rect 42476 9886 42590 9938
rect 42642 9886 42644 9938
rect 42476 9884 42644 9886
rect 40572 9202 40628 9212
rect 41468 9826 41524 9838
rect 41468 9774 41470 9826
rect 41522 9774 41524 9826
rect 41468 8428 41524 9774
rect 42476 9380 42532 9884
rect 42588 9828 42644 9884
rect 42588 9762 42644 9772
rect 41916 9324 42532 9380
rect 41916 9266 41972 9324
rect 41916 9214 41918 9266
rect 41970 9214 41972 9266
rect 41916 9202 41972 9214
rect 42476 9266 42532 9324
rect 42476 9214 42478 9266
rect 42530 9214 42532 9266
rect 42476 9202 42532 9214
rect 42140 9154 42196 9166
rect 42140 9102 42142 9154
rect 42194 9102 42196 9154
rect 41468 8372 41972 8428
rect 40460 8194 40516 8204
rect 40012 8082 40068 8092
rect 41916 8036 41972 8372
rect 41916 7970 41972 7980
rect 39900 7858 39956 7868
rect 40796 7924 40852 7934
rect 40012 7700 40068 7710
rect 40012 7606 40068 7644
rect 39788 7534 39790 7586
rect 39842 7534 39844 7586
rect 39788 7522 39844 7534
rect 40124 7588 40180 7598
rect 40124 7494 40180 7532
rect 40348 7474 40404 7486
rect 40348 7422 40350 7474
rect 40402 7422 40404 7474
rect 40348 6804 40404 7422
rect 40684 7476 40740 7486
rect 40684 6916 40740 7420
rect 40796 7474 40852 7868
rect 41244 7868 41860 7924
rect 41244 7698 41300 7868
rect 41244 7646 41246 7698
rect 41298 7646 41300 7698
rect 41244 7634 41300 7646
rect 41468 7700 41524 7710
rect 40796 7422 40798 7474
rect 40850 7422 40852 7474
rect 40796 7410 40852 7422
rect 41356 7362 41412 7374
rect 41356 7310 41358 7362
rect 41410 7310 41412 7362
rect 41356 7028 41412 7310
rect 40908 6972 41412 7028
rect 40796 6916 40852 6926
rect 40684 6914 40852 6916
rect 40684 6862 40798 6914
rect 40850 6862 40852 6914
rect 40684 6860 40852 6862
rect 40124 6748 40404 6804
rect 40124 6692 40180 6748
rect 40012 6636 40180 6692
rect 40460 6692 40516 6702
rect 40796 6692 40852 6860
rect 40908 6914 40964 6972
rect 40908 6862 40910 6914
rect 40962 6862 40964 6914
rect 40908 6850 40964 6862
rect 41468 6916 41524 7644
rect 41580 7588 41636 7598
rect 41636 7532 41748 7588
rect 41580 7522 41636 7532
rect 41580 6916 41636 6926
rect 41468 6914 41636 6916
rect 41468 6862 41582 6914
rect 41634 6862 41636 6914
rect 41468 6860 41636 6862
rect 41580 6850 41636 6860
rect 41244 6692 41300 6702
rect 40796 6690 41300 6692
rect 40796 6638 41246 6690
rect 41298 6638 41300 6690
rect 40796 6636 41300 6638
rect 40012 6578 40068 6636
rect 40012 6526 40014 6578
rect 40066 6526 40068 6578
rect 40012 6132 40068 6526
rect 40236 6580 40292 6590
rect 40236 6486 40292 6524
rect 40460 6578 40516 6636
rect 41244 6626 41300 6636
rect 40460 6526 40462 6578
rect 40514 6526 40516 6578
rect 40460 6514 40516 6526
rect 40012 6066 40068 6076
rect 40124 6466 40180 6478
rect 40124 6414 40126 6466
rect 40178 6414 40180 6466
rect 40124 5796 40180 6414
rect 40124 5740 40740 5796
rect 39620 5292 39844 5348
rect 39564 5254 39620 5292
rect 39788 5236 39844 5292
rect 40348 5236 40404 5246
rect 39788 5180 40348 5236
rect 38220 5124 38276 5134
rect 38220 4562 38276 5068
rect 39116 5124 39172 5134
rect 39116 5030 39172 5068
rect 39788 5122 39844 5180
rect 40348 5142 40404 5180
rect 40684 5234 40740 5740
rect 41244 5794 41300 5806
rect 41244 5742 41246 5794
rect 41298 5742 41300 5794
rect 40684 5182 40686 5234
rect 40738 5182 40740 5234
rect 40684 5170 40740 5182
rect 40908 5236 40964 5246
rect 39788 5070 39790 5122
rect 39842 5070 39844 5122
rect 39788 5058 39844 5070
rect 38220 4510 38222 4562
rect 38274 4510 38276 4562
rect 38220 4498 38276 4510
rect 40796 4898 40852 4910
rect 40796 4846 40798 4898
rect 40850 4846 40852 4898
rect 38108 4398 38110 4450
rect 38162 4398 38164 4450
rect 38108 4386 38164 4398
rect 40796 4452 40852 4846
rect 40796 4386 40852 4396
rect 37212 4286 37214 4338
rect 37266 4286 37268 4338
rect 37212 4274 37268 4286
rect 40908 4338 40964 5180
rect 41244 5236 41300 5742
rect 41580 5796 41636 5806
rect 41692 5796 41748 7532
rect 41804 6692 41860 7868
rect 42140 7812 42196 9102
rect 42140 7746 42196 7756
rect 42588 7364 42644 7374
rect 42700 7364 42756 12796
rect 43036 11508 43092 11518
rect 42812 11452 43036 11508
rect 42812 10834 42868 11452
rect 42812 10782 42814 10834
rect 42866 10782 42868 10834
rect 42812 10770 42868 10782
rect 42924 10724 42980 10734
rect 42924 10164 42980 10668
rect 43036 10612 43092 11452
rect 43148 10612 43204 10622
rect 43036 10556 43148 10612
rect 43148 10518 43204 10556
rect 43820 10164 43876 14588
rect 44044 14420 44100 14430
rect 44044 13858 44100 14364
rect 44156 13970 44212 14588
rect 44156 13918 44158 13970
rect 44210 13918 44212 13970
rect 44156 13906 44212 13918
rect 44044 13806 44046 13858
rect 44098 13806 44100 13858
rect 44044 13794 44100 13806
rect 44156 13748 44212 13758
rect 44044 12852 44100 12862
rect 44044 12758 44100 12796
rect 43932 10724 43988 10734
rect 43932 10630 43988 10668
rect 42924 9826 42980 10108
rect 43708 10108 43876 10164
rect 43484 9940 43540 9950
rect 43708 9940 43764 10108
rect 43540 9884 43764 9940
rect 43484 9846 43540 9884
rect 42924 9774 42926 9826
rect 42978 9774 42980 9826
rect 42924 9762 42980 9774
rect 43820 9828 43876 9838
rect 43820 9734 43876 9772
rect 44156 9602 44212 13692
rect 44156 9550 44158 9602
rect 44210 9550 44212 9602
rect 42812 9268 42868 9278
rect 42812 9174 42868 9212
rect 43484 9268 43540 9278
rect 43484 9174 43540 9212
rect 43148 9154 43204 9166
rect 43148 9102 43150 9154
rect 43202 9102 43204 9154
rect 43148 8428 43204 9102
rect 43820 9154 43876 9166
rect 43820 9102 43822 9154
rect 43874 9102 43876 9154
rect 43820 8428 43876 9102
rect 43036 8372 43204 8428
rect 43708 8372 43876 8428
rect 42924 7474 42980 7486
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42924 7364 42980 7422
rect 42588 7362 42980 7364
rect 42588 7310 42590 7362
rect 42642 7310 42980 7362
rect 42588 7308 42980 7310
rect 42588 7252 42644 7308
rect 42588 7186 42644 7196
rect 41804 6598 41860 6636
rect 42924 6580 42980 6590
rect 43036 6580 43092 8372
rect 43596 7700 43652 7710
rect 43708 7700 43764 8372
rect 43596 7698 43708 7700
rect 43596 7646 43598 7698
rect 43650 7646 43708 7698
rect 43596 7644 43708 7646
rect 43596 7634 43652 7644
rect 43708 7606 43764 7644
rect 43260 7588 43316 7598
rect 43260 6804 43316 7532
rect 43820 7476 43876 7486
rect 43820 7382 43876 7420
rect 44156 7474 44212 9550
rect 44156 7422 44158 7474
rect 44210 7422 44212 7474
rect 43708 7362 43764 7374
rect 43708 7310 43710 7362
rect 43762 7310 43764 7362
rect 43708 6916 43764 7310
rect 44156 7362 44212 7422
rect 44156 7310 44158 7362
rect 44210 7310 44212 7362
rect 44156 7298 44212 7310
rect 43260 6738 43316 6748
rect 43484 6860 43764 6916
rect 43484 6690 43540 6860
rect 43484 6638 43486 6690
rect 43538 6638 43540 6690
rect 43484 6626 43540 6638
rect 43932 6692 43988 6702
rect 44268 6692 44324 15092
rect 44492 13972 44548 17388
rect 45052 15876 45108 15886
rect 45052 15426 45108 15820
rect 45052 15374 45054 15426
rect 45106 15374 45108 15426
rect 45052 15362 45108 15374
rect 45276 15314 45332 17836
rect 45388 15876 45444 15886
rect 45388 15782 45444 15820
rect 45724 15876 45780 15886
rect 45724 15782 45780 15820
rect 45276 15262 45278 15314
rect 45330 15262 45332 15314
rect 45276 15250 45332 15262
rect 45612 15316 45668 15326
rect 45724 15316 45780 15326
rect 45612 15314 45724 15316
rect 45612 15262 45614 15314
rect 45666 15262 45724 15314
rect 45612 15260 45724 15262
rect 44716 15204 44772 15242
rect 44716 15138 44772 15148
rect 45164 15202 45220 15214
rect 45164 15150 45166 15202
rect 45218 15150 45220 15202
rect 45052 14532 45108 14542
rect 45164 14532 45220 15150
rect 45052 14530 45220 14532
rect 45052 14478 45054 14530
rect 45106 14478 45220 14530
rect 45052 14476 45220 14478
rect 45052 14466 45108 14476
rect 44716 14420 44772 14430
rect 44716 14326 44772 14364
rect 44492 13906 44548 13916
rect 44940 14306 44996 14318
rect 44940 14254 44942 14306
rect 44994 14254 44996 14306
rect 44940 13860 44996 14254
rect 44940 13794 44996 13804
rect 45164 13858 45220 14476
rect 45164 13806 45166 13858
rect 45218 13806 45220 13858
rect 45164 13794 45220 13806
rect 44380 13748 44436 13758
rect 44380 13746 44884 13748
rect 44380 13694 44382 13746
rect 44434 13694 44884 13746
rect 44380 13692 44884 13694
rect 44380 13682 44436 13692
rect 44828 13186 44884 13692
rect 44828 13134 44830 13186
rect 44882 13134 44884 13186
rect 44828 13122 44884 13134
rect 44940 13634 44996 13646
rect 44940 13582 44942 13634
rect 44994 13582 44996 13634
rect 44940 13186 44996 13582
rect 44940 13134 44942 13186
rect 44994 13134 44996 13186
rect 44940 13122 44996 13134
rect 45612 12964 45668 15260
rect 45724 15250 45780 15260
rect 45836 12964 45892 12974
rect 45612 12962 46116 12964
rect 45612 12910 45838 12962
rect 45890 12910 46116 12962
rect 45612 12908 46116 12910
rect 45836 12898 45892 12908
rect 45276 12852 45332 12862
rect 45276 12758 45332 12796
rect 45500 12850 45556 12862
rect 45500 12798 45502 12850
rect 45554 12798 45556 12850
rect 44716 12740 44772 12750
rect 44716 12290 44772 12684
rect 45500 12628 45556 12798
rect 45612 12740 45668 12750
rect 45612 12646 45668 12684
rect 45500 12562 45556 12572
rect 44716 12238 44718 12290
rect 44770 12238 44772 12290
rect 44716 12226 44772 12238
rect 44604 11954 44660 11966
rect 44604 11902 44606 11954
rect 44658 11902 44660 11954
rect 44604 10724 44660 11902
rect 44604 10658 44660 10668
rect 43932 6690 44324 6692
rect 43932 6638 43934 6690
rect 43986 6638 44324 6690
rect 43932 6636 44324 6638
rect 44380 10612 44436 10622
rect 44380 9268 44436 10556
rect 46060 10498 46116 12908
rect 46060 10446 46062 10498
rect 46114 10446 46116 10498
rect 46060 10434 46116 10446
rect 44380 9266 44772 9268
rect 44380 9214 44382 9266
rect 44434 9214 44772 9266
rect 44380 9212 44772 9214
rect 42980 6524 43092 6580
rect 43260 6578 43316 6590
rect 43260 6526 43262 6578
rect 43314 6526 43316 6578
rect 42924 6486 42980 6524
rect 43148 6466 43204 6478
rect 43148 6414 43150 6466
rect 43202 6414 43204 6466
rect 43148 6244 43204 6414
rect 43260 6468 43316 6526
rect 43260 6402 43316 6412
rect 43932 6468 43988 6636
rect 43932 6402 43988 6412
rect 43148 6188 43540 6244
rect 43484 6132 43540 6188
rect 43820 6132 43876 6142
rect 43484 6076 43764 6132
rect 43708 6018 43764 6076
rect 43708 5966 43710 6018
rect 43762 5966 43764 6018
rect 43708 5954 43764 5966
rect 41580 5794 41748 5796
rect 41580 5742 41582 5794
rect 41634 5742 41748 5794
rect 41580 5740 41748 5742
rect 41580 5730 41636 5740
rect 41244 5170 41300 5180
rect 41692 4452 41748 4462
rect 41692 4358 41748 4396
rect 40908 4286 40910 4338
rect 40962 4286 40964 4338
rect 40908 4274 40964 4286
rect 34300 4226 35140 4228
rect 34300 4174 34302 4226
rect 34354 4174 35140 4226
rect 34300 4172 35140 4174
rect 43820 4226 43876 6076
rect 44380 5908 44436 9212
rect 44716 9042 44772 9212
rect 44716 8990 44718 9042
rect 44770 8990 44772 9042
rect 44716 8978 44772 8990
rect 45500 8930 45556 8942
rect 45500 8878 45502 8930
rect 45554 8878 45556 8930
rect 44940 8260 44996 8270
rect 45164 8260 45220 8270
rect 44940 8166 44996 8204
rect 45052 8258 45220 8260
rect 45052 8206 45166 8258
rect 45218 8206 45220 8258
rect 45052 8204 45220 8206
rect 44044 5906 44436 5908
rect 44044 5854 44382 5906
rect 44434 5854 44436 5906
rect 44044 5852 44436 5854
rect 44044 5234 44100 5852
rect 44380 5842 44436 5852
rect 44604 7362 44660 7374
rect 44604 7310 44606 7362
rect 44658 7310 44660 7362
rect 44604 7250 44660 7310
rect 44604 7198 44606 7250
rect 44658 7198 44660 7250
rect 44044 5182 44046 5234
rect 44098 5182 44100 5234
rect 44044 4340 44100 5182
rect 44604 5124 44660 7198
rect 45052 6580 45108 8204
rect 45164 8194 45220 8204
rect 45500 8034 45556 8878
rect 46284 8428 46340 19854
rect 46396 15540 46452 21758
rect 46620 20132 46676 20142
rect 46732 20132 46788 22316
rect 46844 21588 46900 23324
rect 47964 23156 48020 23166
rect 47180 22708 47236 22718
rect 47068 22258 47124 22270
rect 47068 22206 47070 22258
rect 47122 22206 47124 22258
rect 46956 22146 47012 22158
rect 46956 22094 46958 22146
rect 47010 22094 47012 22146
rect 46956 21812 47012 22094
rect 46956 21746 47012 21756
rect 47068 21810 47124 22206
rect 47180 22258 47236 22652
rect 47180 22206 47182 22258
rect 47234 22206 47236 22258
rect 47180 22194 47236 22206
rect 47516 22482 47572 22494
rect 47516 22430 47518 22482
rect 47570 22430 47572 22482
rect 47516 22148 47572 22430
rect 47964 22370 48020 23100
rect 50428 23156 50484 23548
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 51436 23266 51492 23660
rect 52220 23492 52276 25564
rect 52332 25554 52388 25564
rect 52444 25396 52500 26348
rect 52556 26338 52612 26348
rect 52668 26402 52724 26852
rect 52668 26350 52670 26402
rect 52722 26350 52724 26402
rect 52668 26338 52724 26350
rect 52332 24612 52388 24622
rect 52444 24612 52500 25340
rect 52556 25506 52612 25518
rect 52556 25454 52558 25506
rect 52610 25454 52612 25506
rect 52556 24946 52612 25454
rect 52780 25284 52836 25294
rect 52780 25190 52836 25228
rect 52556 24894 52558 24946
rect 52610 24894 52612 24946
rect 52556 24882 52612 24894
rect 52780 24836 52836 24846
rect 52332 24610 52500 24612
rect 52332 24558 52334 24610
rect 52386 24558 52500 24610
rect 52332 24556 52500 24558
rect 52668 24834 52836 24836
rect 52668 24782 52782 24834
rect 52834 24782 52836 24834
rect 52668 24780 52836 24782
rect 52332 24546 52388 24556
rect 52668 23828 52724 24780
rect 52780 24770 52836 24780
rect 52892 24836 52948 26852
rect 53116 26852 53284 26908
rect 53452 26964 53508 27002
rect 53452 26898 53508 26908
rect 53116 25732 53172 26852
rect 53116 25676 53396 25732
rect 53004 25508 53060 25518
rect 53004 25414 53060 25452
rect 53116 25508 53172 25518
rect 53340 25508 53396 25676
rect 53564 25620 53620 28252
rect 53676 27860 53732 27870
rect 53676 27076 53732 27804
rect 54236 27748 54292 27758
rect 53788 27076 53844 27086
rect 53676 27074 53844 27076
rect 53676 27022 53790 27074
rect 53842 27022 53844 27074
rect 53676 27020 53844 27022
rect 53676 26852 53732 26862
rect 53676 26758 53732 26796
rect 53564 25554 53620 25564
rect 53116 25506 53396 25508
rect 53116 25454 53118 25506
rect 53170 25454 53396 25506
rect 53116 25452 53396 25454
rect 53452 25508 53508 25518
rect 52892 24770 52948 24780
rect 53116 24612 53172 25452
rect 53452 25414 53508 25452
rect 53788 25506 53844 27020
rect 54236 26964 54292 27692
rect 54460 27076 54516 28588
rect 55132 28532 55188 30380
rect 55244 30212 55300 31726
rect 55356 31106 55412 31118
rect 55356 31054 55358 31106
rect 55410 31054 55412 31106
rect 55356 30996 55412 31054
rect 55356 30930 55412 30940
rect 55356 30212 55412 30222
rect 55244 30210 55412 30212
rect 55244 30158 55358 30210
rect 55410 30158 55412 30210
rect 55244 30156 55412 30158
rect 55132 28466 55188 28476
rect 55356 28756 55412 30156
rect 54684 28084 54740 28094
rect 55356 28084 55412 28700
rect 54684 28082 55412 28084
rect 54684 28030 54686 28082
rect 54738 28030 55412 28082
rect 54684 28028 55412 28030
rect 54684 28018 54740 28028
rect 55132 27860 55188 27870
rect 55132 27766 55188 27804
rect 54460 27010 54516 27020
rect 55356 27074 55412 28028
rect 55468 27972 55524 27982
rect 55468 27878 55524 27916
rect 55356 27022 55358 27074
rect 55410 27022 55412 27074
rect 55356 27010 55412 27022
rect 54236 26898 54292 26908
rect 53788 25454 53790 25506
rect 53842 25454 53844 25506
rect 53564 25396 53620 25406
rect 53620 25340 53732 25396
rect 53564 25330 53620 25340
rect 53676 25282 53732 25340
rect 53676 25230 53678 25282
rect 53730 25230 53732 25282
rect 53676 25218 53732 25230
rect 53340 25004 53620 25060
rect 53340 24890 53396 25004
rect 53340 24838 53342 24890
rect 53394 24838 53396 24890
rect 53340 24826 53396 24838
rect 53452 24834 53508 24846
rect 53452 24782 53454 24834
rect 53506 24782 53508 24834
rect 53340 24724 53396 24734
rect 53452 24724 53508 24782
rect 53396 24668 53508 24724
rect 53340 24658 53396 24668
rect 52780 24556 53172 24612
rect 52780 23938 52836 24556
rect 53340 24498 53396 24510
rect 53340 24446 53342 24498
rect 53394 24446 53396 24498
rect 52780 23886 52782 23938
rect 52834 23886 52836 23938
rect 52780 23874 52836 23886
rect 53004 23940 53060 23950
rect 53004 23938 53172 23940
rect 53004 23886 53006 23938
rect 53058 23886 53172 23938
rect 53004 23884 53172 23886
rect 53004 23874 53060 23884
rect 52668 23762 52724 23772
rect 53004 23716 53060 23726
rect 53116 23716 53172 23884
rect 53340 23938 53396 24446
rect 53340 23886 53342 23938
rect 53394 23886 53396 23938
rect 53340 23874 53396 23886
rect 53452 23716 53508 23726
rect 53116 23714 53508 23716
rect 53116 23662 53454 23714
rect 53506 23662 53508 23714
rect 53116 23660 53508 23662
rect 53004 23622 53060 23660
rect 53452 23650 53508 23660
rect 52220 23436 52612 23492
rect 51436 23214 51438 23266
rect 51490 23214 51492 23266
rect 51436 23202 51492 23214
rect 52220 23268 52276 23278
rect 50428 23090 50484 23100
rect 50764 23154 50820 23166
rect 50764 23102 50766 23154
rect 50818 23102 50820 23154
rect 48188 23044 48244 23054
rect 48188 22484 48244 22988
rect 50764 23044 50820 23102
rect 50764 22978 50820 22988
rect 51212 23044 51268 23054
rect 48188 22418 48244 22428
rect 50204 22484 50260 22494
rect 47964 22318 47966 22370
rect 48018 22318 48020 22370
rect 47964 22306 48020 22318
rect 48636 22260 48692 22270
rect 48076 22258 48692 22260
rect 48076 22206 48638 22258
rect 48690 22206 48692 22258
rect 48076 22204 48692 22206
rect 48076 22148 48132 22204
rect 48636 22194 48692 22204
rect 47516 22092 48132 22148
rect 47068 21758 47070 21810
rect 47122 21758 47124 21810
rect 47068 21746 47124 21758
rect 47292 21812 47348 21822
rect 49644 21812 49700 21822
rect 47292 21810 47908 21812
rect 47292 21758 47294 21810
rect 47346 21758 47908 21810
rect 47292 21756 47908 21758
rect 47292 21746 47348 21756
rect 47404 21588 47460 21598
rect 46844 21586 47572 21588
rect 46844 21534 47406 21586
rect 47458 21534 47572 21586
rect 46844 21532 47572 21534
rect 47404 21522 47460 21532
rect 46620 20130 46788 20132
rect 46620 20078 46622 20130
rect 46674 20078 46788 20130
rect 46620 20076 46788 20078
rect 47292 20578 47348 20590
rect 47292 20526 47294 20578
rect 47346 20526 47348 20578
rect 46620 20066 46676 20076
rect 46844 20020 46900 20030
rect 46844 19926 46900 19964
rect 47068 20018 47124 20030
rect 47068 19966 47070 20018
rect 47122 19966 47124 20018
rect 46732 19908 46788 19918
rect 46732 19814 46788 19852
rect 46956 19796 47012 19806
rect 46732 18564 46788 18574
rect 46620 17444 46676 17454
rect 46620 17350 46676 17388
rect 46396 15484 46564 15540
rect 45612 8372 46340 8428
rect 45612 8260 45668 8372
rect 45612 8166 45668 8204
rect 45836 8260 45892 8270
rect 46284 8260 46340 8270
rect 45836 8258 46340 8260
rect 45836 8206 45838 8258
rect 45890 8206 46286 8258
rect 46338 8206 46340 8258
rect 45836 8204 46340 8206
rect 45836 8194 45892 8204
rect 46284 8194 46340 8204
rect 46396 8260 46452 8270
rect 46396 8166 46452 8204
rect 45500 7982 45502 8034
rect 45554 7982 45556 8034
rect 45500 7970 45556 7982
rect 46172 8034 46228 8046
rect 46172 7982 46174 8034
rect 46226 7982 46228 8034
rect 45836 7812 45892 7822
rect 45836 7698 45892 7756
rect 45836 7646 45838 7698
rect 45890 7646 45892 7698
rect 45836 7634 45892 7646
rect 46172 7700 46228 7982
rect 45052 5908 45108 6524
rect 46172 6020 46228 7644
rect 46396 6804 46452 6814
rect 46508 6804 46564 15484
rect 46620 15204 46676 15242
rect 46620 15138 46676 15148
rect 46732 15092 46788 18508
rect 46956 17666 47012 19740
rect 47068 17778 47124 19966
rect 47292 20020 47348 20526
rect 47180 19236 47236 19246
rect 47180 19142 47236 19180
rect 47068 17726 47070 17778
rect 47122 17726 47124 17778
rect 47068 17714 47124 17726
rect 46956 17614 46958 17666
rect 47010 17614 47012 17666
rect 46956 17602 47012 17614
rect 47180 17668 47236 17678
rect 47180 17574 47236 17612
rect 47292 17444 47348 19964
rect 47516 20018 47572 21532
rect 47852 21474 47908 21756
rect 49644 21718 49700 21756
rect 49756 21700 49812 21710
rect 49756 21606 49812 21644
rect 47852 21422 47854 21474
rect 47906 21422 47908 21474
rect 47852 20356 47908 21422
rect 47852 20300 48132 20356
rect 47964 20130 48020 20142
rect 47964 20078 47966 20130
rect 48018 20078 48020 20130
rect 47516 19966 47518 20018
rect 47570 19966 47572 20018
rect 47516 19796 47572 19966
rect 47740 20018 47796 20030
rect 47740 19966 47742 20018
rect 47794 19966 47796 20018
rect 47516 19730 47572 19740
rect 47628 19906 47684 19918
rect 47628 19854 47630 19906
rect 47682 19854 47684 19906
rect 47628 19460 47684 19854
rect 47628 19394 47684 19404
rect 47740 19348 47796 19966
rect 47964 20020 48020 20078
rect 47964 19954 48020 19964
rect 47740 18340 47796 19292
rect 47852 19908 47908 19918
rect 47852 19346 47908 19852
rect 47852 19294 47854 19346
rect 47906 19294 47908 19346
rect 47852 19282 47908 19294
rect 47964 18340 48020 18350
rect 47740 18338 48020 18340
rect 47740 18286 47966 18338
rect 48018 18286 48020 18338
rect 47740 18284 48020 18286
rect 47964 18274 48020 18284
rect 47404 17444 47460 17454
rect 47292 17388 47404 17444
rect 47404 17350 47460 17388
rect 47852 15988 47908 15998
rect 47852 15894 47908 15932
rect 47180 15876 47236 15886
rect 47180 15428 47236 15820
rect 47740 15876 47796 15886
rect 46844 15316 46900 15326
rect 46844 15222 46900 15260
rect 47068 15202 47124 15214
rect 47068 15150 47070 15202
rect 47122 15150 47124 15202
rect 47068 15148 47124 15150
rect 46956 15092 47124 15148
rect 46732 15036 46900 15092
rect 46732 14530 46788 14542
rect 46732 14478 46734 14530
rect 46786 14478 46788 14530
rect 46732 14308 46788 14478
rect 46844 14530 46900 15036
rect 46844 14478 46846 14530
rect 46898 14478 46900 14530
rect 46844 14466 46900 14478
rect 46956 14308 47012 15092
rect 47180 14418 47236 15372
rect 47292 15540 47348 15550
rect 47292 15314 47348 15484
rect 47740 15538 47796 15820
rect 47740 15486 47742 15538
rect 47794 15486 47796 15538
rect 47740 15474 47796 15486
rect 47292 15262 47294 15314
rect 47346 15262 47348 15314
rect 47292 15250 47348 15262
rect 48076 15148 48132 20300
rect 49980 19346 50036 19358
rect 49980 19294 49982 19346
rect 50034 19294 50036 19346
rect 49980 17668 50036 19294
rect 49980 17602 50036 17612
rect 48972 16994 49028 17006
rect 48972 16942 48974 16994
rect 49026 16942 49028 16994
rect 48972 15764 49028 16942
rect 49308 16884 49364 16894
rect 48860 15708 49028 15764
rect 49084 16772 49140 16782
rect 48860 15428 48916 15708
rect 48860 15362 48916 15372
rect 48972 15540 49028 15550
rect 48972 15314 49028 15484
rect 49084 15426 49140 16716
rect 49308 16210 49364 16828
rect 50204 16660 50260 22428
rect 50764 22484 50820 22494
rect 50764 22482 50932 22484
rect 50764 22430 50766 22482
rect 50818 22430 50932 22482
rect 50764 22428 50932 22430
rect 50764 22418 50820 22428
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50876 21700 50932 22428
rect 51212 22482 51268 22988
rect 51212 22430 51214 22482
rect 51266 22430 51268 22482
rect 51212 22418 51268 22430
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 19906 50372 19918
rect 50316 19854 50318 19906
rect 50370 19854 50372 19906
rect 50316 19236 50372 19854
rect 50316 19170 50372 19180
rect 50764 19348 50820 19358
rect 50764 19234 50820 19292
rect 50764 19182 50766 19234
rect 50818 19182 50820 19234
rect 50764 19170 50820 19182
rect 50540 19124 50596 19134
rect 50428 19122 50596 19124
rect 50428 19070 50542 19122
rect 50594 19070 50596 19122
rect 50428 19068 50596 19070
rect 50316 18788 50372 18798
rect 50316 18452 50372 18732
rect 50428 18676 50484 19068
rect 50540 19058 50596 19068
rect 50764 19012 50820 19050
rect 50764 18946 50820 18956
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50428 18610 50484 18620
rect 50876 18562 50932 21644
rect 52220 21474 52276 23212
rect 52220 21422 52222 21474
rect 52274 21422 52276 21474
rect 52220 21410 52276 21422
rect 51212 19908 51268 19918
rect 51212 19906 51940 19908
rect 51212 19854 51214 19906
rect 51266 19854 51940 19906
rect 51212 19852 51940 19854
rect 51212 19842 51268 19852
rect 50876 18510 50878 18562
rect 50930 18510 50932 18562
rect 50876 18498 50932 18510
rect 50988 19234 51044 19246
rect 50988 19182 50990 19234
rect 51042 19182 51044 19234
rect 50428 18452 50484 18462
rect 50316 18450 50484 18452
rect 50316 18398 50430 18450
rect 50482 18398 50484 18450
rect 50316 18396 50484 18398
rect 50316 17666 50372 18396
rect 50428 18386 50484 18396
rect 50988 18004 51044 19182
rect 51324 19180 51716 19236
rect 51324 18674 51380 19180
rect 51324 18622 51326 18674
rect 51378 18622 51380 18674
rect 51324 18610 51380 18622
rect 51436 19010 51492 19022
rect 51436 18958 51438 19010
rect 51490 18958 51492 19010
rect 51324 18450 51380 18462
rect 51324 18398 51326 18450
rect 51378 18398 51380 18450
rect 51324 18116 51380 18398
rect 51324 18050 51380 18060
rect 50876 17948 51044 18004
rect 50316 17614 50318 17666
rect 50370 17614 50372 17666
rect 50316 16884 50372 17614
rect 50652 17668 50708 17678
rect 50652 17574 50708 17612
rect 50876 17668 50932 17948
rect 51436 17892 51492 18958
rect 51548 19010 51604 19022
rect 51548 18958 51550 19010
rect 51602 18958 51604 19010
rect 51548 18452 51604 18958
rect 51548 18386 51604 18396
rect 51660 19010 51716 19180
rect 51884 19124 51940 19852
rect 51660 18958 51662 19010
rect 51714 18958 51716 19010
rect 51548 17892 51604 17902
rect 51324 17890 51604 17892
rect 51324 17838 51550 17890
rect 51602 17838 51604 17890
rect 51324 17836 51604 17838
rect 50876 17602 50932 17612
rect 50988 17780 51044 17790
rect 51324 17780 51380 17836
rect 51548 17826 51604 17836
rect 50988 17666 51044 17724
rect 50988 17614 50990 17666
rect 51042 17614 51044 17666
rect 50988 17602 51044 17614
rect 51100 17724 51380 17780
rect 50652 17444 50708 17454
rect 51100 17444 51156 17724
rect 51660 17668 51716 18958
rect 50652 17442 51156 17444
rect 50652 17390 50654 17442
rect 50706 17390 51156 17442
rect 50652 17388 51156 17390
rect 51324 17612 51716 17668
rect 51772 19122 51940 19124
rect 51772 19070 51886 19122
rect 51938 19070 51940 19122
rect 51772 19068 51940 19070
rect 51324 17610 51380 17612
rect 51324 17558 51326 17610
rect 51378 17558 51380 17610
rect 50652 17378 50708 17388
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50316 16818 50372 16828
rect 51212 17108 51268 17118
rect 50204 16604 50372 16660
rect 49308 16158 49310 16210
rect 49362 16158 49364 16210
rect 49308 16146 49364 16158
rect 49532 16098 49588 16110
rect 49532 16046 49534 16098
rect 49586 16046 49588 16098
rect 49084 15374 49086 15426
rect 49138 15374 49140 15426
rect 49084 15362 49140 15374
rect 49420 15428 49476 15438
rect 49420 15334 49476 15372
rect 48972 15262 48974 15314
rect 49026 15262 49028 15314
rect 48972 15250 49028 15262
rect 49308 15202 49364 15214
rect 49308 15150 49310 15202
rect 49362 15150 49364 15202
rect 48076 15092 48468 15148
rect 47852 14644 47908 14654
rect 47180 14366 47182 14418
rect 47234 14366 47236 14418
rect 47180 14354 47236 14366
rect 47404 14642 47908 14644
rect 47404 14590 47854 14642
rect 47906 14590 47908 14642
rect 47404 14588 47908 14590
rect 46732 14252 47012 14308
rect 47068 14306 47124 14318
rect 47068 14254 47070 14306
rect 47122 14254 47124 14306
rect 46732 12964 46788 14252
rect 47068 14196 47124 14254
rect 47404 14196 47460 14588
rect 47628 14420 47684 14430
rect 47068 14140 47460 14196
rect 47516 14306 47572 14318
rect 47516 14254 47518 14306
rect 47570 14254 47572 14306
rect 47404 13858 47460 13870
rect 47404 13806 47406 13858
rect 47458 13806 47460 13858
rect 47404 13748 47460 13806
rect 47292 13692 47404 13748
rect 47180 12964 47236 12974
rect 46732 12962 47236 12964
rect 46732 12910 47182 12962
rect 47234 12910 47236 12962
rect 46732 12908 47236 12910
rect 46732 11506 46788 12908
rect 47180 12898 47236 12908
rect 46732 11454 46734 11506
rect 46786 11454 46788 11506
rect 46732 11442 46788 11454
rect 46956 11620 47012 11630
rect 46956 10948 47012 11564
rect 46844 10610 46900 10622
rect 46844 10558 46846 10610
rect 46898 10558 46900 10610
rect 46844 10164 46900 10558
rect 46844 10098 46900 10108
rect 46956 8428 47012 10892
rect 47180 10836 47236 10846
rect 47292 10836 47348 13692
rect 47404 13682 47460 13692
rect 47516 13860 47572 14254
rect 47628 13970 47684 14364
rect 47628 13918 47630 13970
rect 47682 13918 47684 13970
rect 47628 13906 47684 13918
rect 47852 13970 47908 14588
rect 48076 14532 48132 14542
rect 48076 14438 48132 14476
rect 47852 13918 47854 13970
rect 47906 13918 47908 13970
rect 47852 13906 47908 13918
rect 48300 14420 48356 14430
rect 47516 13076 47572 13804
rect 47740 13634 47796 13646
rect 47740 13582 47742 13634
rect 47794 13582 47796 13634
rect 47740 13300 47796 13582
rect 47740 13244 48244 13300
rect 48188 13186 48244 13244
rect 48188 13134 48190 13186
rect 48242 13134 48244 13186
rect 48188 13122 48244 13134
rect 48076 13076 48132 13086
rect 47516 13074 48132 13076
rect 47516 13022 48078 13074
rect 48130 13022 48132 13074
rect 47516 13020 48132 13022
rect 48076 13010 48132 13020
rect 48300 12964 48356 14364
rect 48188 12908 48356 12964
rect 47516 12850 47572 12862
rect 47516 12798 47518 12850
rect 47570 12798 47572 12850
rect 47404 12738 47460 12750
rect 47404 12686 47406 12738
rect 47458 12686 47460 12738
rect 47404 12404 47460 12686
rect 47516 12628 47572 12798
rect 47852 12852 47908 12862
rect 48188 12852 48244 12908
rect 47908 12796 48244 12852
rect 47852 12758 47908 12796
rect 47516 12562 47572 12572
rect 47404 12348 47796 12404
rect 47740 12290 47796 12348
rect 47740 12238 47742 12290
rect 47794 12238 47796 12290
rect 47740 12226 47796 12238
rect 47852 11954 47908 11966
rect 47852 11902 47854 11954
rect 47906 11902 47908 11954
rect 47852 11508 47908 11902
rect 48412 11620 48468 15092
rect 49308 14756 49364 15150
rect 49308 14690 49364 14700
rect 49532 12516 49588 16046
rect 49980 15428 50036 15438
rect 49980 15314 50036 15372
rect 49980 15262 49982 15314
rect 50034 15262 50036 15314
rect 49980 15250 50036 15262
rect 50316 15314 50372 16604
rect 50540 15988 50596 15998
rect 50540 15894 50596 15932
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50316 15262 50318 15314
rect 50370 15262 50372 15314
rect 50316 15250 50372 15262
rect 50652 15314 50708 15326
rect 50652 15262 50654 15314
rect 50706 15262 50708 15314
rect 50204 15204 50260 15242
rect 50204 15138 50260 15148
rect 50652 15092 50708 15262
rect 51100 15092 51156 15102
rect 50652 15026 50708 15036
rect 50988 15090 51156 15092
rect 50988 15038 51102 15090
rect 51154 15038 51156 15090
rect 50988 15036 51156 15038
rect 50540 14756 50596 14766
rect 50428 14644 50484 14654
rect 50204 14532 50260 14542
rect 50204 14438 50260 14476
rect 50428 13972 50484 14588
rect 50540 14308 50596 14700
rect 50764 14644 50820 14654
rect 50988 14644 51044 15036
rect 51100 15026 51156 15036
rect 51212 14868 51268 17052
rect 51212 14802 51268 14812
rect 50820 14588 51044 14644
rect 50764 14550 50820 14588
rect 51100 14532 51156 14542
rect 50540 14242 50596 14252
rect 50876 14530 51156 14532
rect 50876 14478 51102 14530
rect 51154 14478 51156 14530
rect 50876 14476 51156 14478
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50652 13972 50708 13982
rect 50428 13970 50708 13972
rect 50428 13918 50654 13970
rect 50706 13918 50708 13970
rect 50428 13916 50708 13918
rect 50652 13906 50708 13916
rect 50764 13972 50820 13982
rect 50876 13972 50932 14476
rect 51100 14466 51156 14476
rect 51212 14532 51268 14542
rect 51212 14438 51268 14476
rect 50764 13970 50932 13972
rect 50764 13918 50766 13970
rect 50818 13918 50932 13970
rect 50764 13916 50932 13918
rect 50988 14308 51044 14318
rect 51324 14308 51380 17558
rect 51660 17108 51716 17118
rect 51772 17108 51828 19068
rect 51884 19058 51940 19068
rect 52220 18452 52276 18462
rect 52220 18358 52276 18396
rect 52444 18340 52500 18350
rect 52332 18228 52388 18238
rect 51716 17052 51828 17108
rect 51884 18172 52332 18228
rect 51884 17890 51940 18172
rect 52332 18134 52388 18172
rect 51884 17838 51886 17890
rect 51938 17838 51940 17890
rect 51884 17106 51940 17838
rect 52108 17892 52164 17902
rect 51884 17054 51886 17106
rect 51938 17054 51940 17106
rect 51660 17014 51716 17052
rect 51884 17042 51940 17054
rect 51996 17108 52052 17118
rect 51660 16884 51716 16894
rect 51660 16098 51716 16828
rect 51996 16770 52052 17052
rect 52108 17106 52164 17836
rect 52108 17054 52110 17106
rect 52162 17054 52164 17106
rect 52108 17042 52164 17054
rect 52332 17892 52388 17902
rect 51996 16718 51998 16770
rect 52050 16718 52052 16770
rect 51996 16706 52052 16718
rect 52220 16772 52276 16782
rect 51660 16046 51662 16098
rect 51714 16046 51716 16098
rect 51660 16034 51716 16046
rect 52108 15874 52164 15886
rect 52108 15822 52110 15874
rect 52162 15822 52164 15874
rect 51660 15540 51716 15550
rect 52108 15540 52164 15822
rect 51660 15314 51716 15484
rect 51660 15262 51662 15314
rect 51714 15262 51716 15314
rect 51660 15250 51716 15262
rect 51884 15538 52164 15540
rect 51884 15486 52110 15538
rect 52162 15486 52164 15538
rect 51884 15484 52164 15486
rect 51436 15204 51492 15242
rect 51436 15138 51492 15148
rect 51884 14868 51940 15484
rect 52108 15474 52164 15484
rect 51884 14802 51940 14812
rect 52108 15316 52164 15326
rect 52108 14532 52164 15260
rect 52108 14438 52164 14476
rect 51772 14420 51828 14430
rect 51660 14364 51772 14420
rect 50764 13906 50820 13916
rect 50204 13748 50260 13758
rect 50204 13654 50260 13692
rect 50876 13748 50932 13758
rect 50988 13748 51044 14252
rect 50876 13746 51044 13748
rect 50876 13694 50878 13746
rect 50930 13694 51044 13746
rect 50876 13692 51044 13694
rect 51212 14252 51380 14308
rect 51548 14308 51604 14318
rect 50876 13682 50932 13692
rect 50316 13636 50372 13646
rect 49532 12450 49588 12460
rect 49756 13076 49812 13086
rect 49756 12404 49812 13020
rect 49756 12310 49812 12348
rect 50204 12628 50260 12638
rect 48412 11554 48468 11564
rect 49868 11620 49924 11630
rect 47852 11442 47908 11452
rect 48860 11508 48916 11518
rect 48860 11414 48916 11452
rect 49644 11508 49700 11518
rect 49644 11394 49700 11452
rect 49644 11342 49646 11394
rect 49698 11342 49700 11394
rect 49644 11330 49700 11342
rect 47180 10834 47348 10836
rect 47180 10782 47182 10834
rect 47234 10782 47348 10834
rect 47180 10780 47348 10782
rect 47180 10770 47236 10780
rect 47292 9268 47348 10780
rect 49868 10610 49924 11564
rect 50092 11508 50148 11518
rect 50092 11414 50148 11452
rect 49868 10558 49870 10610
rect 49922 10558 49924 10610
rect 49532 10500 49588 10510
rect 49868 10500 49924 10558
rect 49532 10498 49924 10500
rect 49532 10446 49534 10498
rect 49586 10446 49924 10498
rect 49532 10444 49924 10446
rect 50204 10722 50260 12572
rect 50316 12292 50372 13580
rect 51100 12738 51156 12750
rect 51100 12686 51102 12738
rect 51154 12686 51156 12738
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50316 12178 50372 12236
rect 50316 12126 50318 12178
rect 50370 12126 50372 12178
rect 50316 12114 50372 12126
rect 50652 12404 50708 12414
rect 50652 11506 50708 12348
rect 50988 12290 51044 12302
rect 50988 12238 50990 12290
rect 51042 12238 51044 12290
rect 50988 11956 51044 12238
rect 50988 11890 51044 11900
rect 51100 11620 51156 12686
rect 51100 11554 51156 11564
rect 50652 11454 50654 11506
rect 50706 11454 50708 11506
rect 50652 11442 50708 11454
rect 50988 11396 51044 11406
rect 51212 11396 51268 14252
rect 51548 14214 51604 14252
rect 51436 12738 51492 12750
rect 51436 12686 51438 12738
rect 51490 12686 51492 12738
rect 51436 12404 51492 12686
rect 51436 12338 51492 12348
rect 51660 12402 51716 14364
rect 51772 14326 51828 14364
rect 51884 14306 51940 14318
rect 51884 14254 51886 14306
rect 51938 14254 51940 14306
rect 51884 13748 51940 14254
rect 52220 14196 52276 16716
rect 52332 15540 52388 17836
rect 52444 17444 52500 18284
rect 52444 17378 52500 17388
rect 52556 16548 52612 23436
rect 53564 23268 53620 25004
rect 53788 23938 53844 25454
rect 53788 23886 53790 23938
rect 53842 23886 53844 23938
rect 53564 23202 53620 23212
rect 53676 23716 53732 23754
rect 53564 23044 53620 23054
rect 53676 23044 53732 23660
rect 53564 23042 53732 23044
rect 53564 22990 53566 23042
rect 53618 22990 53732 23042
rect 53564 22988 53732 22990
rect 53564 22978 53620 22988
rect 53788 22820 53844 23886
rect 53900 24610 53956 24622
rect 53900 24558 53902 24610
rect 53954 24558 53956 24610
rect 53900 23044 53956 24558
rect 55916 24500 55972 38612
rect 56700 38052 56756 38612
rect 57708 38500 57764 44942
rect 57820 43650 57876 59052
rect 58156 58548 58212 59164
rect 58268 58548 58324 58558
rect 58156 58546 58324 58548
rect 58156 58494 58270 58546
rect 58322 58494 58324 58546
rect 58156 58492 58324 58494
rect 58268 58482 58324 58492
rect 58156 55300 58212 55310
rect 58156 55206 58212 55244
rect 58156 54292 58212 54302
rect 58156 53842 58212 54236
rect 58156 53790 58158 53842
rect 58210 53790 58212 53842
rect 58156 53778 58212 53790
rect 58156 52946 58212 52958
rect 58156 52894 58158 52946
rect 58210 52894 58212 52946
rect 58156 52836 58212 52894
rect 58156 52276 58212 52780
rect 58156 52210 58212 52220
rect 58156 51604 58212 51614
rect 58156 50706 58212 51548
rect 58156 50654 58158 50706
rect 58210 50654 58212 50706
rect 58156 50642 58212 50654
rect 58156 49252 58212 49262
rect 58156 49138 58212 49196
rect 58156 49086 58158 49138
rect 58210 49086 58212 49138
rect 58156 49074 58212 49086
rect 58044 45892 58100 45902
rect 58044 45798 58100 45836
rect 58156 45332 58212 45342
rect 58212 45276 58324 45332
rect 58156 45238 58212 45276
rect 58268 44434 58324 45276
rect 58268 44382 58270 44434
rect 58322 44382 58324 44434
rect 58268 44370 58324 44382
rect 57820 43598 57822 43650
rect 57874 43598 57876 43650
rect 57820 43314 57876 43598
rect 57820 43262 57822 43314
rect 57874 43262 57876 43314
rect 57820 43250 57876 43262
rect 58156 43314 58212 43326
rect 58156 43262 58158 43314
rect 58210 43262 58212 43314
rect 58156 42194 58212 43262
rect 58156 42142 58158 42194
rect 58210 42142 58212 42194
rect 58156 40628 58212 42142
rect 57820 40626 58212 40628
rect 57820 40574 58158 40626
rect 58210 40574 58212 40626
rect 57820 40572 58212 40574
rect 57820 39842 57876 40572
rect 58156 40562 58212 40572
rect 57820 39790 57822 39842
rect 57874 39790 57876 39842
rect 57820 39778 57876 39790
rect 58380 40068 58436 40078
rect 57708 38434 57764 38444
rect 57820 38946 57876 38958
rect 57820 38894 57822 38946
rect 57874 38894 57876 38946
rect 57820 38276 57876 38894
rect 58044 38836 58100 38846
rect 58044 38388 58100 38780
rect 58044 38322 58100 38332
rect 58268 38500 58324 38510
rect 56028 37938 56084 37950
rect 56028 37886 56030 37938
rect 56082 37886 56084 37938
rect 56028 36260 56084 37886
rect 56700 37490 56756 37996
rect 56700 37438 56702 37490
rect 56754 37438 56756 37490
rect 56700 37426 56756 37438
rect 57596 38220 57876 38276
rect 56140 36596 56196 36606
rect 56140 36594 56644 36596
rect 56140 36542 56142 36594
rect 56194 36542 56644 36594
rect 56140 36540 56644 36542
rect 56140 36530 56196 36540
rect 56028 36194 56084 36204
rect 56588 35924 56644 36540
rect 57036 36484 57092 36494
rect 57036 36390 57092 36428
rect 57372 36484 57428 36494
rect 57372 36482 57540 36484
rect 57372 36430 57374 36482
rect 57426 36430 57540 36482
rect 57372 36428 57540 36430
rect 57372 36418 57428 36428
rect 56700 36372 56756 36382
rect 56700 36278 56756 36316
rect 57148 36260 57204 36270
rect 57148 36166 57204 36204
rect 56700 35924 56756 35934
rect 57260 35924 57316 35934
rect 56588 35922 57316 35924
rect 56588 35870 56702 35922
rect 56754 35870 57262 35922
rect 57314 35870 57316 35922
rect 56588 35868 57316 35870
rect 56700 35858 56756 35868
rect 57260 35858 57316 35868
rect 57484 35922 57540 36428
rect 57484 35870 57486 35922
rect 57538 35870 57540 35922
rect 57484 35858 57540 35870
rect 56476 35700 56532 35710
rect 56476 35606 56532 35644
rect 56812 35698 56868 35710
rect 56812 35646 56814 35698
rect 56866 35646 56868 35698
rect 56812 35364 56868 35646
rect 56812 35298 56868 35308
rect 56924 35700 56980 35710
rect 56924 34802 56980 35644
rect 57148 35698 57204 35710
rect 57148 35646 57150 35698
rect 57202 35646 57204 35698
rect 56924 34750 56926 34802
rect 56978 34750 56980 34802
rect 56924 34738 56980 34750
rect 57036 34804 57092 34814
rect 57148 34804 57204 35646
rect 57036 34802 57204 34804
rect 57036 34750 57038 34802
rect 57090 34750 57204 34802
rect 57036 34748 57204 34750
rect 57036 34738 57092 34748
rect 56700 34690 56756 34702
rect 56700 34638 56702 34690
rect 56754 34638 56756 34690
rect 56700 34242 56756 34638
rect 56700 34190 56702 34242
rect 56754 34190 56756 34242
rect 56700 34178 56756 34190
rect 56924 34132 56980 34142
rect 56812 34020 56868 34030
rect 56140 34018 56868 34020
rect 56140 33966 56814 34018
rect 56866 33966 56868 34018
rect 56140 33964 56868 33966
rect 56028 33122 56084 33134
rect 56028 33070 56030 33122
rect 56082 33070 56084 33122
rect 56028 32116 56084 33070
rect 56028 32050 56084 32060
rect 56028 31892 56084 31902
rect 56140 31892 56196 33964
rect 56812 33954 56868 33964
rect 56924 32900 56980 34076
rect 57036 34130 57092 34142
rect 57036 34078 57038 34130
rect 57090 34078 57092 34130
rect 57036 33570 57092 34078
rect 57036 33518 57038 33570
rect 57090 33518 57092 33570
rect 57036 33506 57092 33518
rect 57148 33460 57204 34748
rect 57260 34132 57316 34142
rect 57260 34038 57316 34076
rect 57596 33796 57652 38220
rect 58156 38164 58212 38174
rect 57820 38162 58212 38164
rect 57820 38110 58158 38162
rect 58210 38110 58212 38162
rect 57820 38108 58212 38110
rect 57820 35922 57876 38108
rect 58156 38098 58212 38108
rect 57932 36484 57988 36494
rect 57988 36428 58100 36484
rect 57932 36418 57988 36428
rect 57820 35870 57822 35922
rect 57874 35870 57876 35922
rect 57708 35698 57764 35710
rect 57708 35646 57710 35698
rect 57762 35646 57764 35698
rect 57708 35364 57764 35646
rect 57820 35700 57876 35870
rect 58044 35922 58100 36428
rect 58044 35870 58046 35922
rect 58098 35870 58100 35922
rect 58044 35858 58100 35870
rect 57820 35634 57876 35644
rect 57708 35298 57764 35308
rect 57596 33740 57764 33796
rect 57596 33572 57652 33582
rect 57148 33394 57204 33404
rect 57260 33570 57652 33572
rect 57260 33518 57598 33570
rect 57650 33518 57652 33570
rect 57260 33516 57652 33518
rect 57148 33236 57204 33246
rect 57148 33142 57204 33180
rect 57036 33124 57092 33134
rect 57036 33030 57092 33068
rect 56924 32844 57092 32900
rect 56028 31890 56196 31892
rect 56028 31838 56030 31890
rect 56082 31838 56196 31890
rect 56028 31836 56196 31838
rect 56028 31826 56084 31836
rect 56924 31220 56980 31230
rect 56028 31218 56980 31220
rect 56028 31166 56926 31218
rect 56978 31166 56980 31218
rect 56028 31164 56980 31166
rect 56028 30322 56084 31164
rect 56924 31154 56980 31164
rect 56588 30996 56644 31006
rect 56812 30996 56868 31006
rect 56588 30902 56644 30940
rect 56700 30994 56868 30996
rect 56700 30942 56814 30994
rect 56866 30942 56868 30994
rect 56700 30940 56868 30942
rect 56028 30270 56030 30322
rect 56082 30270 56084 30322
rect 56028 30258 56084 30270
rect 56700 29650 56756 30940
rect 56812 30930 56868 30940
rect 56924 30996 56980 31006
rect 57036 30996 57092 32844
rect 56980 30940 57092 30996
rect 57260 30994 57316 33516
rect 57596 33506 57652 33516
rect 57484 33348 57540 33358
rect 57484 33254 57540 33292
rect 57596 33124 57652 33134
rect 57596 33030 57652 33068
rect 57708 32788 57764 33740
rect 57260 30942 57262 30994
rect 57314 30942 57316 30994
rect 56924 30930 56980 30940
rect 57260 30930 57316 30942
rect 57484 32732 57764 32788
rect 58044 33124 58100 33134
rect 57036 29988 57092 29998
rect 56700 29598 56702 29650
rect 56754 29598 56756 29650
rect 56700 29586 56756 29598
rect 56924 29652 56980 29662
rect 56924 29558 56980 29596
rect 57036 29538 57092 29932
rect 57036 29486 57038 29538
rect 57090 29486 57092 29538
rect 57036 29474 57092 29486
rect 57372 29652 57428 29662
rect 56588 28756 56644 28794
rect 56588 28690 56644 28700
rect 56588 28532 56644 28542
rect 56588 28082 56644 28476
rect 56588 28030 56590 28082
rect 56642 28030 56644 28082
rect 56588 28018 56644 28030
rect 57372 28082 57428 29596
rect 57372 28030 57374 28082
rect 57426 28030 57428 28082
rect 57372 28018 57428 28030
rect 56924 27972 56980 27982
rect 57260 27972 57316 27982
rect 56700 27970 56980 27972
rect 56700 27918 56926 27970
rect 56978 27918 56980 27970
rect 56700 27916 56980 27918
rect 56028 26962 56084 26974
rect 56028 26910 56030 26962
rect 56082 26910 56084 26962
rect 56028 26516 56084 26910
rect 56700 26908 56756 27916
rect 56924 27906 56980 27916
rect 57148 27916 57260 27972
rect 56924 27636 56980 27646
rect 56028 26450 56084 26460
rect 56588 26852 56756 26908
rect 56812 27188 56868 27198
rect 56588 26292 56644 26852
rect 56476 26290 56644 26292
rect 56476 26238 56590 26290
rect 56642 26238 56644 26290
rect 56476 26236 56644 26238
rect 56364 25282 56420 25294
rect 56364 25230 56366 25282
rect 56418 25230 56420 25282
rect 56364 24724 56420 25230
rect 56476 25172 56532 26236
rect 56588 26226 56644 26236
rect 56812 25620 56868 27132
rect 56924 26290 56980 27580
rect 57036 26516 57092 26526
rect 57036 26422 57092 26460
rect 57148 26292 57204 27916
rect 57260 27878 57316 27916
rect 57372 27634 57428 27646
rect 57372 27582 57374 27634
rect 57426 27582 57428 27634
rect 57372 26908 57428 27582
rect 56924 26238 56926 26290
rect 56978 26238 56980 26290
rect 56924 26226 56980 26238
rect 57036 26236 57204 26292
rect 57260 26852 57428 26908
rect 57260 26290 57316 26852
rect 57260 26238 57262 26290
rect 57314 26238 57316 26290
rect 56588 25564 56868 25620
rect 56588 25394 56644 25564
rect 56588 25342 56590 25394
rect 56642 25342 56644 25394
rect 56588 25330 56644 25342
rect 56700 25396 56756 25406
rect 57036 25396 57092 26236
rect 57260 26226 57316 26238
rect 57484 25732 57540 32732
rect 58044 31892 58100 33068
rect 58156 32450 58212 32462
rect 58156 32398 58158 32450
rect 58210 32398 58212 32450
rect 58156 32116 58212 32398
rect 58156 32050 58212 32060
rect 58156 31892 58212 31902
rect 58044 31890 58212 31892
rect 58044 31838 58158 31890
rect 58210 31838 58212 31890
rect 58044 31836 58212 31838
rect 58156 31826 58212 31836
rect 58156 31444 58212 31454
rect 57820 31108 57876 31118
rect 58156 31108 58212 31388
rect 57596 31106 57876 31108
rect 57596 31054 57822 31106
rect 57874 31054 57876 31106
rect 57596 31052 57876 31054
rect 57596 26180 57652 31052
rect 57820 31042 57876 31052
rect 57932 31106 58212 31108
rect 57932 31054 58158 31106
rect 58210 31054 58212 31106
rect 57932 31052 58212 31054
rect 57708 29988 57764 29998
rect 57708 28196 57764 29932
rect 57820 29652 57876 29662
rect 57932 29652 57988 31052
rect 58156 31042 58212 31052
rect 57820 29650 57988 29652
rect 57820 29598 57822 29650
rect 57874 29598 57988 29650
rect 57820 29596 57988 29598
rect 58156 30322 58212 30334
rect 58156 30270 58158 30322
rect 58210 30270 58212 30322
rect 58156 29652 58212 30270
rect 57820 29586 57876 29596
rect 58156 29586 58212 29596
rect 58156 29316 58212 29326
rect 58044 29314 58212 29316
rect 58044 29262 58158 29314
rect 58210 29262 58212 29314
rect 58044 29260 58212 29262
rect 58044 28756 58100 29260
rect 58156 29250 58212 29260
rect 57708 28140 57876 28196
rect 57820 27858 57876 28140
rect 57932 27972 57988 27982
rect 57932 27878 57988 27916
rect 57820 27806 57822 27858
rect 57874 27806 57876 27858
rect 57820 26908 57876 27806
rect 57932 27636 57988 27646
rect 57932 27542 57988 27580
rect 57820 26852 57988 26908
rect 57596 26114 57652 26124
rect 57484 25666 57540 25676
rect 56700 25394 57092 25396
rect 56700 25342 56702 25394
rect 56754 25342 57092 25394
rect 56700 25340 57092 25342
rect 56476 25116 56644 25172
rect 56476 24724 56532 24734
rect 56364 24722 56532 24724
rect 56364 24670 56478 24722
rect 56530 24670 56532 24722
rect 56364 24668 56532 24670
rect 56476 24658 56532 24668
rect 56588 24724 56644 25116
rect 56588 24658 56644 24668
rect 55916 24434 55972 24444
rect 56700 24164 56756 25340
rect 57596 25284 57652 25294
rect 57596 25190 57652 25228
rect 57820 25282 57876 25294
rect 57820 25230 57822 25282
rect 57874 25230 57876 25282
rect 56812 24948 56868 24958
rect 56812 24946 57316 24948
rect 56812 24894 56814 24946
rect 56866 24894 57316 24946
rect 56812 24892 57316 24894
rect 56812 24882 56868 24892
rect 56924 24722 56980 24734
rect 56924 24670 56926 24722
rect 56978 24670 56980 24722
rect 56700 24108 56868 24164
rect 55132 24050 55188 24062
rect 55132 23998 55134 24050
rect 55186 23998 55188 24050
rect 55132 23380 55188 23998
rect 55132 23314 55188 23324
rect 56700 23380 56756 23390
rect 54124 23268 54180 23278
rect 54124 23174 54180 23212
rect 54348 23268 54404 23278
rect 56588 23268 56644 23278
rect 54348 23266 54964 23268
rect 54348 23214 54350 23266
rect 54402 23214 54964 23266
rect 54348 23212 54964 23214
rect 54348 23202 54404 23212
rect 53900 22978 53956 22988
rect 54012 23154 54068 23166
rect 54012 23102 54014 23154
rect 54066 23102 54068 23154
rect 54012 22820 54068 23102
rect 54684 23044 54740 23054
rect 54740 22988 54852 23044
rect 54684 22950 54740 22988
rect 53788 22764 54068 22820
rect 54572 22260 54628 22270
rect 54572 22166 54628 22204
rect 54684 22146 54740 22158
rect 54684 22094 54686 22146
rect 54738 22094 54740 22146
rect 54684 21812 54740 22094
rect 54348 21756 54740 21812
rect 54348 21698 54404 21756
rect 54348 21646 54350 21698
rect 54402 21646 54404 21698
rect 54348 21634 54404 21646
rect 54796 21588 54852 22988
rect 54908 22370 54964 23212
rect 56588 23174 56644 23212
rect 54908 22318 54910 22370
rect 54962 22318 54964 22370
rect 54908 22306 54964 22318
rect 55132 22258 55188 22270
rect 55132 22206 55134 22258
rect 55186 22206 55188 22258
rect 55132 22036 55188 22206
rect 56700 22258 56756 23324
rect 56812 22372 56868 24108
rect 56924 23378 56980 24670
rect 56924 23326 56926 23378
rect 56978 23326 56980 23378
rect 56924 23314 56980 23326
rect 57148 24724 57204 24734
rect 56812 22278 56868 22316
rect 56700 22206 56702 22258
rect 56754 22206 56756 22258
rect 56700 22194 56756 22206
rect 57036 22260 57092 22270
rect 57036 22166 57092 22204
rect 55132 21970 55188 21980
rect 56476 22146 56532 22158
rect 56476 22094 56478 22146
rect 56530 22094 56532 22146
rect 55132 21588 55188 21598
rect 55580 21588 55636 21598
rect 54796 21586 55636 21588
rect 54796 21534 55134 21586
rect 55186 21534 55582 21586
rect 55634 21534 55636 21586
rect 54796 21532 55636 21534
rect 55132 21522 55188 21532
rect 55244 20802 55300 21532
rect 55580 21522 55636 21532
rect 56476 21586 56532 22094
rect 56924 22148 56980 22158
rect 56924 21698 56980 22092
rect 56924 21646 56926 21698
rect 56978 21646 56980 21698
rect 56924 21634 56980 21646
rect 57148 22036 57204 24668
rect 57260 24050 57316 24892
rect 57820 24834 57876 25230
rect 57820 24782 57822 24834
rect 57874 24782 57876 24834
rect 57820 24770 57876 24782
rect 57260 23998 57262 24050
rect 57314 23998 57316 24050
rect 57260 23986 57316 23998
rect 57484 24610 57540 24622
rect 57484 24558 57486 24610
rect 57538 24558 57540 24610
rect 57484 23492 57540 24558
rect 57484 23426 57540 23436
rect 57932 23268 57988 26852
rect 57372 22372 57428 22382
rect 57372 22278 57428 22316
rect 57932 22370 57988 23212
rect 58044 26180 58100 28700
rect 58268 28532 58324 38444
rect 58268 28466 58324 28476
rect 58156 27972 58212 27982
rect 58156 27188 58212 27916
rect 58156 27094 58212 27132
rect 58380 26292 58436 40012
rect 58380 26226 58436 26236
rect 58156 26180 58212 26190
rect 58044 26178 58212 26180
rect 58044 26126 58158 26178
rect 58210 26126 58212 26178
rect 58044 26124 58212 26126
rect 58044 23938 58100 26124
rect 58156 26114 58212 26124
rect 58156 25394 58212 25406
rect 58156 25342 58158 25394
rect 58210 25342 58212 25394
rect 58156 25284 58212 25342
rect 58156 24500 58212 25228
rect 58156 24434 58212 24444
rect 58044 23886 58046 23938
rect 58098 23886 58100 23938
rect 58044 23044 58100 23886
rect 58156 23044 58212 23054
rect 58044 23042 58324 23044
rect 58044 22990 58158 23042
rect 58210 22990 58324 23042
rect 58044 22988 58324 22990
rect 58156 22978 58212 22988
rect 57932 22318 57934 22370
rect 57986 22318 57988 22370
rect 57932 22306 57988 22318
rect 57148 21698 57204 21980
rect 57260 22146 57316 22158
rect 57260 22094 57262 22146
rect 57314 22094 57316 22146
rect 57260 21924 57316 22094
rect 57596 22148 57652 22158
rect 57596 22054 57652 22092
rect 57820 22146 57876 22158
rect 57820 22094 57822 22146
rect 57874 22094 57876 22146
rect 57820 21924 57876 22094
rect 57260 21868 57876 21924
rect 57148 21646 57150 21698
rect 57202 21646 57204 21698
rect 57148 21634 57204 21646
rect 56476 21534 56478 21586
rect 56530 21534 56532 21586
rect 56476 21522 56532 21534
rect 56700 21476 56756 21486
rect 56588 21474 56756 21476
rect 56588 21422 56702 21474
rect 56754 21422 56756 21474
rect 56588 21420 56756 21422
rect 56588 21028 56644 21420
rect 56700 21410 56756 21420
rect 56028 20972 56644 21028
rect 56028 20914 56084 20972
rect 56028 20862 56030 20914
rect 56082 20862 56084 20914
rect 56028 20850 56084 20862
rect 57820 20916 57876 21868
rect 58156 20916 58212 20926
rect 57820 20914 58212 20916
rect 57820 20862 58158 20914
rect 58210 20862 58212 20914
rect 57820 20860 58212 20862
rect 58156 20850 58212 20860
rect 55244 20750 55246 20802
rect 55298 20750 55300 20802
rect 55244 20738 55300 20750
rect 58156 20244 58212 20254
rect 58268 20244 58324 22988
rect 58156 20242 58324 20244
rect 58156 20190 58158 20242
rect 58210 20190 58324 20242
rect 58156 20188 58324 20190
rect 58156 20178 58212 20188
rect 54908 19236 54964 19246
rect 52780 19010 52836 19022
rect 52780 18958 52782 19010
rect 52834 18958 52836 19010
rect 52668 18564 52724 18574
rect 52780 18564 52836 18958
rect 52668 18562 52836 18564
rect 52668 18510 52670 18562
rect 52722 18510 52836 18562
rect 52668 18508 52836 18510
rect 53788 19012 53844 19022
rect 52668 18340 52724 18508
rect 52668 18274 52724 18284
rect 52892 18450 52948 18462
rect 52892 18398 52894 18450
rect 52946 18398 52948 18450
rect 52780 17892 52836 17902
rect 52780 17798 52836 17836
rect 52668 17666 52724 17678
rect 52668 17614 52670 17666
rect 52722 17614 52724 17666
rect 52668 17108 52724 17614
rect 52668 17042 52724 17052
rect 52780 17444 52836 17454
rect 52668 16884 52724 16894
rect 52780 16884 52836 17388
rect 52892 17220 52948 18398
rect 53116 18450 53172 18462
rect 53116 18398 53118 18450
rect 53170 18398 53172 18450
rect 53116 17780 53172 18398
rect 53788 18450 53844 18956
rect 53788 18398 53790 18450
rect 53842 18398 53844 18450
rect 53788 18386 53844 18398
rect 53228 18340 53284 18350
rect 53228 18246 53284 18284
rect 53564 18338 53620 18350
rect 53564 18286 53566 18338
rect 53618 18286 53620 18338
rect 53564 18228 53620 18286
rect 54460 18340 54516 18350
rect 54460 18246 54516 18284
rect 53564 18162 53620 18172
rect 54124 18226 54180 18238
rect 54124 18174 54126 18226
rect 54178 18174 54180 18226
rect 54124 17892 54180 18174
rect 54572 18228 54628 18238
rect 54572 18134 54628 18172
rect 53340 17836 53732 17892
rect 53340 17780 53396 17836
rect 53116 17724 53340 17780
rect 53340 17714 53396 17724
rect 53340 17610 53396 17622
rect 53340 17558 53342 17610
rect 53394 17558 53396 17610
rect 53340 17556 53396 17558
rect 53228 17500 53396 17556
rect 53564 17556 53620 17566
rect 53116 17444 53172 17454
rect 53116 17350 53172 17388
rect 53228 17220 53284 17500
rect 53564 17462 53620 17500
rect 53452 17444 53508 17454
rect 53340 17442 53508 17444
rect 53340 17390 53454 17442
rect 53506 17390 53508 17442
rect 53340 17388 53508 17390
rect 53340 17332 53396 17388
rect 53452 17378 53508 17388
rect 53340 17266 53396 17276
rect 52892 17164 53284 17220
rect 52668 16882 52836 16884
rect 52668 16830 52670 16882
rect 52722 16830 52836 16882
rect 52668 16828 52836 16830
rect 52892 16884 52948 16894
rect 52668 16818 52724 16828
rect 52892 16790 52948 16828
rect 52556 16492 53060 16548
rect 52332 15446 52388 15484
rect 52556 15314 52612 15326
rect 52556 15262 52558 15314
rect 52610 15262 52612 15314
rect 52444 15202 52500 15214
rect 52444 15150 52446 15202
rect 52498 15150 52500 15202
rect 52444 14756 52500 15150
rect 52556 15204 52612 15262
rect 52556 15138 52612 15148
rect 52668 14756 52724 14766
rect 53004 14756 53060 16492
rect 53116 15148 53172 17164
rect 53564 16884 53620 16894
rect 53676 16884 53732 17836
rect 54124 17826 54180 17836
rect 54348 17780 54404 17790
rect 54348 17686 54404 17724
rect 54908 17668 54964 19180
rect 53564 16882 53732 16884
rect 53564 16830 53566 16882
rect 53618 16830 53732 16882
rect 53564 16828 53732 16830
rect 53788 17444 53844 17454
rect 53788 16884 53844 17388
rect 53564 16818 53620 16828
rect 53340 16772 53396 16782
rect 53340 16678 53396 16716
rect 53788 16770 53844 16828
rect 53788 16718 53790 16770
rect 53842 16718 53844 16770
rect 53788 16706 53844 16718
rect 54012 16772 54068 16782
rect 54012 16770 54404 16772
rect 54012 16718 54014 16770
rect 54066 16718 54404 16770
rect 54012 16716 54404 16718
rect 54012 16706 54068 16716
rect 54124 15202 54180 15214
rect 54124 15150 54126 15202
rect 54178 15150 54180 15202
rect 54124 15148 54180 15150
rect 53116 15092 53508 15148
rect 52444 14754 52724 14756
rect 52444 14702 52670 14754
rect 52722 14702 52724 14754
rect 52444 14700 52724 14702
rect 52668 14690 52724 14700
rect 52892 14700 53060 14756
rect 52780 14644 52836 14654
rect 52780 14550 52836 14588
rect 51884 13682 51940 13692
rect 52108 14140 52276 14196
rect 51660 12350 51662 12402
rect 51714 12350 51716 12402
rect 51660 12338 51716 12350
rect 52108 12402 52164 14140
rect 52668 13748 52724 13758
rect 52668 13654 52724 13692
rect 52780 13636 52836 13646
rect 52780 13542 52836 13580
rect 52892 13188 52948 14700
rect 53004 14532 53060 14542
rect 53004 13636 53060 14476
rect 53340 14420 53396 14430
rect 53452 14420 53508 15092
rect 53564 15092 53620 15102
rect 53564 14644 53620 15036
rect 53564 14530 53620 14588
rect 53676 15092 54180 15148
rect 54236 15092 54292 15102
rect 53676 14642 53732 15092
rect 54236 14998 54292 15036
rect 53676 14590 53678 14642
rect 53730 14590 53732 14642
rect 53676 14578 53732 14590
rect 54348 14644 54404 16716
rect 54908 16210 54964 17612
rect 55132 18338 55188 18350
rect 55132 18286 55134 18338
rect 55186 18286 55188 18338
rect 55132 17332 55188 18286
rect 55132 17266 55188 17276
rect 55244 18226 55300 18238
rect 55244 18174 55246 18226
rect 55298 18174 55300 18226
rect 55020 16884 55076 16894
rect 55076 16828 55188 16884
rect 55020 16818 55076 16828
rect 54908 16158 54910 16210
rect 54962 16158 54964 16210
rect 54908 16146 54964 16158
rect 55132 16212 55188 16828
rect 55244 16772 55300 18174
rect 56476 18228 56532 18238
rect 56476 17778 56532 18172
rect 56476 17726 56478 17778
rect 56530 17726 56532 17778
rect 56476 17714 56532 17726
rect 57820 18004 57876 18014
rect 57148 17668 57204 17678
rect 57204 17612 57540 17668
rect 57148 17574 57204 17612
rect 57484 17108 57540 17612
rect 57820 17554 57876 17948
rect 57820 17502 57822 17554
rect 57874 17502 57876 17554
rect 57820 17490 57876 17502
rect 58156 17556 58212 17566
rect 58212 17500 58324 17556
rect 58156 17462 58212 17500
rect 57484 17106 58100 17108
rect 57484 17054 57486 17106
rect 57538 17054 58100 17106
rect 57484 17052 58100 17054
rect 57484 17042 57540 17052
rect 55244 16706 55300 16716
rect 57372 16772 57428 16782
rect 55244 16212 55300 16222
rect 55132 16210 55300 16212
rect 55132 16158 55246 16210
rect 55298 16158 55300 16210
rect 55132 16156 55300 16158
rect 55244 16146 55300 16156
rect 57372 16210 57428 16716
rect 57372 16158 57374 16210
rect 57426 16158 57428 16210
rect 57372 16146 57428 16158
rect 54348 14550 54404 14588
rect 56476 15092 56532 15102
rect 56476 14642 56532 15036
rect 57708 14644 57764 17052
rect 58044 16098 58100 17052
rect 58268 17106 58324 17500
rect 58268 17054 58270 17106
rect 58322 17054 58324 17106
rect 58268 17042 58324 17054
rect 58044 16046 58046 16098
rect 58098 16046 58100 16098
rect 58044 16034 58100 16046
rect 56476 14590 56478 14642
rect 56530 14590 56532 14642
rect 56476 14578 56532 14590
rect 57260 14642 57764 14644
rect 57260 14590 57710 14642
rect 57762 14590 57764 14642
rect 57260 14588 57764 14590
rect 57260 14532 57316 14588
rect 57708 14578 57764 14588
rect 53564 14478 53566 14530
rect 53618 14478 53620 14530
rect 53564 14466 53620 14478
rect 56700 14530 57316 14532
rect 56700 14478 57262 14530
rect 57314 14478 57316 14530
rect 56700 14476 57316 14478
rect 53396 14364 53508 14420
rect 53340 14326 53396 14364
rect 53116 14308 53172 14318
rect 53116 14214 53172 14252
rect 56700 13970 56756 14476
rect 57260 14466 57316 14476
rect 56700 13918 56702 13970
rect 56754 13918 56756 13970
rect 55356 13748 55412 13758
rect 53116 13636 53172 13646
rect 53004 13634 53172 13636
rect 53004 13582 53118 13634
rect 53170 13582 53172 13634
rect 53004 13580 53172 13582
rect 53116 13570 53172 13580
rect 55244 13636 55300 13646
rect 55244 13542 55300 13580
rect 52108 12350 52110 12402
rect 52162 12350 52164 12402
rect 51324 12178 51380 12190
rect 51324 12126 51326 12178
rect 51378 12126 51380 12178
rect 51324 11620 51380 12126
rect 51884 12178 51940 12190
rect 51884 12126 51886 12178
rect 51938 12126 51940 12178
rect 51324 11554 51380 11564
rect 51660 11956 51716 11966
rect 50988 11394 51268 11396
rect 50988 11342 50990 11394
rect 51042 11342 51268 11394
rect 50988 11340 51268 11342
rect 50988 11330 51044 11340
rect 51324 11284 51380 11294
rect 51548 11284 51604 11294
rect 51324 11282 51604 11284
rect 51324 11230 51326 11282
rect 51378 11230 51550 11282
rect 51602 11230 51604 11282
rect 51324 11228 51604 11230
rect 51324 11218 51380 11228
rect 51548 11218 51604 11228
rect 51100 11170 51156 11182
rect 51100 11118 51102 11170
rect 51154 11118 51156 11170
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50204 10670 50206 10722
rect 50258 10670 50260 10722
rect 49532 10388 49588 10444
rect 49532 10322 49588 10332
rect 50204 10052 50260 10670
rect 50652 10500 50708 10510
rect 51100 10500 51156 11118
rect 51660 11060 51716 11900
rect 51884 11394 51940 12126
rect 52108 12068 52164 12350
rect 52780 13132 52948 13188
rect 52220 12292 52276 12302
rect 52220 12198 52276 12236
rect 52668 12292 52724 12302
rect 52668 12198 52724 12236
rect 52108 12012 52724 12068
rect 52668 11506 52724 12012
rect 52668 11454 52670 11506
rect 52722 11454 52724 11506
rect 52668 11442 52724 11454
rect 52108 11396 52164 11406
rect 51884 11342 51886 11394
rect 51938 11342 51940 11394
rect 51884 11330 51940 11342
rect 51996 11340 52108 11396
rect 51772 11284 51828 11294
rect 51772 11170 51828 11228
rect 51772 11118 51774 11170
rect 51826 11118 51828 11170
rect 51772 11106 51828 11118
rect 50708 10444 51156 10500
rect 51324 11004 51716 11060
rect 51324 10722 51380 11004
rect 51996 10836 52052 11340
rect 52108 11302 52164 11340
rect 52780 11396 52836 13132
rect 52892 12964 52948 12974
rect 52948 12908 53284 12964
rect 52892 12870 52948 12908
rect 53228 12178 53284 12908
rect 53228 12126 53230 12178
rect 53282 12126 53284 12178
rect 53228 12114 53284 12126
rect 55356 12066 55412 13692
rect 56028 13748 56084 13758
rect 56028 13654 56084 13692
rect 56700 13748 56756 13918
rect 56700 13682 56756 13692
rect 55356 12014 55358 12066
rect 55410 12014 55412 12066
rect 55356 11620 55412 12014
rect 55356 11554 55412 11564
rect 57260 11732 57316 11742
rect 57260 11618 57316 11676
rect 57260 11566 57262 11618
rect 57314 11566 57316 11618
rect 57260 11554 57316 11566
rect 52780 11330 52836 11340
rect 55580 11508 55636 11518
rect 55580 11394 55636 11452
rect 56028 11508 56084 11518
rect 56028 11414 56084 11452
rect 55580 11342 55582 11394
rect 55634 11342 55636 11394
rect 54796 11284 54852 11294
rect 54796 11190 54852 11228
rect 52052 10780 52164 10836
rect 51996 10742 52052 10780
rect 51324 10670 51326 10722
rect 51378 10670 51380 10722
rect 50652 10406 50708 10444
rect 50204 9986 50260 9996
rect 50764 9828 50820 9838
rect 50204 9826 50820 9828
rect 50204 9774 50766 9826
rect 50818 9774 50820 9826
rect 50204 9772 50820 9774
rect 47292 9202 47348 9212
rect 49756 9268 49812 9278
rect 49756 9042 49812 9212
rect 49756 8990 49758 9042
rect 49810 8990 49812 9042
rect 47628 8930 47684 8942
rect 47628 8878 47630 8930
rect 47682 8878 47684 8930
rect 46844 8372 47236 8428
rect 46620 8034 46676 8046
rect 46620 7982 46622 8034
rect 46674 7982 46676 8034
rect 46620 7812 46676 7982
rect 46620 7746 46676 7756
rect 46396 6802 46564 6804
rect 46396 6750 46398 6802
rect 46450 6750 46564 6802
rect 46396 6748 46564 6750
rect 46396 6580 46452 6748
rect 46844 6692 46900 8372
rect 47180 8260 47236 8372
rect 47404 8372 47460 8382
rect 46396 6514 46452 6524
rect 46732 6690 46900 6692
rect 46732 6638 46846 6690
rect 46898 6638 46900 6690
rect 46732 6636 46900 6638
rect 46732 6244 46788 6636
rect 46844 6626 46900 6636
rect 46956 8204 47236 8260
rect 47292 8260 47348 8270
rect 47404 8260 47460 8316
rect 47292 8258 47460 8260
rect 47292 8206 47294 8258
rect 47346 8206 47460 8258
rect 47292 8204 47460 8206
rect 47516 8370 47572 8382
rect 47516 8318 47518 8370
rect 47570 8318 47572 8370
rect 46956 6468 47012 8204
rect 47292 8148 47348 8204
rect 47292 8082 47348 8092
rect 47516 8148 47572 8318
rect 47628 8260 47684 8878
rect 49756 8428 49812 8990
rect 50204 9266 50260 9772
rect 50764 9762 50820 9772
rect 50876 9714 50932 10444
rect 51212 10052 51268 10062
rect 50876 9662 50878 9714
rect 50930 9662 50932 9714
rect 50428 9604 50484 9614
rect 50876 9604 50932 9662
rect 51100 9716 51156 9726
rect 51100 9622 51156 9660
rect 50428 9602 50932 9604
rect 50428 9550 50430 9602
rect 50482 9550 50932 9602
rect 50428 9548 50932 9550
rect 50428 9538 50484 9548
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50204 9214 50206 9266
rect 50258 9214 50260 9266
rect 48636 8372 48692 8382
rect 48524 8260 48580 8270
rect 47628 8166 47684 8204
rect 48412 8258 48580 8260
rect 48412 8206 48526 8258
rect 48578 8206 48580 8258
rect 48412 8204 48580 8206
rect 47516 8082 47572 8092
rect 47964 8146 48020 8158
rect 47964 8094 47966 8146
rect 48018 8094 48020 8146
rect 47964 7700 48020 8094
rect 47964 7634 48020 7644
rect 48300 8146 48356 8158
rect 48300 8094 48302 8146
rect 48354 8094 48356 8146
rect 46284 6188 46788 6244
rect 46844 6412 47012 6468
rect 47180 6580 47236 6590
rect 46284 6130 46340 6188
rect 46284 6078 46286 6130
rect 46338 6078 46340 6130
rect 46284 6066 46340 6078
rect 46060 6018 46228 6020
rect 46060 5966 46174 6018
rect 46226 5966 46228 6018
rect 46060 5964 46228 5966
rect 45052 5814 45108 5852
rect 45276 5906 45332 5918
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45164 5794 45220 5806
rect 45164 5742 45166 5794
rect 45218 5742 45220 5794
rect 44940 5684 44996 5694
rect 44940 5234 44996 5628
rect 44940 5182 44942 5234
rect 44994 5182 44996 5234
rect 44940 5170 44996 5182
rect 44604 5058 44660 5068
rect 44940 4452 44996 4462
rect 45164 4452 45220 5742
rect 45276 5684 45332 5854
rect 45612 5908 45668 5918
rect 45612 5906 45780 5908
rect 45612 5854 45614 5906
rect 45666 5854 45780 5906
rect 45612 5852 45780 5854
rect 45612 5842 45668 5852
rect 45276 5618 45332 5628
rect 45500 5124 45556 5134
rect 45500 5030 45556 5068
rect 45724 4900 45780 5852
rect 45836 5124 45892 5134
rect 46060 5124 46116 5964
rect 46172 5954 46228 5964
rect 46508 6020 46564 6030
rect 46508 5926 46564 5964
rect 46732 5908 46788 5918
rect 46732 5814 46788 5852
rect 45836 5122 46116 5124
rect 45836 5070 45838 5122
rect 45890 5070 46116 5122
rect 45836 5068 46116 5070
rect 46396 5124 46452 5134
rect 45836 5058 45892 5068
rect 46396 5030 46452 5068
rect 45948 4900 46004 4910
rect 45724 4898 46004 4900
rect 45724 4846 45950 4898
rect 46002 4846 46004 4898
rect 45724 4844 46004 4846
rect 45948 4834 46004 4844
rect 46060 4898 46116 4910
rect 46060 4846 46062 4898
rect 46114 4846 46116 4898
rect 44940 4450 45220 4452
rect 44940 4398 44942 4450
rect 44994 4398 45220 4450
rect 44940 4396 45220 4398
rect 44940 4386 44996 4396
rect 44156 4340 44212 4350
rect 43820 4174 43822 4226
rect 43874 4174 43876 4226
rect 34300 4162 34356 4172
rect 43820 4162 43876 4174
rect 43932 4338 44212 4340
rect 43932 4286 44158 4338
rect 44210 4286 44212 4338
rect 43932 4284 44212 4286
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 21644 3614 21646 3666
rect 21698 3614 21700 3666
rect 21644 3602 21700 3614
rect 43932 3666 43988 4284
rect 44156 4274 44212 4284
rect 46060 4228 46116 4846
rect 46844 4340 46900 6412
rect 46956 6018 47012 6030
rect 46956 5966 46958 6018
rect 47010 5966 47012 6018
rect 46956 4564 47012 5966
rect 47068 6020 47124 6030
rect 47068 5926 47124 5964
rect 47180 6018 47236 6524
rect 48300 6132 48356 8094
rect 48412 6690 48468 8204
rect 48524 8194 48580 8204
rect 48412 6638 48414 6690
rect 48466 6638 48468 6690
rect 48412 6468 48468 6638
rect 48412 6402 48468 6412
rect 48524 6578 48580 6590
rect 48524 6526 48526 6578
rect 48578 6526 48580 6578
rect 48300 6066 48356 6076
rect 47180 5966 47182 6018
rect 47234 5966 47236 6018
rect 47180 5954 47236 5966
rect 47516 5796 47572 5806
rect 47516 5794 47796 5796
rect 47516 5742 47518 5794
rect 47570 5742 47796 5794
rect 47516 5740 47796 5742
rect 47516 5730 47572 5740
rect 47740 5234 47796 5740
rect 47740 5182 47742 5234
rect 47794 5182 47796 5234
rect 47740 5170 47796 5182
rect 47068 5124 47124 5134
rect 47068 5030 47124 5068
rect 46956 4498 47012 4508
rect 46956 4340 47012 4350
rect 46844 4284 46956 4340
rect 46956 4274 47012 4284
rect 46060 4162 46116 4172
rect 47068 4228 47124 4238
rect 47068 4134 47124 4172
rect 48524 4228 48580 6526
rect 48636 6580 48692 8316
rect 49644 8372 49700 8382
rect 49756 8372 50148 8428
rect 48748 8258 48804 8270
rect 48748 8206 48750 8258
rect 48802 8206 48804 8258
rect 48748 7700 48804 8206
rect 48972 8260 49028 8270
rect 48972 8166 49028 8204
rect 49644 8258 49700 8316
rect 49644 8206 49646 8258
rect 49698 8206 49700 8258
rect 49644 8194 49700 8206
rect 49980 8146 50036 8158
rect 49980 8094 49982 8146
rect 50034 8094 50036 8146
rect 49420 8036 49476 8046
rect 49420 7942 49476 7980
rect 48748 7634 48804 7644
rect 49644 7474 49700 7486
rect 49644 7422 49646 7474
rect 49698 7422 49700 7474
rect 48748 6804 48804 6814
rect 49644 6804 49700 7422
rect 49868 7476 49924 7486
rect 49868 7382 49924 7420
rect 49756 7364 49812 7374
rect 49756 7270 49812 7308
rect 49980 6916 50036 8094
rect 50092 7698 50148 8372
rect 50204 8372 50260 9214
rect 50428 9042 50484 9054
rect 50428 8990 50430 9042
rect 50482 8990 50484 9042
rect 50204 8278 50260 8316
rect 50316 8930 50372 8942
rect 50316 8878 50318 8930
rect 50370 8878 50372 8930
rect 50092 7646 50094 7698
rect 50146 7646 50148 7698
rect 50092 7634 50148 7646
rect 50316 7476 50372 8878
rect 50428 8148 50484 8990
rect 51100 8372 51156 8382
rect 51100 8278 51156 8316
rect 50764 8260 50820 8270
rect 50764 8166 50820 8204
rect 50428 8082 50484 8092
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50876 7588 50932 7598
rect 51212 7588 51268 9996
rect 51324 9716 51380 10670
rect 51436 10722 51492 10734
rect 51436 10670 51438 10722
rect 51490 10670 51492 10722
rect 51436 9940 51492 10670
rect 51436 9874 51492 9884
rect 51660 10610 51716 10622
rect 51660 10558 51662 10610
rect 51714 10558 51716 10610
rect 51660 9828 51716 10558
rect 52108 10164 52164 10780
rect 52108 9938 52164 10108
rect 53228 10164 53284 10174
rect 52108 9886 52110 9938
rect 52162 9886 52164 9938
rect 52108 9874 52164 9886
rect 52332 9940 52388 9950
rect 51660 9762 51716 9772
rect 51436 9716 51492 9726
rect 51324 9714 51492 9716
rect 51324 9662 51438 9714
rect 51490 9662 51492 9714
rect 51324 9660 51492 9662
rect 51436 9650 51492 9660
rect 52332 8930 52388 9884
rect 52556 9826 52612 9838
rect 52556 9774 52558 9826
rect 52610 9774 52612 9826
rect 52556 9716 52612 9774
rect 52892 9828 52948 9866
rect 52892 9762 52948 9772
rect 53228 9826 53284 10108
rect 53228 9774 53230 9826
rect 53282 9774 53284 9826
rect 53228 9762 53284 9774
rect 52556 9650 52612 9660
rect 52892 9604 52948 9614
rect 52892 9510 52948 9548
rect 54460 9604 54516 9614
rect 54460 9154 54516 9548
rect 54460 9102 54462 9154
rect 54514 9102 54516 9154
rect 54460 9090 54516 9102
rect 55580 9268 55636 11342
rect 57372 11284 57428 11294
rect 57820 11284 57876 11294
rect 57372 11282 57876 11284
rect 57372 11230 57374 11282
rect 57426 11230 57822 11282
rect 57874 11230 57876 11282
rect 57372 11228 57876 11230
rect 57372 11218 57428 11228
rect 57820 11218 57876 11228
rect 58156 11282 58212 11294
rect 58156 11230 58158 11282
rect 58210 11230 58212 11282
rect 58156 10612 58212 11230
rect 58156 10518 58212 10556
rect 55692 9268 55748 9278
rect 55580 9266 55748 9268
rect 55580 9214 55694 9266
rect 55746 9214 55748 9266
rect 55580 9212 55748 9214
rect 52332 8878 52334 8930
rect 52386 8878 52388 8930
rect 52332 8428 52388 8878
rect 55244 9042 55300 9054
rect 55244 8990 55246 9042
rect 55298 8990 55300 9042
rect 55244 8932 55300 8990
rect 55580 8932 55636 9212
rect 55244 8876 55636 8932
rect 51996 8372 52388 8428
rect 51324 8258 51380 8270
rect 51324 8206 51326 8258
rect 51378 8206 51380 8258
rect 51324 8148 51380 8206
rect 51996 8260 52052 8372
rect 51996 8194 52052 8204
rect 51324 8082 51380 8092
rect 51660 8034 51716 8046
rect 51660 7982 51662 8034
rect 51714 7982 51716 8034
rect 50764 7532 50876 7588
rect 50540 7476 50596 7486
rect 50316 7474 50596 7476
rect 50316 7422 50542 7474
rect 50594 7422 50596 7474
rect 50316 7420 50596 7422
rect 50540 7410 50596 7420
rect 50652 7476 50708 7486
rect 50092 7364 50148 7374
rect 50148 7308 50372 7364
rect 50092 7298 50148 7308
rect 49868 6860 50036 6916
rect 50316 6914 50372 7308
rect 50316 6862 50318 6914
rect 50370 6862 50372 6914
rect 49756 6804 49812 6814
rect 48748 6802 49812 6804
rect 48748 6750 48750 6802
rect 48802 6750 49758 6802
rect 49810 6750 49812 6802
rect 48748 6748 49812 6750
rect 48748 6738 48804 6748
rect 49756 6738 49812 6748
rect 48860 6580 48916 6590
rect 48636 6578 48916 6580
rect 48636 6526 48862 6578
rect 48914 6526 48916 6578
rect 48636 6524 48916 6526
rect 48860 6514 48916 6524
rect 49420 6580 49476 6590
rect 49420 6486 49476 6524
rect 49868 5236 49924 6860
rect 50316 6850 50372 6862
rect 50204 6804 50260 6814
rect 49980 6748 50204 6804
rect 49980 6690 50036 6748
rect 50204 6738 50260 6748
rect 50428 6802 50484 6814
rect 50428 6750 50430 6802
rect 50482 6750 50484 6802
rect 49980 6638 49982 6690
rect 50034 6638 50036 6690
rect 49980 6626 50036 6638
rect 50428 6692 50484 6750
rect 50652 6804 50708 7420
rect 50652 6738 50708 6748
rect 50428 6626 50484 6636
rect 50764 6578 50820 7532
rect 50876 7494 50932 7532
rect 51100 7586 51268 7588
rect 51100 7534 51214 7586
rect 51266 7534 51268 7586
rect 51100 7532 51268 7534
rect 50988 6692 51044 6702
rect 51100 6692 51156 7532
rect 51212 7522 51268 7532
rect 51436 7700 51492 7710
rect 51436 7474 51492 7644
rect 51436 7422 51438 7474
rect 51490 7422 51492 7474
rect 51436 6804 51492 7422
rect 51660 7476 51716 7982
rect 51660 7410 51716 7420
rect 51548 7364 51604 7374
rect 51548 7270 51604 7308
rect 52444 7364 52500 7374
rect 52444 7270 52500 7308
rect 52556 7250 52612 7262
rect 52556 7198 52558 7250
rect 52610 7198 52612 7250
rect 51548 6804 51604 6814
rect 51436 6748 51548 6804
rect 51548 6738 51604 6748
rect 50988 6690 51156 6692
rect 50988 6638 50990 6690
rect 51042 6638 51156 6690
rect 50988 6636 51156 6638
rect 52556 6692 52612 7198
rect 52668 6804 52724 6814
rect 52668 6710 52724 6748
rect 50988 6626 51044 6636
rect 52556 6626 52612 6636
rect 54796 6692 54852 6702
rect 54796 6598 54852 6636
rect 55468 6692 55524 6702
rect 55692 6692 55748 9212
rect 56028 6692 56084 6702
rect 55468 6690 56084 6692
rect 55468 6638 55470 6690
rect 55522 6638 56030 6690
rect 56082 6638 56084 6690
rect 55468 6636 56084 6638
rect 50764 6526 50766 6578
rect 50818 6526 50820 6578
rect 50764 6514 50820 6526
rect 51212 6578 51268 6590
rect 51212 6526 51214 6578
rect 51266 6526 51268 6578
rect 48860 5234 49924 5236
rect 48860 5182 49870 5234
rect 49922 5182 49924 5234
rect 48860 5180 49924 5182
rect 48748 4564 48804 4574
rect 48748 4470 48804 4508
rect 48860 4450 48916 5180
rect 49868 5170 49924 5180
rect 50428 6468 50484 6478
rect 50316 5124 50372 5134
rect 50316 5030 50372 5068
rect 48860 4398 48862 4450
rect 48914 4398 48916 4450
rect 48860 4386 48916 4398
rect 50428 4228 50484 6412
rect 51100 6466 51156 6478
rect 51100 6414 51102 6466
rect 51154 6414 51156 6466
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 51100 5236 51156 6414
rect 51212 6468 51268 6526
rect 51212 6402 51268 6412
rect 51212 5236 51268 5246
rect 51100 5234 51268 5236
rect 51100 5182 51214 5234
rect 51266 5182 51268 5234
rect 51100 5180 51268 5182
rect 51212 5170 51268 5180
rect 53340 5012 53396 5022
rect 51324 4900 51380 4910
rect 51324 4806 51380 4844
rect 52668 4900 52724 4910
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 52668 4450 52724 4844
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 53340 4564 53396 4956
rect 55468 5012 55524 6636
rect 56028 6626 56084 6636
rect 55468 4946 55524 4956
rect 53900 4564 53956 4574
rect 53340 4562 53956 4564
rect 53340 4510 53902 4562
rect 53954 4510 53956 4562
rect 53340 4508 53956 4510
rect 53340 4338 53396 4508
rect 53900 4498 53956 4508
rect 53340 4286 53342 4338
rect 53394 4286 53396 4338
rect 53340 4274 53396 4286
rect 57596 4340 57652 4350
rect 57596 4246 57652 4284
rect 58156 4338 58212 4350
rect 58156 4286 58158 4338
rect 58210 4286 58212 4338
rect 50540 4228 50596 4238
rect 50428 4226 50596 4228
rect 50428 4174 50542 4226
rect 50594 4174 50596 4226
rect 50428 4172 50596 4174
rect 48524 4162 48580 4172
rect 50540 4162 50596 4172
rect 57372 4228 57428 4238
rect 57372 4134 57428 4172
rect 58156 4228 58212 4286
rect 43932 3614 43934 3666
rect 43986 3614 43988 3666
rect 43932 3602 43988 3614
rect 58156 3668 58212 4172
rect 58156 3602 58212 3612
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
<< via2 >>
rect 4732 66780 4788 66836
rect 5516 66780 5572 66836
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 8764 64652 8820 64708
rect 5740 63868 5796 63924
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 10108 64818 10164 64820
rect 10108 64766 10110 64818
rect 10110 64766 10162 64818
rect 10162 64766 10164 64818
rect 10108 64764 10164 64766
rect 9436 64706 9492 64708
rect 9436 64654 9438 64706
rect 9438 64654 9490 64706
rect 9490 64654 9492 64706
rect 9436 64652 9492 64654
rect 11340 64540 11396 64596
rect 8764 63868 8820 63924
rect 6524 63026 6580 63028
rect 6524 62974 6526 63026
rect 6526 62974 6578 63026
rect 6578 62974 6580 63026
rect 6524 62972 6580 62974
rect 7308 62972 7364 63028
rect 7644 63026 7700 63028
rect 7644 62974 7646 63026
rect 7646 62974 7698 63026
rect 7698 62974 7700 63026
rect 7644 62972 7700 62974
rect 6748 62300 6804 62356
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 7868 62466 7924 62468
rect 7868 62414 7870 62466
rect 7870 62414 7922 62466
rect 7922 62414 7924 62466
rect 7868 62412 7924 62414
rect 8540 62578 8596 62580
rect 8540 62526 8542 62578
rect 8542 62526 8594 62578
rect 8594 62526 8596 62578
rect 8540 62524 8596 62526
rect 7084 62354 7140 62356
rect 7084 62302 7086 62354
rect 7086 62302 7138 62354
rect 7138 62302 7140 62354
rect 7084 62300 7140 62302
rect 7980 62300 8036 62356
rect 6188 61346 6244 61348
rect 6188 61294 6190 61346
rect 6190 61294 6242 61346
rect 6242 61294 6244 61346
rect 6188 61292 6244 61294
rect 2828 60060 2884 60116
rect 1708 58322 1764 58324
rect 1708 58270 1710 58322
rect 1710 58270 1762 58322
rect 1762 58270 1764 58322
rect 1708 58268 1764 58270
rect 1820 57708 1876 57764
rect 1820 47516 1876 47572
rect 2492 58156 2548 58212
rect 5628 60674 5684 60676
rect 5628 60622 5630 60674
rect 5630 60622 5682 60674
rect 5682 60622 5684 60674
rect 5628 60620 5684 60622
rect 6300 60620 6356 60676
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 6860 61346 6916 61348
rect 6860 61294 6862 61346
rect 6862 61294 6914 61346
rect 6914 61294 6916 61346
rect 6860 61292 6916 61294
rect 3500 59388 3556 59444
rect 5852 59778 5908 59780
rect 5852 59726 5854 59778
rect 5854 59726 5906 59778
rect 5906 59726 5908 59778
rect 5852 59724 5908 59726
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 2828 57708 2884 57764
rect 3948 58210 4004 58212
rect 3948 58158 3950 58210
rect 3950 58158 4002 58210
rect 4002 58158 4004 58210
rect 3948 58156 4004 58158
rect 3836 57708 3892 57764
rect 4060 56812 4116 56868
rect 4172 57708 4228 57764
rect 5516 58156 5572 58212
rect 5068 58044 5124 58100
rect 4956 57762 5012 57764
rect 4956 57710 4958 57762
rect 4958 57710 5010 57762
rect 5010 57710 5012 57762
rect 4956 57708 5012 57710
rect 4620 57538 4676 57540
rect 4620 57486 4622 57538
rect 4622 57486 4674 57538
rect 4674 57486 4676 57538
rect 4620 57484 4676 57486
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4508 56866 4564 56868
rect 4508 56814 4510 56866
rect 4510 56814 4562 56866
rect 4562 56814 4564 56866
rect 4508 56812 4564 56814
rect 4844 56812 4900 56868
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4396 55468 4452 55524
rect 5740 58210 5796 58212
rect 5740 58158 5742 58210
rect 5742 58158 5794 58210
rect 5794 58158 5796 58210
rect 5740 58156 5796 58158
rect 5852 58044 5908 58100
rect 5628 57484 5684 57540
rect 5516 56866 5572 56868
rect 5516 56814 5518 56866
rect 5518 56814 5570 56866
rect 5570 56814 5572 56866
rect 5516 56812 5572 56814
rect 5852 57036 5908 57092
rect 6188 57036 6244 57092
rect 5292 56700 5348 56756
rect 5068 55580 5124 55636
rect 2828 55020 2884 55076
rect 3052 55020 3108 55076
rect 3724 55074 3780 55076
rect 3724 55022 3726 55074
rect 3726 55022 3778 55074
rect 3778 55022 3780 55074
rect 3724 55020 3780 55022
rect 3164 54572 3220 54628
rect 3948 54572 4004 54628
rect 4620 54460 4676 54516
rect 3388 53900 3444 53956
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4284 53900 4340 53956
rect 4284 52668 4340 52724
rect 5180 54514 5236 54516
rect 5180 54462 5182 54514
rect 5182 54462 5234 54514
rect 5234 54462 5236 54514
rect 5180 54460 5236 54462
rect 6860 56812 6916 56868
rect 6636 56700 6692 56756
rect 6188 55468 6244 55524
rect 6636 55580 6692 55636
rect 5404 54626 5460 54628
rect 5404 54574 5406 54626
rect 5406 54574 5458 54626
rect 5458 54574 5460 54626
rect 5404 54572 5460 54574
rect 4956 52668 5012 52724
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3948 52220 4004 52276
rect 4620 52274 4676 52276
rect 4620 52222 4622 52274
rect 4622 52222 4674 52274
rect 4674 52222 4676 52274
rect 4620 52220 4676 52222
rect 3388 51490 3444 51492
rect 3388 51438 3390 51490
rect 3390 51438 3442 51490
rect 3442 51438 3444 51490
rect 3388 51436 3444 51438
rect 3276 51212 3332 51268
rect 2492 49980 2548 50036
rect 3612 50540 3668 50596
rect 2716 46562 2772 46564
rect 2716 46510 2718 46562
rect 2718 46510 2770 46562
rect 2770 46510 2772 46562
rect 2716 46508 2772 46510
rect 3388 46562 3444 46564
rect 3388 46510 3390 46562
rect 3390 46510 3442 46562
rect 3442 46510 3444 46562
rect 3388 46508 3444 46510
rect 3388 44380 3444 44436
rect 2380 43708 2436 43764
rect 1820 43538 1876 43540
rect 1820 43486 1822 43538
rect 1822 43486 1874 43538
rect 1874 43486 1876 43538
rect 1820 43484 1876 43486
rect 1820 39676 1876 39732
rect 1820 35026 1876 35028
rect 1820 34974 1822 35026
rect 1822 34974 1874 35026
rect 1874 34974 1876 35026
rect 1820 34972 1876 34974
rect 2604 43708 2660 43764
rect 3612 43484 3668 43540
rect 3612 42924 3668 42980
rect 2828 41692 2884 41748
rect 3276 41692 3332 41748
rect 5068 51436 5124 51492
rect 3948 51212 4004 51268
rect 3948 50652 4004 50708
rect 4396 51378 4452 51380
rect 4396 51326 4398 51378
rect 4398 51326 4450 51378
rect 4450 51326 4452 51378
rect 4396 51324 4452 51326
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4172 50428 4228 50484
rect 5964 53452 6020 53508
rect 5516 50652 5572 50708
rect 5628 50594 5684 50596
rect 5628 50542 5630 50594
rect 5630 50542 5682 50594
rect 5682 50542 5684 50594
rect 5628 50540 5684 50542
rect 5740 50482 5796 50484
rect 5740 50430 5742 50482
rect 5742 50430 5794 50482
rect 5794 50430 5796 50482
rect 5740 50428 5796 50430
rect 4284 50316 4340 50372
rect 4732 50204 4788 50260
rect 4508 50034 4564 50036
rect 4508 49982 4510 50034
rect 4510 49982 4562 50034
rect 4562 49982 4564 50034
rect 4508 49980 4564 49982
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 5404 48972 5460 49028
rect 4956 48130 5012 48132
rect 4956 48078 4958 48130
rect 4958 48078 5010 48130
rect 5010 48078 5012 48130
rect 4956 48076 5012 48078
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 6076 49026 6132 49028
rect 6076 48974 6078 49026
rect 6078 48974 6130 49026
rect 6130 48974 6132 49026
rect 6076 48972 6132 48974
rect 5628 48076 5684 48132
rect 5068 47570 5124 47572
rect 5068 47518 5070 47570
rect 5070 47518 5122 47570
rect 5122 47518 5124 47570
rect 5068 47516 5124 47518
rect 4620 47292 4676 47348
rect 5292 47292 5348 47348
rect 5404 46956 5460 47012
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4508 44380 4564 44436
rect 4844 44268 4900 44324
rect 5180 44492 5236 44548
rect 5740 47346 5796 47348
rect 5740 47294 5742 47346
rect 5742 47294 5794 47346
rect 5794 47294 5796 47346
rect 5740 47292 5796 47294
rect 6188 46956 6244 47012
rect 6076 45106 6132 45108
rect 6076 45054 6078 45106
rect 6078 45054 6130 45106
rect 6130 45054 6132 45106
rect 6076 45052 6132 45054
rect 5628 44434 5684 44436
rect 5628 44382 5630 44434
rect 5630 44382 5682 44434
rect 5682 44382 5684 44434
rect 5628 44380 5684 44382
rect 5964 44434 6020 44436
rect 5964 44382 5966 44434
rect 5966 44382 6018 44434
rect 6018 44382 6020 44434
rect 5964 44380 6020 44382
rect 6188 44322 6244 44324
rect 6188 44270 6190 44322
rect 6190 44270 6242 44322
rect 6242 44270 6244 44322
rect 6188 44268 6244 44270
rect 5068 43484 5124 43540
rect 5516 43650 5572 43652
rect 5516 43598 5518 43650
rect 5518 43598 5570 43650
rect 5570 43598 5572 43650
rect 5516 43596 5572 43598
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 3948 42924 4004 42980
rect 3052 40460 3108 40516
rect 4060 40460 4116 40516
rect 3948 40402 4004 40404
rect 3948 40350 3950 40402
rect 3950 40350 4002 40402
rect 4002 40350 4004 40402
rect 3948 40348 4004 40350
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4284 40908 4340 40964
rect 5180 41186 5236 41188
rect 5180 41134 5182 41186
rect 5182 41134 5234 41186
rect 5234 41134 5236 41186
rect 5180 41132 5236 41134
rect 5292 41020 5348 41076
rect 5068 40908 5124 40964
rect 5292 40348 5348 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5068 39730 5124 39732
rect 5068 39678 5070 39730
rect 5070 39678 5122 39730
rect 5122 39678 5124 39730
rect 5068 39676 5124 39678
rect 4172 38668 4228 38724
rect 6076 42476 6132 42532
rect 5516 41186 5572 41188
rect 5516 41134 5518 41186
rect 5518 41134 5570 41186
rect 5570 41134 5572 41186
rect 5516 41132 5572 41134
rect 5852 41074 5908 41076
rect 5852 41022 5854 41074
rect 5854 41022 5906 41074
rect 5906 41022 5908 41074
rect 5852 41020 5908 41022
rect 5740 40962 5796 40964
rect 5740 40910 5742 40962
rect 5742 40910 5794 40962
rect 5794 40910 5796 40962
rect 5740 40908 5796 40910
rect 5404 39676 5460 39732
rect 7644 59442 7700 59444
rect 7644 59390 7646 59442
rect 7646 59390 7698 59442
rect 7698 59390 7700 59442
rect 7644 59388 7700 59390
rect 7532 59330 7588 59332
rect 7532 59278 7534 59330
rect 7534 59278 7586 59330
rect 7586 59278 7588 59330
rect 7532 59276 7588 59278
rect 10556 62412 10612 62468
rect 9548 62300 9604 62356
rect 10220 62354 10276 62356
rect 10220 62302 10222 62354
rect 10222 62302 10274 62354
rect 10274 62302 10276 62354
rect 10220 62300 10276 62302
rect 10892 62466 10948 62468
rect 10892 62414 10894 62466
rect 10894 62414 10946 62466
rect 10946 62414 10948 62466
rect 10892 62412 10948 62414
rect 12796 64818 12852 64820
rect 12796 64766 12798 64818
rect 12798 64766 12850 64818
rect 12850 64766 12852 64818
rect 12796 64764 12852 64766
rect 12684 64652 12740 64708
rect 12572 64594 12628 64596
rect 12572 64542 12574 64594
rect 12574 64542 12626 64594
rect 12626 64542 12628 64594
rect 12572 64540 12628 64542
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 20188 65490 20244 65492
rect 20188 65438 20190 65490
rect 20190 65438 20242 65490
rect 20242 65438 20244 65490
rect 20188 65436 20244 65438
rect 17612 65324 17668 65380
rect 13580 64706 13636 64708
rect 13580 64654 13582 64706
rect 13582 64654 13634 64706
rect 13634 64654 13636 64706
rect 13580 64652 13636 64654
rect 12236 63868 12292 63924
rect 12572 64092 12628 64148
rect 11900 62300 11956 62356
rect 10220 60732 10276 60788
rect 9100 60002 9156 60004
rect 9100 59950 9102 60002
rect 9102 59950 9154 60002
rect 9154 59950 9156 60002
rect 9100 59948 9156 59950
rect 8428 59724 8484 59780
rect 8204 59330 8260 59332
rect 8204 59278 8206 59330
rect 8206 59278 8258 59330
rect 8258 59278 8260 59330
rect 8204 59276 8260 59278
rect 11788 61628 11844 61684
rect 11004 60898 11060 60900
rect 11004 60846 11006 60898
rect 11006 60846 11058 60898
rect 11058 60846 11060 60898
rect 11004 60844 11060 60846
rect 10780 60786 10836 60788
rect 10780 60734 10782 60786
rect 10782 60734 10834 60786
rect 10834 60734 10836 60786
rect 10780 60732 10836 60734
rect 10556 60060 10612 60116
rect 12236 61682 12292 61684
rect 12236 61630 12238 61682
rect 12238 61630 12290 61682
rect 12290 61630 12292 61682
rect 12236 61628 12292 61630
rect 13804 64092 13860 64148
rect 12796 63980 12852 64036
rect 13692 64034 13748 64036
rect 13692 63982 13694 64034
rect 13694 63982 13746 64034
rect 13746 63982 13748 64034
rect 13692 63980 13748 63982
rect 14140 64034 14196 64036
rect 14140 63982 14142 64034
rect 14142 63982 14194 64034
rect 14194 63982 14196 64034
rect 14140 63980 14196 63982
rect 12908 63868 12964 63924
rect 14252 63922 14308 63924
rect 14252 63870 14254 63922
rect 14254 63870 14306 63922
rect 14306 63870 14308 63922
rect 14252 63868 14308 63870
rect 13132 63084 13188 63140
rect 13580 62300 13636 62356
rect 15484 63138 15540 63140
rect 15484 63086 15486 63138
rect 15486 63086 15538 63138
rect 15538 63086 15540 63138
rect 15484 63084 15540 63086
rect 16828 64706 16884 64708
rect 16828 64654 16830 64706
rect 16830 64654 16882 64706
rect 16882 64654 16884 64706
rect 16828 64652 16884 64654
rect 19516 65378 19572 65380
rect 19516 65326 19518 65378
rect 19518 65326 19570 65378
rect 19570 65326 19572 65378
rect 19516 65324 19572 65326
rect 17948 64706 18004 64708
rect 17948 64654 17950 64706
rect 17950 64654 18002 64706
rect 18002 64654 18004 64706
rect 17948 64652 18004 64654
rect 20860 65436 20916 65492
rect 20188 64652 20244 64708
rect 16716 63868 16772 63924
rect 16492 62972 16548 63028
rect 16268 62860 16324 62916
rect 17612 63922 17668 63924
rect 17612 63870 17614 63922
rect 17614 63870 17666 63922
rect 17666 63870 17668 63922
rect 17612 63868 17668 63870
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 20860 64428 20916 64484
rect 17276 63084 17332 63140
rect 17612 63026 17668 63028
rect 17612 62974 17614 63026
rect 17614 62974 17666 63026
rect 17666 62974 17668 63026
rect 17612 62972 17668 62974
rect 17388 62914 17444 62916
rect 17388 62862 17390 62914
rect 17390 62862 17442 62914
rect 17442 62862 17444 62914
rect 17388 62860 17444 62862
rect 17948 62860 18004 62916
rect 12684 61628 12740 61684
rect 15596 61628 15652 61684
rect 13244 60898 13300 60900
rect 13244 60846 13246 60898
rect 13246 60846 13298 60898
rect 13298 60846 13300 60898
rect 13244 60844 13300 60846
rect 13356 60786 13412 60788
rect 13356 60734 13358 60786
rect 13358 60734 13410 60786
rect 13410 60734 13412 60786
rect 13356 60732 13412 60734
rect 12572 60508 12628 60564
rect 13804 60508 13860 60564
rect 11788 59948 11844 60004
rect 11340 59724 11396 59780
rect 12796 60114 12852 60116
rect 12796 60062 12798 60114
rect 12798 60062 12850 60114
rect 12850 60062 12852 60114
rect 12796 60060 12852 60062
rect 12460 60002 12516 60004
rect 12460 59950 12462 60002
rect 12462 59950 12514 60002
rect 12514 59950 12516 60002
rect 12460 59948 12516 59950
rect 11004 58268 11060 58324
rect 8428 57596 8484 57652
rect 8204 56252 8260 56308
rect 8316 56194 8372 56196
rect 8316 56142 8318 56194
rect 8318 56142 8370 56194
rect 8370 56142 8372 56194
rect 8316 56140 8372 56142
rect 9436 57650 9492 57652
rect 9436 57598 9438 57650
rect 9438 57598 9490 57650
rect 9490 57598 9492 57650
rect 9436 57596 9492 57598
rect 10108 57650 10164 57652
rect 10108 57598 10110 57650
rect 10110 57598 10162 57650
rect 10162 57598 10164 57650
rect 10108 57596 10164 57598
rect 9996 57036 10052 57092
rect 9772 56700 9828 56756
rect 8764 56306 8820 56308
rect 8764 56254 8766 56306
rect 8766 56254 8818 56306
rect 8818 56254 8820 56306
rect 8764 56252 8820 56254
rect 9884 56252 9940 56308
rect 8988 56140 9044 56196
rect 7196 55580 7252 55636
rect 6860 54348 6916 54404
rect 7196 53506 7252 53508
rect 7196 53454 7198 53506
rect 7198 53454 7250 53506
rect 7250 53454 7252 53506
rect 7196 53452 7252 53454
rect 7420 53452 7476 53508
rect 8092 53506 8148 53508
rect 8092 53454 8094 53506
rect 8094 53454 8146 53506
rect 8146 53454 8148 53506
rect 8092 53452 8148 53454
rect 7644 53116 7700 53172
rect 8652 53452 8708 53508
rect 7308 52780 7364 52836
rect 6860 52220 6916 52276
rect 8540 53170 8596 53172
rect 8540 53118 8542 53170
rect 8542 53118 8594 53170
rect 8594 53118 8596 53170
rect 8540 53116 8596 53118
rect 8428 52780 8484 52836
rect 8204 52444 8260 52500
rect 7980 51996 8036 52052
rect 8652 52444 8708 52500
rect 10444 57036 10500 57092
rect 10668 57650 10724 57652
rect 10668 57598 10670 57650
rect 10670 57598 10722 57650
rect 10722 57598 10724 57650
rect 10668 57596 10724 57598
rect 10780 57036 10836 57092
rect 10332 55468 10388 55524
rect 11788 58268 11844 58324
rect 12236 58828 12292 58884
rect 11900 57484 11956 57540
rect 11228 56700 11284 56756
rect 11004 55468 11060 55524
rect 11788 55468 11844 55524
rect 11340 55298 11396 55300
rect 11340 55246 11342 55298
rect 11342 55246 11394 55298
rect 11394 55246 11396 55298
rect 11340 55244 11396 55246
rect 8764 52050 8820 52052
rect 8764 51998 8766 52050
rect 8766 51998 8818 52050
rect 8818 51998 8820 52050
rect 8764 51996 8820 51998
rect 8988 49868 9044 49924
rect 8876 49810 8932 49812
rect 8876 49758 8878 49810
rect 8878 49758 8930 49810
rect 8930 49758 8932 49810
rect 8876 49756 8932 49758
rect 8540 49084 8596 49140
rect 6748 48914 6804 48916
rect 6748 48862 6750 48914
rect 6750 48862 6802 48914
rect 6802 48862 6804 48914
rect 6748 48860 6804 48862
rect 8428 48748 8484 48804
rect 8316 48466 8372 48468
rect 8316 48414 8318 48466
rect 8318 48414 8370 48466
rect 8370 48414 8372 48466
rect 8316 48412 8372 48414
rect 8092 48354 8148 48356
rect 8092 48302 8094 48354
rect 8094 48302 8146 48354
rect 8146 48302 8148 48354
rect 8092 48300 8148 48302
rect 9100 49084 9156 49140
rect 10668 52834 10724 52836
rect 10668 52782 10670 52834
rect 10670 52782 10722 52834
rect 10722 52782 10724 52834
rect 10668 52780 10724 52782
rect 10108 52444 10164 52500
rect 10220 52668 10276 52724
rect 10780 52162 10836 52164
rect 10780 52110 10782 52162
rect 10782 52110 10834 52162
rect 10834 52110 10836 52162
rect 10780 52108 10836 52110
rect 11452 52444 11508 52500
rect 9324 49756 9380 49812
rect 9324 48914 9380 48916
rect 9324 48862 9326 48914
rect 9326 48862 9378 48914
rect 9378 48862 9380 48914
rect 9324 48860 9380 48862
rect 10220 49922 10276 49924
rect 10220 49870 10222 49922
rect 10222 49870 10274 49922
rect 10274 49870 10276 49922
rect 10220 49868 10276 49870
rect 10332 49810 10388 49812
rect 10332 49758 10334 49810
rect 10334 49758 10386 49810
rect 10386 49758 10388 49810
rect 10332 49756 10388 49758
rect 9212 48300 9268 48356
rect 9660 48748 9716 48804
rect 10108 48972 10164 49028
rect 9548 48412 9604 48468
rect 9548 47628 9604 47684
rect 9660 47404 9716 47460
rect 7532 45164 7588 45220
rect 8204 45164 8260 45220
rect 8764 45724 8820 45780
rect 9996 46002 10052 46004
rect 9996 45950 9998 46002
rect 9998 45950 10050 46002
rect 10050 45950 10052 46002
rect 9996 45948 10052 45950
rect 8876 45276 8932 45332
rect 9436 45388 9492 45444
rect 9996 45724 10052 45780
rect 9772 45330 9828 45332
rect 9772 45278 9774 45330
rect 9774 45278 9826 45330
rect 9826 45278 9828 45330
rect 9772 45276 9828 45278
rect 9436 45052 9492 45108
rect 10108 45164 10164 45220
rect 8764 42754 8820 42756
rect 8764 42702 8766 42754
rect 8766 42702 8818 42754
rect 8818 42702 8820 42754
rect 8764 42700 8820 42702
rect 8316 42588 8372 42644
rect 8204 41916 8260 41972
rect 8204 41132 8260 41188
rect 5852 38780 5908 38836
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4060 38050 4116 38052
rect 4060 37998 4062 38050
rect 4062 37998 4114 38050
rect 4114 37998 4116 38050
rect 4060 37996 4116 37998
rect 2716 37436 2772 37492
rect 3612 37490 3668 37492
rect 3612 37438 3614 37490
rect 3614 37438 3666 37490
rect 3666 37438 3668 37490
rect 3612 37436 3668 37438
rect 3052 37378 3108 37380
rect 3052 37326 3054 37378
rect 3054 37326 3106 37378
rect 3106 37326 3108 37378
rect 3052 37324 3108 37326
rect 3948 37324 4004 37380
rect 3164 37266 3220 37268
rect 3164 37214 3166 37266
rect 3166 37214 3218 37266
rect 3218 37214 3220 37266
rect 3164 37212 3220 37214
rect 3724 37266 3780 37268
rect 3724 37214 3726 37266
rect 3726 37214 3778 37266
rect 3778 37214 3780 37266
rect 3724 37212 3780 37214
rect 4620 37266 4676 37268
rect 4620 37214 4622 37266
rect 4622 37214 4674 37266
rect 4674 37214 4676 37266
rect 4620 37212 4676 37214
rect 6636 38834 6692 38836
rect 6636 38782 6638 38834
rect 6638 38782 6690 38834
rect 6690 38782 6692 38834
rect 6636 38780 6692 38782
rect 6412 38556 6468 38612
rect 7868 39004 7924 39060
rect 9100 42642 9156 42644
rect 9100 42590 9102 42642
rect 9102 42590 9154 42642
rect 9154 42590 9156 42642
rect 9100 42588 9156 42590
rect 8988 42530 9044 42532
rect 8988 42478 8990 42530
rect 8990 42478 9042 42530
rect 9042 42478 9044 42530
rect 8988 42476 9044 42478
rect 8876 42252 8932 42308
rect 8764 41916 8820 41972
rect 9660 42252 9716 42308
rect 9884 42140 9940 42196
rect 9548 41244 9604 41300
rect 9660 41916 9716 41972
rect 8652 41186 8708 41188
rect 8652 41134 8654 41186
rect 8654 41134 8706 41186
rect 8706 41134 8708 41186
rect 8652 41132 8708 41134
rect 9996 41298 10052 41300
rect 9996 41246 9998 41298
rect 9998 41246 10050 41298
rect 10050 41246 10052 41298
rect 9996 41244 10052 41246
rect 10108 41132 10164 41188
rect 7868 38780 7924 38836
rect 7532 38722 7588 38724
rect 7532 38670 7534 38722
rect 7534 38670 7586 38722
rect 7586 38670 7588 38722
rect 7532 38668 7588 38670
rect 7420 38556 7476 38612
rect 7084 38444 7140 38500
rect 5180 37212 5236 37268
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 7980 38556 8036 38612
rect 9884 38274 9940 38276
rect 9884 38222 9886 38274
rect 9886 38222 9938 38274
rect 9938 38222 9940 38274
rect 9884 38220 9940 38222
rect 8428 37324 8484 37380
rect 7868 37266 7924 37268
rect 7868 37214 7870 37266
rect 7870 37214 7922 37266
rect 7922 37214 7924 37266
rect 7868 37212 7924 37214
rect 8540 37212 8596 37268
rect 8764 37378 8820 37380
rect 8764 37326 8766 37378
rect 8766 37326 8818 37378
rect 8818 37326 8820 37378
rect 8764 37324 8820 37326
rect 8764 37154 8820 37156
rect 8764 37102 8766 37154
rect 8766 37102 8818 37154
rect 8818 37102 8820 37154
rect 8764 37100 8820 37102
rect 9100 36988 9156 37044
rect 8764 36540 8820 36596
rect 2268 35586 2324 35588
rect 2268 35534 2270 35586
rect 2270 35534 2322 35586
rect 2322 35534 2324 35586
rect 2268 35532 2324 35534
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 7868 34914 7924 34916
rect 7868 34862 7870 34914
rect 7870 34862 7922 34914
rect 7922 34862 7924 34914
rect 7868 34860 7924 34862
rect 8652 35644 8708 35700
rect 8764 35308 8820 35364
rect 8876 36316 8932 36372
rect 8428 34914 8484 34916
rect 8428 34862 8430 34914
rect 8430 34862 8482 34914
rect 8482 34862 8484 34914
rect 8428 34860 8484 34862
rect 5852 33964 5908 34020
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 5068 29314 5124 29316
rect 5068 29262 5070 29314
rect 5070 29262 5122 29314
rect 5122 29262 5124 29314
rect 5068 29260 5124 29262
rect 5516 28364 5572 28420
rect 4844 27858 4900 27860
rect 4844 27806 4846 27858
rect 4846 27806 4898 27858
rect 4898 27806 4900 27858
rect 4844 27804 4900 27806
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2268 26460 2324 26516
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 7980 31836 8036 31892
rect 8540 32620 8596 32676
rect 8764 34188 8820 34244
rect 9324 37212 9380 37268
rect 9436 37100 9492 37156
rect 9884 37378 9940 37380
rect 9884 37326 9886 37378
rect 9886 37326 9938 37378
rect 9938 37326 9940 37378
rect 9884 37324 9940 37326
rect 9548 36988 9604 37044
rect 10220 36988 10276 37044
rect 9772 36540 9828 36596
rect 9436 35308 9492 35364
rect 9548 34914 9604 34916
rect 9548 34862 9550 34914
rect 9550 34862 9602 34914
rect 9602 34862 9604 34914
rect 9548 34860 9604 34862
rect 8764 32396 8820 32452
rect 8092 31666 8148 31668
rect 8092 31614 8094 31666
rect 8094 31614 8146 31666
rect 8146 31614 8148 31666
rect 8092 31612 8148 31614
rect 7644 30994 7700 30996
rect 7644 30942 7646 30994
rect 7646 30942 7698 30994
rect 7698 30942 7700 30994
rect 7644 30940 7700 30942
rect 8204 30380 8260 30436
rect 8092 30268 8148 30324
rect 8540 30994 8596 30996
rect 8540 30942 8542 30994
rect 8542 30942 8594 30994
rect 8594 30942 8596 30994
rect 8540 30940 8596 30942
rect 8428 30268 8484 30324
rect 8876 31836 8932 31892
rect 8988 31666 9044 31668
rect 8988 31614 8990 31666
rect 8990 31614 9042 31666
rect 9042 31614 9044 31666
rect 8988 31612 9044 31614
rect 8876 30994 8932 30996
rect 8876 30942 8878 30994
rect 8878 30942 8930 30994
rect 8930 30942 8932 30994
rect 8876 30940 8932 30942
rect 8988 30380 9044 30436
rect 9324 30716 9380 30772
rect 9212 30322 9268 30324
rect 9212 30270 9214 30322
rect 9214 30270 9266 30322
rect 9266 30270 9268 30322
rect 9212 30268 9268 30270
rect 6076 27804 6132 27860
rect 7196 27804 7252 27860
rect 8316 28028 8372 28084
rect 8092 27858 8148 27860
rect 8092 27806 8094 27858
rect 8094 27806 8146 27858
rect 8146 27806 8148 27858
rect 8092 27804 8148 27806
rect 7644 27746 7700 27748
rect 7644 27694 7646 27746
rect 7646 27694 7698 27746
rect 7698 27694 7700 27746
rect 7644 27692 7700 27694
rect 8988 29596 9044 29652
rect 9884 36092 9940 36148
rect 10780 49980 10836 50036
rect 10556 48354 10612 48356
rect 10556 48302 10558 48354
rect 10558 48302 10610 48354
rect 10610 48302 10612 48354
rect 10556 48300 10612 48302
rect 10556 46732 10612 46788
rect 10556 45948 10612 46004
rect 10556 42140 10612 42196
rect 10780 38668 10836 38724
rect 11788 51548 11844 51604
rect 11676 50706 11732 50708
rect 11676 50654 11678 50706
rect 11678 50654 11730 50706
rect 11730 50654 11732 50706
rect 11676 50652 11732 50654
rect 11116 49980 11172 50036
rect 11116 48076 11172 48132
rect 11116 47682 11172 47684
rect 11116 47630 11118 47682
rect 11118 47630 11170 47682
rect 11170 47630 11172 47682
rect 11116 47628 11172 47630
rect 11340 48300 11396 48356
rect 11116 47458 11172 47460
rect 11116 47406 11118 47458
rect 11118 47406 11170 47458
rect 11170 47406 11172 47458
rect 11116 47404 11172 47406
rect 11788 47404 11844 47460
rect 11676 45276 11732 45332
rect 11788 47180 11844 47236
rect 14140 60002 14196 60004
rect 14140 59950 14142 60002
rect 14142 59950 14194 60002
rect 14194 59950 14196 60002
rect 14140 59948 14196 59950
rect 15148 59948 15204 60004
rect 12796 59724 12852 59780
rect 12796 59106 12852 59108
rect 12796 59054 12798 59106
rect 12798 59054 12850 59106
rect 12850 59054 12852 59106
rect 12796 59052 12852 59054
rect 15036 59724 15092 59780
rect 13804 58434 13860 58436
rect 13804 58382 13806 58434
rect 13806 58382 13858 58434
rect 13858 58382 13860 58434
rect 13804 58380 13860 58382
rect 12460 57484 12516 57540
rect 13356 57538 13412 57540
rect 13356 57486 13358 57538
rect 13358 57486 13410 57538
rect 13410 57486 13412 57538
rect 13356 57484 13412 57486
rect 13916 57484 13972 57540
rect 12236 57090 12292 57092
rect 12236 57038 12238 57090
rect 12238 57038 12290 57090
rect 12290 57038 12292 57090
rect 12236 57036 12292 57038
rect 12012 56754 12068 56756
rect 12012 56702 12014 56754
rect 12014 56702 12066 56754
rect 12066 56702 12068 56754
rect 12012 56700 12068 56702
rect 13692 56700 13748 56756
rect 12572 56642 12628 56644
rect 12572 56590 12574 56642
rect 12574 56590 12626 56642
rect 12626 56590 12628 56642
rect 12572 56588 12628 56590
rect 12908 56252 12964 56308
rect 14364 58828 14420 58884
rect 14924 58380 14980 58436
rect 14252 56754 14308 56756
rect 14252 56702 14254 56754
rect 14254 56702 14306 56754
rect 14306 56702 14308 56754
rect 14252 56700 14308 56702
rect 13916 56588 13972 56644
rect 13356 56194 13412 56196
rect 13356 56142 13358 56194
rect 13358 56142 13410 56194
rect 13410 56142 13412 56194
rect 13356 56140 13412 56142
rect 13020 55468 13076 55524
rect 12684 55074 12740 55076
rect 12684 55022 12686 55074
rect 12686 55022 12738 55074
rect 12738 55022 12740 55074
rect 12684 55020 12740 55022
rect 12572 54460 12628 54516
rect 12908 53004 12964 53060
rect 12348 52780 12404 52836
rect 12796 52108 12852 52164
rect 12236 50652 12292 50708
rect 13132 55356 13188 55412
rect 14028 56194 14084 56196
rect 14028 56142 14030 56194
rect 14030 56142 14082 56194
rect 14082 56142 14084 56194
rect 14028 56140 14084 56142
rect 14252 56082 14308 56084
rect 14252 56030 14254 56082
rect 14254 56030 14306 56082
rect 14306 56030 14308 56082
rect 14252 56028 14308 56030
rect 14028 55356 14084 55412
rect 15708 60732 15764 60788
rect 15596 59948 15652 60004
rect 16268 60844 16324 60900
rect 16156 59890 16212 59892
rect 16156 59838 16158 59890
rect 16158 59838 16210 59890
rect 16210 59838 16212 59890
rect 16156 59836 16212 59838
rect 17500 60898 17556 60900
rect 17500 60846 17502 60898
rect 17502 60846 17554 60898
rect 17554 60846 17556 60898
rect 17500 60844 17556 60846
rect 18172 62300 18228 62356
rect 17612 60226 17668 60228
rect 17612 60174 17614 60226
rect 17614 60174 17666 60226
rect 17666 60174 17668 60226
rect 17612 60172 17668 60174
rect 16940 59724 16996 59780
rect 15932 59164 15988 59220
rect 14924 57708 14980 57764
rect 16380 59218 16436 59220
rect 16380 59166 16382 59218
rect 16382 59166 16434 59218
rect 16434 59166 16436 59218
rect 16380 59164 16436 59166
rect 16492 59052 16548 59108
rect 16380 58434 16436 58436
rect 16380 58382 16382 58434
rect 16382 58382 16434 58434
rect 16434 58382 16436 58434
rect 16380 58380 16436 58382
rect 15484 57708 15540 57764
rect 15148 56754 15204 56756
rect 15148 56702 15150 56754
rect 15150 56702 15202 56754
rect 15202 56702 15204 56754
rect 15148 56700 15204 56702
rect 14588 56588 14644 56644
rect 14588 56306 14644 56308
rect 14588 56254 14590 56306
rect 14590 56254 14642 56306
rect 14642 56254 14644 56306
rect 14588 56252 14644 56254
rect 15148 56082 15204 56084
rect 15148 56030 15150 56082
rect 15150 56030 15202 56082
rect 15202 56030 15204 56082
rect 15148 56028 15204 56030
rect 14924 55356 14980 55412
rect 13468 55244 13524 55300
rect 14476 55298 14532 55300
rect 14476 55246 14478 55298
rect 14478 55246 14530 55298
rect 14530 55246 14532 55298
rect 14476 55244 14532 55246
rect 13580 55074 13636 55076
rect 13580 55022 13582 55074
rect 13582 55022 13634 55074
rect 13634 55022 13636 55074
rect 13580 55020 13636 55022
rect 12348 50034 12404 50036
rect 12348 49982 12350 50034
rect 12350 49982 12402 50034
rect 12402 49982 12404 50034
rect 12348 49980 12404 49982
rect 12684 49810 12740 49812
rect 12684 49758 12686 49810
rect 12686 49758 12738 49810
rect 12738 49758 12740 49810
rect 12684 49756 12740 49758
rect 12684 47234 12740 47236
rect 12684 47182 12686 47234
rect 12686 47182 12738 47234
rect 12738 47182 12740 47234
rect 12684 47180 12740 47182
rect 12348 46844 12404 46900
rect 13356 52108 13412 52164
rect 13244 51602 13300 51604
rect 13244 51550 13246 51602
rect 13246 51550 13298 51602
rect 13298 51550 13300 51602
rect 13244 51548 13300 51550
rect 13468 51548 13524 51604
rect 13244 49810 13300 49812
rect 13244 49758 13246 49810
rect 13246 49758 13298 49810
rect 13298 49758 13300 49810
rect 13244 49756 13300 49758
rect 12908 48076 12964 48132
rect 12796 46786 12852 46788
rect 12796 46734 12798 46786
rect 12798 46734 12850 46786
rect 12850 46734 12852 46786
rect 12796 46732 12852 46734
rect 13020 47180 13076 47236
rect 12796 45388 12852 45444
rect 12124 43932 12180 43988
rect 11788 42700 11844 42756
rect 11788 41244 11844 41300
rect 11004 41020 11060 41076
rect 12572 44044 12628 44100
rect 12348 41074 12404 41076
rect 12348 41022 12350 41074
rect 12350 41022 12402 41074
rect 12402 41022 12404 41074
rect 12348 41020 12404 41022
rect 11004 40348 11060 40404
rect 12460 40908 12516 40964
rect 11452 38834 11508 38836
rect 11452 38782 11454 38834
rect 11454 38782 11506 38834
rect 11506 38782 11508 38834
rect 11452 38780 11508 38782
rect 11676 38722 11732 38724
rect 11676 38670 11678 38722
rect 11678 38670 11730 38722
rect 11730 38670 11732 38722
rect 11676 38668 11732 38670
rect 11788 38332 11844 38388
rect 12684 43932 12740 43988
rect 12012 38946 12068 38948
rect 12012 38894 12014 38946
rect 12014 38894 12066 38946
rect 12066 38894 12068 38946
rect 12012 38892 12068 38894
rect 11900 38220 11956 38276
rect 11116 37996 11172 38052
rect 10892 37324 10948 37380
rect 11340 37378 11396 37380
rect 11340 37326 11342 37378
rect 11342 37326 11394 37378
rect 11394 37326 11396 37378
rect 11340 37324 11396 37326
rect 10556 36988 10612 37044
rect 11004 36988 11060 37044
rect 10780 36258 10836 36260
rect 10780 36206 10782 36258
rect 10782 36206 10834 36258
rect 10834 36206 10836 36258
rect 10780 36204 10836 36206
rect 11004 36092 11060 36148
rect 9996 34914 10052 34916
rect 9996 34862 9998 34914
rect 9998 34862 10050 34914
rect 10050 34862 10052 34914
rect 9996 34860 10052 34862
rect 11340 35698 11396 35700
rect 11340 35646 11342 35698
rect 11342 35646 11394 35698
rect 11394 35646 11396 35698
rect 11340 35644 11396 35646
rect 11564 36370 11620 36372
rect 11564 36318 11566 36370
rect 11566 36318 11618 36370
rect 11618 36318 11620 36370
rect 11564 36316 11620 36318
rect 11900 36988 11956 37044
rect 12572 39394 12628 39396
rect 12572 39342 12574 39394
rect 12574 39342 12626 39394
rect 12626 39342 12628 39394
rect 12572 39340 12628 39342
rect 12236 38556 12292 38612
rect 12348 39004 12404 39060
rect 12572 38834 12628 38836
rect 12572 38782 12574 38834
rect 12574 38782 12626 38834
rect 12626 38782 12628 38834
rect 12572 38780 12628 38782
rect 12460 38668 12516 38724
rect 12572 38556 12628 38612
rect 13020 43036 13076 43092
rect 12796 40572 12852 40628
rect 12908 39564 12964 39620
rect 12908 38892 12964 38948
rect 13132 38780 13188 38836
rect 12460 37378 12516 37380
rect 12460 37326 12462 37378
rect 12462 37326 12514 37378
rect 12514 37326 12516 37378
rect 12460 37324 12516 37326
rect 11900 36316 11956 36372
rect 10556 34636 10612 34692
rect 9884 34130 9940 34132
rect 9884 34078 9886 34130
rect 9886 34078 9938 34130
rect 9938 34078 9940 34130
rect 9884 34076 9940 34078
rect 10556 33628 10612 33684
rect 10780 34242 10836 34244
rect 10780 34190 10782 34242
rect 10782 34190 10834 34242
rect 10834 34190 10836 34242
rect 10780 34188 10836 34190
rect 9884 32450 9940 32452
rect 9884 32398 9886 32450
rect 9886 32398 9938 32450
rect 9938 32398 9940 32450
rect 9884 32396 9940 32398
rect 9772 31612 9828 31668
rect 9772 30268 9828 30324
rect 10892 33292 10948 33348
rect 10220 30828 10276 30884
rect 9996 29372 10052 29428
rect 11116 34860 11172 34916
rect 12684 36258 12740 36260
rect 12684 36206 12686 36258
rect 12686 36206 12738 36258
rect 12738 36206 12740 36258
rect 12684 36204 12740 36206
rect 13356 46898 13412 46900
rect 13356 46846 13358 46898
rect 13358 46846 13410 46898
rect 13410 46846 13412 46898
rect 13356 46844 13412 46846
rect 13692 52108 13748 52164
rect 13804 51548 13860 51604
rect 14476 54514 14532 54516
rect 14476 54462 14478 54514
rect 14478 54462 14530 54514
rect 14530 54462 14532 54514
rect 14476 54460 14532 54462
rect 15372 54514 15428 54516
rect 15372 54462 15374 54514
rect 15374 54462 15426 54514
rect 15426 54462 15428 54514
rect 15372 54460 15428 54462
rect 14812 53058 14868 53060
rect 14812 53006 14814 53058
rect 14814 53006 14866 53058
rect 14866 53006 14868 53058
rect 14812 53004 14868 53006
rect 14924 52220 14980 52276
rect 14476 52162 14532 52164
rect 14476 52110 14478 52162
rect 14478 52110 14530 52162
rect 14530 52110 14532 52162
rect 14476 52108 14532 52110
rect 15260 52162 15316 52164
rect 15260 52110 15262 52162
rect 15262 52110 15314 52162
rect 15314 52110 15316 52162
rect 15260 52108 15316 52110
rect 14028 49980 14084 50036
rect 14252 49810 14308 49812
rect 14252 49758 14254 49810
rect 14254 49758 14306 49810
rect 14306 49758 14308 49810
rect 14252 49756 14308 49758
rect 14028 48242 14084 48244
rect 14028 48190 14030 48242
rect 14030 48190 14082 48242
rect 14082 48190 14084 48242
rect 14028 48188 14084 48190
rect 13804 48076 13860 48132
rect 14140 48130 14196 48132
rect 14140 48078 14142 48130
rect 14142 48078 14194 48130
rect 14194 48078 14196 48130
rect 14140 48076 14196 48078
rect 14700 49586 14756 49588
rect 14700 49534 14702 49586
rect 14702 49534 14754 49586
rect 14754 49534 14756 49586
rect 14700 49532 14756 49534
rect 13692 46956 13748 47012
rect 13580 45948 13636 46004
rect 13580 45388 13636 45444
rect 13468 44268 13524 44324
rect 13244 38332 13300 38388
rect 13468 41916 13524 41972
rect 10444 30716 10500 30772
rect 10332 29596 10388 29652
rect 11452 34636 11508 34692
rect 11676 33346 11732 33348
rect 11676 33294 11678 33346
rect 11678 33294 11730 33346
rect 11730 33294 11732 33346
rect 11676 33292 11732 33294
rect 11116 30716 11172 30772
rect 11004 30380 11060 30436
rect 10668 29708 10724 29764
rect 8652 27692 8708 27748
rect 9548 27692 9604 27748
rect 9660 27804 9716 27860
rect 9996 27746 10052 27748
rect 9996 27694 9998 27746
rect 9998 27694 10050 27746
rect 10050 27694 10052 27746
rect 9996 27692 10052 27694
rect 8876 26852 8932 26908
rect 8988 26124 9044 26180
rect 8876 25900 8932 25956
rect 8204 25394 8260 25396
rect 8204 25342 8206 25394
rect 8206 25342 8258 25394
rect 8258 25342 8260 25394
rect 8204 25340 8260 25342
rect 9548 26124 9604 26180
rect 9660 25900 9716 25956
rect 9436 25618 9492 25620
rect 9436 25566 9438 25618
rect 9438 25566 9490 25618
rect 9490 25566 9492 25618
rect 9436 25564 9492 25566
rect 8988 25340 9044 25396
rect 11116 30322 11172 30324
rect 11116 30270 11118 30322
rect 11118 30270 11170 30322
rect 11170 30270 11172 30322
rect 11116 30268 11172 30270
rect 12012 33628 12068 33684
rect 12684 34690 12740 34692
rect 12684 34638 12686 34690
rect 12686 34638 12738 34690
rect 12738 34638 12740 34690
rect 12684 34636 12740 34638
rect 14252 46620 14308 46676
rect 14476 46508 14532 46564
rect 16716 59442 16772 59444
rect 16716 59390 16718 59442
rect 16718 59390 16770 59442
rect 16770 59390 16772 59442
rect 16716 59388 16772 59390
rect 17612 59330 17668 59332
rect 17612 59278 17614 59330
rect 17614 59278 17666 59330
rect 17666 59278 17668 59330
rect 17612 59276 17668 59278
rect 18060 59836 18116 59892
rect 18172 60060 18228 60116
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 24892 66444 24948 66500
rect 26124 66498 26180 66500
rect 26124 66446 26126 66498
rect 26126 66446 26178 66498
rect 26178 66446 26180 66498
rect 26124 66444 26180 66446
rect 21420 64482 21476 64484
rect 21420 64430 21422 64482
rect 21422 64430 21474 64482
rect 21474 64430 21476 64482
rect 21420 64428 21476 64430
rect 22540 64876 22596 64932
rect 21868 64428 21924 64484
rect 23548 64930 23604 64932
rect 23548 64878 23550 64930
rect 23550 64878 23602 64930
rect 23602 64878 23604 64930
rect 23548 64876 23604 64878
rect 23212 64482 23268 64484
rect 23212 64430 23214 64482
rect 23214 64430 23266 64482
rect 23266 64430 23268 64482
rect 23212 64428 23268 64430
rect 21084 63308 21140 63364
rect 22316 63362 22372 63364
rect 22316 63310 22318 63362
rect 22318 63310 22370 63362
rect 22370 63310 22372 63362
rect 22316 63308 22372 63310
rect 18956 62466 19012 62468
rect 18956 62414 18958 62466
rect 18958 62414 19010 62466
rect 19010 62414 19012 62466
rect 18956 62412 19012 62414
rect 20412 62412 20468 62468
rect 19516 62354 19572 62356
rect 19516 62302 19518 62354
rect 19518 62302 19570 62354
rect 19570 62302 19572 62354
rect 19516 62300 19572 62302
rect 20860 62466 20916 62468
rect 20860 62414 20862 62466
rect 20862 62414 20914 62466
rect 20914 62414 20916 62466
rect 20860 62412 20916 62414
rect 18844 60284 18900 60340
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 20188 60284 20244 60340
rect 19852 60060 19908 60116
rect 18172 59388 18228 59444
rect 18060 59276 18116 59332
rect 18060 59106 18116 59108
rect 18060 59054 18062 59106
rect 18062 59054 18114 59106
rect 18114 59054 18116 59106
rect 18060 59052 18116 59054
rect 16604 58268 16660 58324
rect 15932 55858 15988 55860
rect 15932 55806 15934 55858
rect 15934 55806 15986 55858
rect 15986 55806 15988 55858
rect 15932 55804 15988 55806
rect 16044 54402 16100 54404
rect 16044 54350 16046 54402
rect 16046 54350 16098 54402
rect 16098 54350 16100 54402
rect 16044 54348 16100 54350
rect 16492 52386 16548 52388
rect 16492 52334 16494 52386
rect 16494 52334 16546 52386
rect 16546 52334 16548 52386
rect 16492 52332 16548 52334
rect 15932 52162 15988 52164
rect 15932 52110 15934 52162
rect 15934 52110 15986 52162
rect 15986 52110 15988 52162
rect 15932 52108 15988 52110
rect 15596 49532 15652 49588
rect 15484 48242 15540 48244
rect 15484 48190 15486 48242
rect 15486 48190 15538 48242
rect 15538 48190 15540 48242
rect 15484 48188 15540 48190
rect 14924 47404 14980 47460
rect 15036 47346 15092 47348
rect 15036 47294 15038 47346
rect 15038 47294 15090 47346
rect 15090 47294 15092 47346
rect 15036 47292 15092 47294
rect 14812 46844 14868 46900
rect 14700 46674 14756 46676
rect 14700 46622 14702 46674
rect 14702 46622 14754 46674
rect 14754 46622 14756 46674
rect 14700 46620 14756 46622
rect 14028 45500 14084 45556
rect 14924 46562 14980 46564
rect 14924 46510 14926 46562
rect 14926 46510 14978 46562
rect 14978 46510 14980 46562
rect 14924 46508 14980 46510
rect 14812 45778 14868 45780
rect 14812 45726 14814 45778
rect 14814 45726 14866 45778
rect 14866 45726 14868 45778
rect 14812 45724 14868 45726
rect 14812 45500 14868 45556
rect 13804 44098 13860 44100
rect 13804 44046 13806 44098
rect 13806 44046 13858 44098
rect 13858 44046 13860 44098
rect 13804 44044 13860 44046
rect 13916 43036 13972 43092
rect 13804 41468 13860 41524
rect 14140 41970 14196 41972
rect 14140 41918 14142 41970
rect 14142 41918 14194 41970
rect 14194 41918 14196 41970
rect 14140 41916 14196 41918
rect 14476 41970 14532 41972
rect 14476 41918 14478 41970
rect 14478 41918 14530 41970
rect 14530 41918 14532 41970
rect 14476 41916 14532 41918
rect 13692 40962 13748 40964
rect 13692 40910 13694 40962
rect 13694 40910 13746 40962
rect 13746 40910 13748 40962
rect 13692 40908 13748 40910
rect 13916 41074 13972 41076
rect 13916 41022 13918 41074
rect 13918 41022 13970 41074
rect 13970 41022 13972 41074
rect 13916 41020 13972 41022
rect 15932 48188 15988 48244
rect 15372 47404 15428 47460
rect 15708 47346 15764 47348
rect 15708 47294 15710 47346
rect 15710 47294 15762 47346
rect 15762 47294 15764 47346
rect 15708 47292 15764 47294
rect 15372 46562 15428 46564
rect 15372 46510 15374 46562
rect 15374 46510 15426 46562
rect 15426 46510 15428 46562
rect 15372 46508 15428 46510
rect 15484 45778 15540 45780
rect 15484 45726 15486 45778
rect 15486 45726 15538 45778
rect 15538 45726 15540 45778
rect 15484 45724 15540 45726
rect 15148 45052 15204 45108
rect 15820 45890 15876 45892
rect 15820 45838 15822 45890
rect 15822 45838 15874 45890
rect 15874 45838 15876 45890
rect 15820 45836 15876 45838
rect 15820 45106 15876 45108
rect 15820 45054 15822 45106
rect 15822 45054 15874 45106
rect 15874 45054 15876 45106
rect 15820 45052 15876 45054
rect 15596 44380 15652 44436
rect 15484 44322 15540 44324
rect 15484 44270 15486 44322
rect 15486 44270 15538 44322
rect 15538 44270 15540 44322
rect 15484 44268 15540 44270
rect 15820 44268 15876 44324
rect 14924 42812 14980 42868
rect 14812 41804 14868 41860
rect 14700 41132 14756 41188
rect 14028 40626 14084 40628
rect 14028 40574 14030 40626
rect 14030 40574 14082 40626
rect 14082 40574 14084 40626
rect 14028 40572 14084 40574
rect 13804 40124 13860 40180
rect 14140 39618 14196 39620
rect 14140 39566 14142 39618
rect 14142 39566 14194 39618
rect 14194 39566 14196 39618
rect 14140 39564 14196 39566
rect 14028 38050 14084 38052
rect 14028 37998 14030 38050
rect 14030 37998 14082 38050
rect 14082 37998 14084 38050
rect 14028 37996 14084 37998
rect 13468 34914 13524 34916
rect 13468 34862 13470 34914
rect 13470 34862 13522 34914
rect 13522 34862 13524 34914
rect 13468 34860 13524 34862
rect 12908 34802 12964 34804
rect 12908 34750 12910 34802
rect 12910 34750 12962 34802
rect 12962 34750 12964 34802
rect 12908 34748 12964 34750
rect 13132 33852 13188 33908
rect 12796 33068 12852 33124
rect 12460 32620 12516 32676
rect 13468 33122 13524 33124
rect 13468 33070 13470 33122
rect 13470 33070 13522 33122
rect 13522 33070 13524 33122
rect 13468 33068 13524 33070
rect 11788 30940 11844 30996
rect 11452 30828 11508 30884
rect 11228 28812 11284 28868
rect 11004 28252 11060 28308
rect 11900 30156 11956 30212
rect 11452 28082 11508 28084
rect 11452 28030 11454 28082
rect 11454 28030 11506 28082
rect 11506 28030 11508 28082
rect 11452 28028 11508 28030
rect 11788 28082 11844 28084
rect 11788 28030 11790 28082
rect 11790 28030 11842 28082
rect 11842 28030 11844 28082
rect 11788 28028 11844 28030
rect 10892 26908 10948 26964
rect 12572 31666 12628 31668
rect 12572 31614 12574 31666
rect 12574 31614 12626 31666
rect 12626 31614 12628 31666
rect 12572 31612 12628 31614
rect 13020 31836 13076 31892
rect 12908 30994 12964 30996
rect 12908 30942 12910 30994
rect 12910 30942 12962 30994
rect 12962 30942 12964 30994
rect 12908 30940 12964 30942
rect 12684 30882 12740 30884
rect 12684 30830 12686 30882
rect 12686 30830 12738 30882
rect 12738 30830 12740 30882
rect 12684 30828 12740 30830
rect 12012 29426 12068 29428
rect 12012 29374 12014 29426
rect 12014 29374 12066 29426
rect 12066 29374 12068 29426
rect 12012 29372 12068 29374
rect 12012 28866 12068 28868
rect 12012 28814 12014 28866
rect 12014 28814 12066 28866
rect 12066 28814 12068 28866
rect 12012 28812 12068 28814
rect 12348 28028 12404 28084
rect 12572 28530 12628 28532
rect 12572 28478 12574 28530
rect 12574 28478 12626 28530
rect 12626 28478 12628 28530
rect 12572 28476 12628 28478
rect 12684 28028 12740 28084
rect 14476 40348 14532 40404
rect 13804 34802 13860 34804
rect 13804 34750 13806 34802
rect 13806 34750 13858 34802
rect 13858 34750 13860 34802
rect 13804 34748 13860 34750
rect 13692 33852 13748 33908
rect 13916 34130 13972 34132
rect 13916 34078 13918 34130
rect 13918 34078 13970 34130
rect 13970 34078 13972 34130
rect 13916 34076 13972 34078
rect 13580 30380 13636 30436
rect 13692 33628 13748 33684
rect 13580 30210 13636 30212
rect 13580 30158 13582 30210
rect 13582 30158 13634 30210
rect 13634 30158 13636 30210
rect 13580 30156 13636 30158
rect 14588 39564 14644 39620
rect 14812 40908 14868 40964
rect 15932 42754 15988 42756
rect 15932 42702 15934 42754
rect 15934 42702 15986 42754
rect 15986 42702 15988 42754
rect 15932 42700 15988 42702
rect 15932 42476 15988 42532
rect 15820 42364 15876 42420
rect 15260 41970 15316 41972
rect 15260 41918 15262 41970
rect 15262 41918 15314 41970
rect 15314 41918 15316 41970
rect 15260 41916 15316 41918
rect 15484 41970 15540 41972
rect 15484 41918 15486 41970
rect 15486 41918 15538 41970
rect 15538 41918 15540 41970
rect 15484 41916 15540 41918
rect 15708 41692 15764 41748
rect 15820 41186 15876 41188
rect 15820 41134 15822 41186
rect 15822 41134 15874 41186
rect 15874 41134 15876 41186
rect 15820 41132 15876 41134
rect 14588 38220 14644 38276
rect 14812 38050 14868 38052
rect 14812 37998 14814 38050
rect 14814 37998 14866 38050
rect 14866 37998 14868 38050
rect 14812 37996 14868 37998
rect 15148 40178 15204 40180
rect 15148 40126 15150 40178
rect 15150 40126 15202 40178
rect 15202 40126 15204 40178
rect 15148 40124 15204 40126
rect 15148 38444 15204 38500
rect 15484 39452 15540 39508
rect 16268 49196 16324 49252
rect 16268 45724 16324 45780
rect 16156 44322 16212 44324
rect 16156 44270 16158 44322
rect 16158 44270 16210 44322
rect 16210 44270 16212 44322
rect 16156 44268 16212 44270
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 20300 59164 20356 59220
rect 21756 60620 21812 60676
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19740 57820 19796 57876
rect 19404 57650 19460 57652
rect 19404 57598 19406 57650
rect 19406 57598 19458 57650
rect 19458 57598 19460 57650
rect 19404 57596 19460 57598
rect 19068 57484 19124 57540
rect 20300 57820 20356 57876
rect 19852 56812 19908 56868
rect 17836 53788 17892 53844
rect 17948 53618 18004 53620
rect 17948 53566 17950 53618
rect 17950 53566 18002 53618
rect 18002 53566 18004 53618
rect 17948 53564 18004 53566
rect 18284 54514 18340 54516
rect 18284 54462 18286 54514
rect 18286 54462 18338 54514
rect 18338 54462 18340 54514
rect 18284 54460 18340 54462
rect 19068 54460 19124 54516
rect 18732 53842 18788 53844
rect 18732 53790 18734 53842
rect 18734 53790 18786 53842
rect 18786 53790 18788 53842
rect 18732 53788 18788 53790
rect 17500 52946 17556 52948
rect 17500 52894 17502 52946
rect 17502 52894 17554 52946
rect 17554 52894 17556 52946
rect 17500 52892 17556 52894
rect 17388 49138 17444 49140
rect 17388 49086 17390 49138
rect 17390 49086 17442 49138
rect 17442 49086 17444 49138
rect 17388 49084 17444 49086
rect 16716 49026 16772 49028
rect 16716 48974 16718 49026
rect 16718 48974 16770 49026
rect 16770 48974 16772 49026
rect 16716 48972 16772 48974
rect 17836 47292 17892 47348
rect 17052 45890 17108 45892
rect 17052 45838 17054 45890
rect 17054 45838 17106 45890
rect 17106 45838 17108 45890
rect 17052 45836 17108 45838
rect 17724 45724 17780 45780
rect 16828 45276 16884 45332
rect 16380 43650 16436 43652
rect 16380 43598 16382 43650
rect 16382 43598 16434 43650
rect 16434 43598 16436 43650
rect 16380 43596 16436 43598
rect 16940 43484 16996 43540
rect 16828 42866 16884 42868
rect 16828 42814 16830 42866
rect 16830 42814 16882 42866
rect 16882 42814 16884 42866
rect 16828 42812 16884 42814
rect 16492 42754 16548 42756
rect 16492 42702 16494 42754
rect 16494 42702 16546 42754
rect 16546 42702 16548 42754
rect 16492 42700 16548 42702
rect 16828 42476 16884 42532
rect 16156 41132 16212 41188
rect 16268 42364 16324 42420
rect 16380 41692 16436 41748
rect 16716 41244 16772 41300
rect 17500 44268 17556 44324
rect 17276 42924 17332 42980
rect 17388 41804 17444 41860
rect 16940 41580 16996 41636
rect 15372 38610 15428 38612
rect 15372 38558 15374 38610
rect 15374 38558 15426 38610
rect 15426 38558 15428 38610
rect 15372 38556 15428 38558
rect 15484 38444 15540 38500
rect 15372 38274 15428 38276
rect 15372 38222 15374 38274
rect 15374 38222 15426 38274
rect 15426 38222 15428 38274
rect 15372 38220 15428 38222
rect 15596 38108 15652 38164
rect 15260 37772 15316 37828
rect 14812 37378 14868 37380
rect 14812 37326 14814 37378
rect 14814 37326 14866 37378
rect 14866 37326 14868 37378
rect 14812 37324 14868 37326
rect 15484 37996 15540 38052
rect 15596 37660 15652 37716
rect 15484 37266 15540 37268
rect 15484 37214 15486 37266
rect 15486 37214 15538 37266
rect 15538 37214 15540 37266
rect 15484 37212 15540 37214
rect 16492 40178 16548 40180
rect 16492 40126 16494 40178
rect 16494 40126 16546 40178
rect 16546 40126 16548 40178
rect 16492 40124 16548 40126
rect 16380 39564 16436 39620
rect 16492 39506 16548 39508
rect 16492 39454 16494 39506
rect 16494 39454 16546 39506
rect 16546 39454 16548 39506
rect 16492 39452 16548 39454
rect 15820 38780 15876 38836
rect 15932 37660 15988 37716
rect 16044 38220 16100 38276
rect 16044 37212 16100 37268
rect 16156 38108 16212 38164
rect 15820 37154 15876 37156
rect 15820 37102 15822 37154
rect 15822 37102 15874 37154
rect 15874 37102 15876 37154
rect 15820 37100 15876 37102
rect 15708 36316 15764 36372
rect 14924 35644 14980 35700
rect 17612 43538 17668 43540
rect 17612 43486 17614 43538
rect 17614 43486 17666 43538
rect 17666 43486 17668 43538
rect 17612 43484 17668 43486
rect 19404 53564 19460 53620
rect 18844 53506 18900 53508
rect 18844 53454 18846 53506
rect 18846 53454 18898 53506
rect 18898 53454 18900 53506
rect 18844 53452 18900 53454
rect 19180 52220 19236 52276
rect 20300 57650 20356 57652
rect 20300 57598 20302 57650
rect 20302 57598 20354 57650
rect 20354 57598 20356 57650
rect 20300 57596 20356 57598
rect 22652 61292 22708 61348
rect 23212 60674 23268 60676
rect 23212 60622 23214 60674
rect 23214 60622 23266 60674
rect 23266 60622 23268 60674
rect 23212 60620 23268 60622
rect 23996 64428 24052 64484
rect 23660 63756 23716 63812
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 39004 66444 39060 66500
rect 40796 66498 40852 66500
rect 40796 66446 40798 66498
rect 40798 66446 40850 66498
rect 40850 66446 40852 66498
rect 40796 66444 40852 66446
rect 33740 65436 33796 65492
rect 30268 64876 30324 64932
rect 25452 64428 25508 64484
rect 27804 64652 27860 64708
rect 26684 64204 26740 64260
rect 26348 63644 26404 63700
rect 24780 63196 24836 63252
rect 26236 63250 26292 63252
rect 26236 63198 26238 63250
rect 26238 63198 26290 63250
rect 26290 63198 26292 63250
rect 26236 63196 26292 63198
rect 26124 62860 26180 62916
rect 25900 62076 25956 62132
rect 23548 60620 23604 60676
rect 23996 59836 24052 59892
rect 21084 59164 21140 59220
rect 20748 57708 20804 57764
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20748 56866 20804 56868
rect 20748 56814 20750 56866
rect 20750 56814 20802 56866
rect 20802 56814 20804 56866
rect 20748 56812 20804 56814
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19628 54460 19684 54516
rect 20524 53788 20580 53844
rect 19852 53730 19908 53732
rect 19852 53678 19854 53730
rect 19854 53678 19906 53730
rect 19906 53678 19908 53730
rect 19852 53676 19908 53678
rect 19628 53506 19684 53508
rect 19628 53454 19630 53506
rect 19630 53454 19682 53506
rect 19682 53454 19684 53506
rect 19628 53452 19684 53454
rect 20076 53506 20132 53508
rect 20076 53454 20078 53506
rect 20078 53454 20130 53506
rect 20130 53454 20132 53506
rect 20076 53452 20132 53454
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20300 52834 20356 52836
rect 20300 52782 20302 52834
rect 20302 52782 20354 52834
rect 20354 52782 20356 52834
rect 20300 52780 20356 52782
rect 20636 53618 20692 53620
rect 20636 53566 20638 53618
rect 20638 53566 20690 53618
rect 20690 53566 20692 53618
rect 20636 53564 20692 53566
rect 20636 53228 20692 53284
rect 20636 52946 20692 52948
rect 20636 52894 20638 52946
rect 20638 52894 20690 52946
rect 20690 52894 20692 52946
rect 20636 52892 20692 52894
rect 20524 52780 20580 52836
rect 20300 52220 20356 52276
rect 20748 52274 20804 52276
rect 20748 52222 20750 52274
rect 20750 52222 20802 52274
rect 20802 52222 20804 52274
rect 20748 52220 20804 52222
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19516 49980 19572 50036
rect 19292 49922 19348 49924
rect 19292 49870 19294 49922
rect 19294 49870 19346 49922
rect 19346 49870 19348 49922
rect 19292 49868 19348 49870
rect 19516 49810 19572 49812
rect 19516 49758 19518 49810
rect 19518 49758 19570 49810
rect 19570 49758 19572 49810
rect 19516 49756 19572 49758
rect 19180 49644 19236 49700
rect 19068 48972 19124 49028
rect 18284 47346 18340 47348
rect 18284 47294 18286 47346
rect 18286 47294 18338 47346
rect 18338 47294 18340 47346
rect 18284 47292 18340 47294
rect 18508 46844 18564 46900
rect 18396 45778 18452 45780
rect 18396 45726 18398 45778
rect 18398 45726 18450 45778
rect 18450 45726 18452 45778
rect 18396 45724 18452 45726
rect 18508 44322 18564 44324
rect 18508 44270 18510 44322
rect 18510 44270 18562 44322
rect 18562 44270 18564 44322
rect 18508 44268 18564 44270
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20188 49868 20244 49924
rect 20076 49138 20132 49140
rect 20076 49086 20078 49138
rect 20078 49086 20130 49138
rect 20130 49086 20132 49138
rect 20076 49084 20132 49086
rect 19964 48914 20020 48916
rect 19964 48862 19966 48914
rect 19966 48862 20018 48914
rect 20018 48862 20020 48914
rect 19964 48860 20020 48862
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20524 49698 20580 49700
rect 20524 49646 20526 49698
rect 20526 49646 20578 49698
rect 20578 49646 20580 49698
rect 20524 49644 20580 49646
rect 20524 48914 20580 48916
rect 20524 48862 20526 48914
rect 20526 48862 20578 48914
rect 20578 48862 20580 48914
rect 20524 48860 20580 48862
rect 20300 48636 20356 48692
rect 20412 48748 20468 48804
rect 20972 48466 21028 48468
rect 20972 48414 20974 48466
rect 20974 48414 21026 48466
rect 21026 48414 21028 48466
rect 20972 48412 21028 48414
rect 21308 55580 21364 55636
rect 21196 53788 21252 53844
rect 26684 63138 26740 63140
rect 26684 63086 26686 63138
rect 26686 63086 26738 63138
rect 26738 63086 26740 63138
rect 26684 63084 26740 63086
rect 26460 63026 26516 63028
rect 26460 62974 26462 63026
rect 26462 62974 26514 63026
rect 26514 62974 26516 63026
rect 26460 62972 26516 62974
rect 27468 64204 27524 64260
rect 28140 64204 28196 64260
rect 27244 63644 27300 63700
rect 27132 63138 27188 63140
rect 27132 63086 27134 63138
rect 27134 63086 27186 63138
rect 27186 63086 27188 63138
rect 27132 63084 27188 63086
rect 27020 62914 27076 62916
rect 27020 62862 27022 62914
rect 27022 62862 27074 62914
rect 27074 62862 27076 62914
rect 27020 62860 27076 62862
rect 27244 62972 27300 63028
rect 27580 62860 27636 62916
rect 27244 62188 27300 62244
rect 28252 63644 28308 63700
rect 29148 64652 29204 64708
rect 28364 62188 28420 62244
rect 28476 62860 28532 62916
rect 27692 62076 27748 62132
rect 25564 61346 25620 61348
rect 25564 61294 25566 61346
rect 25566 61294 25618 61346
rect 25618 61294 25620 61346
rect 25564 61292 25620 61294
rect 25452 61010 25508 61012
rect 25452 60958 25454 61010
rect 25454 60958 25506 61010
rect 25506 60958 25508 61010
rect 25452 60956 25508 60958
rect 26012 61010 26068 61012
rect 26012 60958 26014 61010
rect 26014 60958 26066 61010
rect 26066 60958 26068 61010
rect 26012 60956 26068 60958
rect 25676 60620 25732 60676
rect 25900 60620 25956 60676
rect 25452 60508 25508 60564
rect 25228 58380 25284 58436
rect 22988 56140 23044 56196
rect 23660 56140 23716 56196
rect 23660 55468 23716 55524
rect 22316 53842 22372 53844
rect 22316 53790 22318 53842
rect 22318 53790 22370 53842
rect 22370 53790 22372 53842
rect 22316 53788 22372 53790
rect 26012 57708 26068 57764
rect 28140 61180 28196 61236
rect 27132 60620 27188 60676
rect 26572 59890 26628 59892
rect 26572 59838 26574 59890
rect 26574 59838 26626 59890
rect 26626 59838 26628 59890
rect 26572 59836 26628 59838
rect 27804 60898 27860 60900
rect 27804 60846 27806 60898
rect 27806 60846 27858 60898
rect 27858 60846 27860 60898
rect 27804 60844 27860 60846
rect 27244 60508 27300 60564
rect 27916 60786 27972 60788
rect 27916 60734 27918 60786
rect 27918 60734 27970 60786
rect 27970 60734 27972 60786
rect 27916 60732 27972 60734
rect 27692 60620 27748 60676
rect 28028 60508 28084 60564
rect 27468 59948 27524 60004
rect 26684 58434 26740 58436
rect 26684 58382 26686 58434
rect 26686 58382 26738 58434
rect 26738 58382 26740 58434
rect 26684 58380 26740 58382
rect 26684 56866 26740 56868
rect 26684 56814 26686 56866
rect 26686 56814 26738 56866
rect 26738 56814 26740 56866
rect 26684 56812 26740 56814
rect 24108 55916 24164 55972
rect 23324 53954 23380 53956
rect 23324 53902 23326 53954
rect 23326 53902 23378 53954
rect 23378 53902 23380 53954
rect 23324 53900 23380 53902
rect 24444 55468 24500 55524
rect 25340 55580 25396 55636
rect 24780 53900 24836 53956
rect 21308 53228 21364 53284
rect 23100 53618 23156 53620
rect 23100 53566 23102 53618
rect 23102 53566 23154 53618
rect 23154 53566 23156 53618
rect 23100 53564 23156 53566
rect 23548 53564 23604 53620
rect 23212 53506 23268 53508
rect 23212 53454 23214 53506
rect 23214 53454 23266 53506
rect 23266 53454 23268 53506
rect 23212 53452 23268 53454
rect 23100 52892 23156 52948
rect 23884 53452 23940 53508
rect 24332 53618 24388 53620
rect 24332 53566 24334 53618
rect 24334 53566 24386 53618
rect 24386 53566 24388 53618
rect 24332 53564 24388 53566
rect 24220 52946 24276 52948
rect 24220 52894 24222 52946
rect 24222 52894 24274 52946
rect 24274 52894 24276 52946
rect 24220 52892 24276 52894
rect 23100 52220 23156 52276
rect 24668 53170 24724 53172
rect 24668 53118 24670 53170
rect 24670 53118 24722 53170
rect 24722 53118 24724 53170
rect 24668 53116 24724 53118
rect 25340 53170 25396 53172
rect 25340 53118 25342 53170
rect 25342 53118 25394 53170
rect 25394 53118 25396 53170
rect 25340 53116 25396 53118
rect 22428 51436 22484 51492
rect 23772 51436 23828 51492
rect 21420 49810 21476 49812
rect 21420 49758 21422 49810
rect 21422 49758 21474 49810
rect 21474 49758 21476 49810
rect 21420 49756 21476 49758
rect 21420 48914 21476 48916
rect 21420 48862 21422 48914
rect 21422 48862 21474 48914
rect 21474 48862 21476 48914
rect 21420 48860 21476 48862
rect 21308 48802 21364 48804
rect 21308 48750 21310 48802
rect 21310 48750 21362 48802
rect 21362 48750 21364 48802
rect 21308 48748 21364 48750
rect 21532 48636 21588 48692
rect 21980 48412 22036 48468
rect 23548 49084 23604 49140
rect 22540 49026 22596 49028
rect 22540 48974 22542 49026
rect 22542 48974 22594 49026
rect 22594 48974 22596 49026
rect 22540 48972 22596 48974
rect 22988 49026 23044 49028
rect 22988 48974 22990 49026
rect 22990 48974 23042 49026
rect 23042 48974 23044 49026
rect 22988 48972 23044 48974
rect 23324 48412 23380 48468
rect 21532 47628 21588 47684
rect 22652 47682 22708 47684
rect 22652 47630 22654 47682
rect 22654 47630 22706 47682
rect 22706 47630 22708 47682
rect 22652 47628 22708 47630
rect 23100 47570 23156 47572
rect 23100 47518 23102 47570
rect 23102 47518 23154 47570
rect 23154 47518 23156 47570
rect 23100 47516 23156 47518
rect 21084 47180 21140 47236
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20188 46844 20244 46900
rect 19404 46674 19460 46676
rect 19404 46622 19406 46674
rect 19406 46622 19458 46674
rect 19458 46622 19460 46674
rect 19404 46620 19460 46622
rect 19740 46450 19796 46452
rect 19740 46398 19742 46450
rect 19742 46398 19794 46450
rect 19794 46398 19796 46450
rect 19740 46396 19796 46398
rect 19068 45948 19124 46004
rect 22988 46060 23044 46116
rect 20748 45666 20804 45668
rect 20748 45614 20750 45666
rect 20750 45614 20802 45666
rect 20802 45614 20804 45666
rect 20748 45612 20804 45614
rect 21420 45666 21476 45668
rect 21420 45614 21422 45666
rect 21422 45614 21474 45666
rect 21474 45614 21476 45666
rect 21420 45612 21476 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22316 45330 22372 45332
rect 22316 45278 22318 45330
rect 22318 45278 22370 45330
rect 22370 45278 22372 45330
rect 22316 45276 22372 45278
rect 21644 45164 21700 45220
rect 20972 44268 21028 44324
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20524 43596 20580 43652
rect 19740 43426 19796 43428
rect 19740 43374 19742 43426
rect 19742 43374 19794 43426
rect 19794 43374 19796 43426
rect 19740 43372 19796 43374
rect 19628 43148 19684 43204
rect 20188 42978 20244 42980
rect 20188 42926 20190 42978
rect 20190 42926 20242 42978
rect 20242 42926 20244 42978
rect 20188 42924 20244 42926
rect 18060 42588 18116 42644
rect 17836 42140 17892 42196
rect 18060 41468 18116 41524
rect 18284 41132 18340 41188
rect 17388 40124 17444 40180
rect 17500 39618 17556 39620
rect 17500 39566 17502 39618
rect 17502 39566 17554 39618
rect 17554 39566 17556 39618
rect 17500 39564 17556 39566
rect 16828 38780 16884 38836
rect 16604 38162 16660 38164
rect 16604 38110 16606 38162
rect 16606 38110 16658 38162
rect 16658 38110 16660 38162
rect 16604 38108 16660 38110
rect 16380 37266 16436 37268
rect 16380 37214 16382 37266
rect 16382 37214 16434 37266
rect 16434 37214 16436 37266
rect 16380 37212 16436 37214
rect 17724 39730 17780 39732
rect 17724 39678 17726 39730
rect 17726 39678 17778 39730
rect 17778 39678 17780 39730
rect 17724 39676 17780 39678
rect 17612 37996 17668 38052
rect 17724 38668 17780 38724
rect 17052 37938 17108 37940
rect 17052 37886 17054 37938
rect 17054 37886 17106 37938
rect 17106 37886 17108 37938
rect 17052 37884 17108 37886
rect 16828 37324 16884 37380
rect 16268 37100 16324 37156
rect 17276 37212 17332 37268
rect 17164 36876 17220 36932
rect 15932 36428 15988 36484
rect 16828 36428 16884 36484
rect 14812 33628 14868 33684
rect 13916 31836 13972 31892
rect 12572 27132 12628 27188
rect 12236 27020 12292 27076
rect 9996 25452 10052 25508
rect 11004 26178 11060 26180
rect 11004 26126 11006 26178
rect 11006 26126 11058 26178
rect 11058 26126 11060 26178
rect 11004 26124 11060 26126
rect 10780 24610 10836 24612
rect 10780 24558 10782 24610
rect 10782 24558 10834 24610
rect 10834 24558 10836 24610
rect 10780 24556 10836 24558
rect 13468 27692 13524 27748
rect 13916 29932 13972 29988
rect 11788 25564 11844 25620
rect 12236 25506 12292 25508
rect 12236 25454 12238 25506
rect 12238 25454 12290 25506
rect 12290 25454 12292 25506
rect 12236 25452 12292 25454
rect 12796 25506 12852 25508
rect 12796 25454 12798 25506
rect 12798 25454 12850 25506
rect 12850 25454 12852 25506
rect 12796 25452 12852 25454
rect 11564 25394 11620 25396
rect 11564 25342 11566 25394
rect 11566 25342 11618 25394
rect 11618 25342 11620 25394
rect 11564 25340 11620 25342
rect 14252 31612 14308 31668
rect 15036 31388 15092 31444
rect 14812 30210 14868 30212
rect 14812 30158 14814 30210
rect 14814 30158 14866 30210
rect 14866 30158 14868 30210
rect 14812 30156 14868 30158
rect 16156 35698 16212 35700
rect 16156 35646 16158 35698
rect 16158 35646 16210 35698
rect 16210 35646 16212 35698
rect 16156 35644 16212 35646
rect 18060 38834 18116 38836
rect 18060 38782 18062 38834
rect 18062 38782 18114 38834
rect 18114 38782 18116 38834
rect 18060 38780 18116 38782
rect 17948 38668 18004 38724
rect 18396 40348 18452 40404
rect 20300 42642 20356 42644
rect 20300 42590 20302 42642
rect 20302 42590 20354 42642
rect 20354 42590 20356 42642
rect 20300 42588 20356 42590
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 21644 44268 21700 44324
rect 23212 45276 23268 45332
rect 22204 45218 22260 45220
rect 22204 45166 22206 45218
rect 22206 45166 22258 45218
rect 22258 45166 22260 45218
rect 22204 45164 22260 45166
rect 21756 45052 21812 45108
rect 22428 45106 22484 45108
rect 22428 45054 22430 45106
rect 22430 45054 22482 45106
rect 22482 45054 22484 45106
rect 22428 45052 22484 45054
rect 22316 44940 22372 44996
rect 22092 44322 22148 44324
rect 22092 44270 22094 44322
rect 22094 44270 22146 44322
rect 22146 44270 22148 44322
rect 22092 44268 22148 44270
rect 20972 43484 21028 43540
rect 22540 43932 22596 43988
rect 23100 44994 23156 44996
rect 23100 44942 23102 44994
rect 23102 44942 23154 44994
rect 23154 44942 23156 44994
rect 23100 44940 23156 44942
rect 23884 48130 23940 48132
rect 23884 48078 23886 48130
rect 23886 48078 23938 48130
rect 23938 48078 23940 48130
rect 23884 48076 23940 48078
rect 23660 47458 23716 47460
rect 23660 47406 23662 47458
rect 23662 47406 23714 47458
rect 23714 47406 23716 47458
rect 23660 47404 23716 47406
rect 24444 49084 24500 49140
rect 25116 48972 25172 49028
rect 24668 48130 24724 48132
rect 24668 48078 24670 48130
rect 24670 48078 24722 48130
rect 24722 48078 24724 48130
rect 24668 48076 24724 48078
rect 24332 47516 24388 47572
rect 24556 47458 24612 47460
rect 24556 47406 24558 47458
rect 24558 47406 24610 47458
rect 24610 47406 24612 47458
rect 24556 47404 24612 47406
rect 24892 48076 24948 48132
rect 24332 47234 24388 47236
rect 24332 47182 24334 47234
rect 24334 47182 24386 47234
rect 24386 47182 24388 47234
rect 24332 47180 24388 47182
rect 24668 47180 24724 47236
rect 23660 47068 23716 47124
rect 24556 46898 24612 46900
rect 24556 46846 24558 46898
rect 24558 46846 24610 46898
rect 24610 46846 24612 46898
rect 24556 46844 24612 46846
rect 23548 46674 23604 46676
rect 23548 46622 23550 46674
rect 23550 46622 23602 46674
rect 23602 46622 23604 46674
rect 23548 46620 23604 46622
rect 23660 46060 23716 46116
rect 24892 47068 24948 47124
rect 25452 47234 25508 47236
rect 25452 47182 25454 47234
rect 25454 47182 25506 47234
rect 25506 47182 25508 47234
rect 25452 47180 25508 47182
rect 25452 46956 25508 47012
rect 25228 46620 25284 46676
rect 23436 44380 23492 44436
rect 24108 44434 24164 44436
rect 24108 44382 24110 44434
rect 24110 44382 24162 44434
rect 24162 44382 24164 44434
rect 24108 44380 24164 44382
rect 22876 43932 22932 43988
rect 22316 43426 22372 43428
rect 22316 43374 22318 43426
rect 22318 43374 22370 43426
rect 22370 43374 22372 43426
rect 22316 43372 22372 43374
rect 20860 43148 20916 43204
rect 19404 41804 19460 41860
rect 17948 38108 18004 38164
rect 17500 35420 17556 35476
rect 16604 34914 16660 34916
rect 16604 34862 16606 34914
rect 16606 34862 16658 34914
rect 16658 34862 16660 34914
rect 16604 34860 16660 34862
rect 15708 30156 15764 30212
rect 17948 36428 18004 36484
rect 17612 34076 17668 34132
rect 15596 29986 15652 29988
rect 15596 29934 15598 29986
rect 15598 29934 15650 29986
rect 15650 29934 15652 29986
rect 15596 29932 15652 29934
rect 15372 29596 15428 29652
rect 14140 28924 14196 28980
rect 14700 29314 14756 29316
rect 14700 29262 14702 29314
rect 14702 29262 14754 29314
rect 14754 29262 14756 29314
rect 14700 29260 14756 29262
rect 14812 29036 14868 29092
rect 13580 27020 13636 27076
rect 13468 26962 13524 26964
rect 13468 26910 13470 26962
rect 13470 26910 13522 26962
rect 13522 26910 13524 26962
rect 13468 26908 13524 26910
rect 14700 28642 14756 28644
rect 14700 28590 14702 28642
rect 14702 28590 14754 28642
rect 14754 28590 14756 28642
rect 14700 28588 14756 28590
rect 14140 28530 14196 28532
rect 14140 28478 14142 28530
rect 14142 28478 14194 28530
rect 14194 28478 14196 28530
rect 14140 28476 14196 28478
rect 14028 28418 14084 28420
rect 14028 28366 14030 28418
rect 14030 28366 14082 28418
rect 14082 28366 14084 28418
rect 14028 28364 14084 28366
rect 14924 28252 14980 28308
rect 14364 27692 14420 27748
rect 14588 27132 14644 27188
rect 14252 27020 14308 27076
rect 15596 29036 15652 29092
rect 15148 28476 15204 28532
rect 15148 27468 15204 27524
rect 13692 26348 13748 26404
rect 13244 25564 13300 25620
rect 13356 25452 13412 25508
rect 13916 25452 13972 25508
rect 14476 26572 14532 26628
rect 14028 25394 14084 25396
rect 14028 25342 14030 25394
rect 14030 25342 14082 25394
rect 14082 25342 14084 25394
rect 14028 25340 14084 25342
rect 14140 25116 14196 25172
rect 13916 24668 13972 24724
rect 14028 24610 14084 24612
rect 14028 24558 14030 24610
rect 14030 24558 14082 24610
rect 14082 24558 14084 24610
rect 14028 24556 14084 24558
rect 14252 24556 14308 24612
rect 15596 26402 15652 26404
rect 15596 26350 15598 26402
rect 15598 26350 15650 26402
rect 15650 26350 15652 26402
rect 15596 26348 15652 26350
rect 15484 25900 15540 25956
rect 15484 25618 15540 25620
rect 15484 25566 15486 25618
rect 15486 25566 15538 25618
rect 15538 25566 15540 25618
rect 15484 25564 15540 25566
rect 14700 25452 14756 25508
rect 15148 25116 15204 25172
rect 17836 34914 17892 34916
rect 17836 34862 17838 34914
rect 17838 34862 17890 34914
rect 17890 34862 17892 34914
rect 17836 34860 17892 34862
rect 17948 34802 18004 34804
rect 17948 34750 17950 34802
rect 17950 34750 18002 34802
rect 18002 34750 18004 34802
rect 17948 34748 18004 34750
rect 18844 39730 18900 39732
rect 18844 39678 18846 39730
rect 18846 39678 18898 39730
rect 18898 39678 18900 39730
rect 18844 39676 18900 39678
rect 18956 41020 19012 41076
rect 19964 41746 20020 41748
rect 19964 41694 19966 41746
rect 19966 41694 20018 41746
rect 20018 41694 20020 41746
rect 19964 41692 20020 41694
rect 20076 41298 20132 41300
rect 20076 41246 20078 41298
rect 20078 41246 20130 41298
rect 20130 41246 20132 41298
rect 20076 41244 20132 41246
rect 19852 41186 19908 41188
rect 19852 41134 19854 41186
rect 19854 41134 19906 41186
rect 19906 41134 19908 41186
rect 19852 41132 19908 41134
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20300 41916 20356 41972
rect 20300 40796 20356 40852
rect 20524 41074 20580 41076
rect 20524 41022 20526 41074
rect 20526 41022 20578 41074
rect 20578 41022 20580 41074
rect 20524 41020 20580 41022
rect 19068 39564 19124 39620
rect 18844 38892 18900 38948
rect 18620 38722 18676 38724
rect 18620 38670 18622 38722
rect 18622 38670 18674 38722
rect 18674 38670 18676 38722
rect 18620 38668 18676 38670
rect 18508 38556 18564 38612
rect 18956 38220 19012 38276
rect 18508 38050 18564 38052
rect 18508 37998 18510 38050
rect 18510 37998 18562 38050
rect 18562 37998 18564 38050
rect 18508 37996 18564 37998
rect 18508 37100 18564 37156
rect 18620 37772 18676 37828
rect 18508 34802 18564 34804
rect 18508 34750 18510 34802
rect 18510 34750 18562 34802
rect 18562 34750 18564 34802
rect 18508 34748 18564 34750
rect 15932 33234 15988 33236
rect 15932 33182 15934 33234
rect 15934 33182 15986 33234
rect 15986 33182 15988 33234
rect 15932 33180 15988 33182
rect 17948 31948 18004 32004
rect 17500 31836 17556 31892
rect 16268 30156 16324 30212
rect 16044 29426 16100 29428
rect 16044 29374 16046 29426
rect 16046 29374 16098 29426
rect 16098 29374 16100 29426
rect 16044 29372 16100 29374
rect 16716 31388 16772 31444
rect 16604 29932 16660 29988
rect 16492 29538 16548 29540
rect 16492 29486 16494 29538
rect 16494 29486 16546 29538
rect 16546 29486 16548 29538
rect 16492 29484 16548 29486
rect 16156 28530 16212 28532
rect 16156 28478 16158 28530
rect 16158 28478 16210 28530
rect 16210 28478 16212 28530
rect 16156 28476 16212 28478
rect 18284 34130 18340 34132
rect 18284 34078 18286 34130
rect 18286 34078 18338 34130
rect 18338 34078 18340 34130
rect 18284 34076 18340 34078
rect 18620 33234 18676 33236
rect 18620 33182 18622 33234
rect 18622 33182 18674 33234
rect 18674 33182 18676 33234
rect 18620 33180 18676 33182
rect 18508 33068 18564 33124
rect 19180 40460 19236 40516
rect 20300 40402 20356 40404
rect 20300 40350 20302 40402
rect 20302 40350 20354 40402
rect 20354 40350 20356 40402
rect 20300 40348 20356 40350
rect 20188 39564 20244 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19292 38892 19348 38948
rect 18956 37884 19012 37940
rect 19068 37212 19124 37268
rect 18844 36316 18900 36372
rect 19180 35420 19236 35476
rect 19180 34130 19236 34132
rect 19180 34078 19182 34130
rect 19182 34078 19234 34130
rect 19234 34078 19236 34130
rect 19180 34076 19236 34078
rect 18844 33346 18900 33348
rect 18844 33294 18846 33346
rect 18846 33294 18898 33346
rect 18898 33294 18900 33346
rect 18844 33292 18900 33294
rect 19068 32956 19124 33012
rect 18956 31836 19012 31892
rect 17948 29708 18004 29764
rect 18060 29932 18116 29988
rect 17276 29538 17332 29540
rect 17276 29486 17278 29538
rect 17278 29486 17330 29538
rect 17330 29486 17332 29538
rect 17276 29484 17332 29486
rect 16492 28418 16548 28420
rect 16492 28366 16494 28418
rect 16494 28366 16546 28418
rect 16546 28366 16548 28418
rect 16492 28364 16548 28366
rect 17612 28476 17668 28532
rect 17724 28364 17780 28420
rect 17612 27970 17668 27972
rect 17612 27918 17614 27970
rect 17614 27918 17666 27970
rect 17666 27918 17668 27970
rect 17612 27916 17668 27918
rect 18172 27580 18228 27636
rect 15932 26796 15988 26852
rect 15932 26402 15988 26404
rect 15932 26350 15934 26402
rect 15934 26350 15986 26402
rect 15986 26350 15988 26402
rect 15932 26348 15988 26350
rect 17836 27468 17892 27524
rect 15932 25618 15988 25620
rect 15932 25566 15934 25618
rect 15934 25566 15986 25618
rect 15986 25566 15988 25618
rect 15932 25564 15988 25566
rect 16268 25506 16324 25508
rect 16268 25454 16270 25506
rect 16270 25454 16322 25506
rect 16322 25454 16324 25506
rect 16268 25452 16324 25454
rect 16044 24946 16100 24948
rect 16044 24894 16046 24946
rect 16046 24894 16098 24946
rect 16098 24894 16100 24946
rect 16044 24892 16100 24894
rect 15820 24668 15876 24724
rect 15596 24610 15652 24612
rect 15596 24558 15598 24610
rect 15598 24558 15650 24610
rect 15650 24558 15652 24610
rect 15596 24556 15652 24558
rect 16380 24668 16436 24724
rect 16828 26124 16884 26180
rect 17388 26236 17444 26292
rect 16716 24892 16772 24948
rect 16268 24556 16324 24612
rect 16716 24444 16772 24500
rect 16268 23772 16324 23828
rect 17388 25452 17444 25508
rect 17724 26124 17780 26180
rect 17724 25452 17780 25508
rect 17388 24946 17444 24948
rect 17388 24894 17390 24946
rect 17390 24894 17442 24946
rect 17442 24894 17444 24946
rect 17388 24892 17444 24894
rect 18844 29372 18900 29428
rect 18620 27916 18676 27972
rect 18956 27580 19012 27636
rect 18060 26290 18116 26292
rect 18060 26238 18062 26290
rect 18062 26238 18114 26290
rect 18114 26238 18116 26290
rect 18060 26236 18116 26238
rect 17612 24834 17668 24836
rect 17612 24782 17614 24834
rect 17614 24782 17666 24834
rect 17666 24782 17668 24834
rect 17612 24780 17668 24782
rect 18060 24892 18116 24948
rect 17836 24722 17892 24724
rect 17836 24670 17838 24722
rect 17838 24670 17890 24722
rect 17890 24670 17892 24722
rect 17836 24668 17892 24670
rect 18732 25116 18788 25172
rect 18620 24834 18676 24836
rect 18620 24782 18622 24834
rect 18622 24782 18674 24834
rect 18674 24782 18676 24834
rect 18620 24780 18676 24782
rect 18172 24668 18228 24724
rect 17836 24444 17892 24500
rect 17276 23826 17332 23828
rect 17276 23774 17278 23826
rect 17278 23774 17330 23826
rect 17330 23774 17332 23826
rect 17276 23772 17332 23774
rect 19852 38556 19908 38612
rect 20412 38946 20468 38948
rect 20412 38894 20414 38946
rect 20414 38894 20466 38946
rect 20466 38894 20468 38946
rect 20412 38892 20468 38894
rect 20188 38332 20244 38388
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19628 37436 19684 37492
rect 19404 37324 19460 37380
rect 20188 37436 20244 37492
rect 19740 37154 19796 37156
rect 19740 37102 19742 37154
rect 19742 37102 19794 37154
rect 19794 37102 19796 37154
rect 19740 37100 19796 37102
rect 20748 41692 20804 41748
rect 20748 40236 20804 40292
rect 20636 38220 20692 38276
rect 22092 43148 22148 43204
rect 21420 42530 21476 42532
rect 21420 42478 21422 42530
rect 21422 42478 21474 42530
rect 21474 42478 21476 42530
rect 21420 42476 21476 42478
rect 20972 42194 21028 42196
rect 20972 42142 20974 42194
rect 20974 42142 21026 42194
rect 21026 42142 21028 42194
rect 20972 42140 21028 42142
rect 21084 41916 21140 41972
rect 20972 40626 21028 40628
rect 20972 40574 20974 40626
rect 20974 40574 21026 40626
rect 21026 40574 21028 40626
rect 20972 40572 21028 40574
rect 21196 41858 21252 41860
rect 21196 41806 21198 41858
rect 21198 41806 21250 41858
rect 21250 41806 21252 41858
rect 21196 41804 21252 41806
rect 21420 41580 21476 41636
rect 21308 41468 21364 41524
rect 22652 42028 22708 42084
rect 22316 40962 22372 40964
rect 22316 40910 22318 40962
rect 22318 40910 22370 40962
rect 22370 40910 22372 40962
rect 22316 40908 22372 40910
rect 21420 40626 21476 40628
rect 21420 40574 21422 40626
rect 21422 40574 21474 40626
rect 21474 40574 21476 40626
rect 21420 40572 21476 40574
rect 22204 39730 22260 39732
rect 22204 39678 22206 39730
rect 22206 39678 22258 39730
rect 22258 39678 22260 39730
rect 22204 39676 22260 39678
rect 22988 40796 23044 40852
rect 22428 39116 22484 39172
rect 20412 37266 20468 37268
rect 20412 37214 20414 37266
rect 20414 37214 20466 37266
rect 20466 37214 20468 37266
rect 20412 37212 20468 37214
rect 20748 37154 20804 37156
rect 20748 37102 20750 37154
rect 20750 37102 20802 37154
rect 20802 37102 20804 37154
rect 20748 37100 20804 37102
rect 20300 36876 20356 36932
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20860 35420 20916 35476
rect 21308 38332 21364 38388
rect 23212 43932 23268 43988
rect 23660 43932 23716 43988
rect 23100 40684 23156 40740
rect 23324 40572 23380 40628
rect 23772 41298 23828 41300
rect 23772 41246 23774 41298
rect 23774 41246 23826 41298
rect 23826 41246 23828 41298
rect 23772 41244 23828 41246
rect 23436 40796 23492 40852
rect 23884 40796 23940 40852
rect 23436 39676 23492 39732
rect 23212 39116 23268 39172
rect 22988 37884 23044 37940
rect 22876 37154 22932 37156
rect 22876 37102 22878 37154
rect 22878 37102 22930 37154
rect 22930 37102 22932 37154
rect 22876 37100 22932 37102
rect 21308 35586 21364 35588
rect 21308 35534 21310 35586
rect 21310 35534 21362 35586
rect 21362 35534 21364 35586
rect 21308 35532 21364 35534
rect 19516 34076 19572 34132
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19516 33292 19572 33348
rect 19404 33122 19460 33124
rect 19404 33070 19406 33122
rect 19406 33070 19458 33122
rect 19458 33070 19460 33122
rect 19404 33068 19460 33070
rect 19516 32956 19572 33012
rect 19404 32450 19460 32452
rect 19404 32398 19406 32450
rect 19406 32398 19458 32450
rect 19458 32398 19460 32450
rect 19404 32396 19460 32398
rect 19180 30156 19236 30212
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20188 32284 20244 32340
rect 20188 31948 20244 32004
rect 20748 32396 20804 32452
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 30828 20356 30884
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19180 28082 19236 28084
rect 19180 28030 19182 28082
rect 19182 28030 19234 28082
rect 19234 28030 19236 28082
rect 19180 28028 19236 28030
rect 19516 28028 19572 28084
rect 19628 27858 19684 27860
rect 19628 27806 19630 27858
rect 19630 27806 19682 27858
rect 19682 27806 19684 27858
rect 19628 27804 19684 27806
rect 21196 30882 21252 30884
rect 21196 30830 21198 30882
rect 21198 30830 21250 30882
rect 21250 30830 21252 30882
rect 21196 30828 21252 30830
rect 20412 29260 20468 29316
rect 21644 33404 21700 33460
rect 21420 33068 21476 33124
rect 22204 33180 22260 33236
rect 21980 30940 22036 30996
rect 22204 31106 22260 31108
rect 22204 31054 22206 31106
rect 22206 31054 22258 31106
rect 22258 31054 22260 31106
rect 22204 31052 22260 31054
rect 22092 30828 22148 30884
rect 22204 30380 22260 30436
rect 21868 30156 21924 30212
rect 21308 29708 21364 29764
rect 21084 29596 21140 29652
rect 21756 29596 21812 29652
rect 22540 30994 22596 30996
rect 22540 30942 22542 30994
rect 22542 30942 22594 30994
rect 22594 30942 22596 30994
rect 22540 30940 22596 30942
rect 22316 30210 22372 30212
rect 22316 30158 22318 30210
rect 22318 30158 22370 30210
rect 22370 30158 22372 30210
rect 22316 30156 22372 30158
rect 22204 29932 22260 29988
rect 22764 35868 22820 35924
rect 22764 35698 22820 35700
rect 22764 35646 22766 35698
rect 22766 35646 22818 35698
rect 22818 35646 22820 35698
rect 22764 35644 22820 35646
rect 22764 33516 22820 33572
rect 22876 30994 22932 30996
rect 22876 30942 22878 30994
rect 22878 30942 22930 30994
rect 22930 30942 22932 30994
rect 22876 30940 22932 30942
rect 24220 41746 24276 41748
rect 24220 41694 24222 41746
rect 24222 41694 24274 41746
rect 24274 41694 24276 41746
rect 24220 41692 24276 41694
rect 24668 44994 24724 44996
rect 24668 44942 24670 44994
rect 24670 44942 24722 44994
rect 24722 44942 24724 44994
rect 24668 44940 24724 44942
rect 24444 44268 24500 44324
rect 24780 44322 24836 44324
rect 24780 44270 24782 44322
rect 24782 44270 24834 44322
rect 24834 44270 24836 44322
rect 24780 44268 24836 44270
rect 25340 44268 25396 44324
rect 25564 44940 25620 44996
rect 25564 44380 25620 44436
rect 24332 40908 24388 40964
rect 23772 40572 23828 40628
rect 24556 42082 24612 42084
rect 24556 42030 24558 42082
rect 24558 42030 24610 42082
rect 24610 42030 24612 42082
rect 24556 42028 24612 42030
rect 25228 41244 25284 41300
rect 26796 56754 26852 56756
rect 26796 56702 26798 56754
rect 26798 56702 26850 56754
rect 26850 56702 26852 56754
rect 26796 56700 26852 56702
rect 26684 54626 26740 54628
rect 26684 54574 26686 54626
rect 26686 54574 26738 54626
rect 26738 54574 26740 54626
rect 26684 54572 26740 54574
rect 26236 50482 26292 50484
rect 26236 50430 26238 50482
rect 26238 50430 26290 50482
rect 26290 50430 26292 50482
rect 26236 50428 26292 50430
rect 28364 60226 28420 60228
rect 28364 60174 28366 60226
rect 28366 60174 28418 60226
rect 28418 60174 28420 60226
rect 28364 60172 28420 60174
rect 28252 57762 28308 57764
rect 28252 57710 28254 57762
rect 28254 57710 28306 57762
rect 28306 57710 28308 57762
rect 28252 57708 28308 57710
rect 27132 56754 27188 56756
rect 27132 56702 27134 56754
rect 27134 56702 27186 56754
rect 27186 56702 27188 56754
rect 27132 56700 27188 56702
rect 27020 55804 27076 55860
rect 27692 56642 27748 56644
rect 27692 56590 27694 56642
rect 27694 56590 27746 56642
rect 27746 56590 27748 56642
rect 27692 56588 27748 56590
rect 28924 62860 28980 62916
rect 29484 64706 29540 64708
rect 29484 64654 29486 64706
rect 29486 64654 29538 64706
rect 29538 64654 29540 64706
rect 29484 64652 29540 64654
rect 30380 64706 30436 64708
rect 30380 64654 30382 64706
rect 30382 64654 30434 64706
rect 30434 64654 30436 64706
rect 30380 64652 30436 64654
rect 30940 64594 30996 64596
rect 30940 64542 30942 64594
rect 30942 64542 30994 64594
rect 30994 64542 30996 64594
rect 30940 64540 30996 64542
rect 30156 63138 30212 63140
rect 30156 63086 30158 63138
rect 30158 63086 30210 63138
rect 30210 63086 30212 63138
rect 30156 63084 30212 63086
rect 29484 62860 29540 62916
rect 29484 62188 29540 62244
rect 30940 63084 30996 63140
rect 31276 63084 31332 63140
rect 31500 62914 31556 62916
rect 31500 62862 31502 62914
rect 31502 62862 31554 62914
rect 31554 62862 31556 62914
rect 31500 62860 31556 62862
rect 32956 64594 33012 64596
rect 32956 64542 32958 64594
rect 32958 64542 33010 64594
rect 33010 64542 33012 64594
rect 32956 64540 33012 64542
rect 33292 64482 33348 64484
rect 33292 64430 33294 64482
rect 33294 64430 33346 64482
rect 33346 64430 33348 64482
rect 33292 64428 33348 64430
rect 32508 63922 32564 63924
rect 32508 63870 32510 63922
rect 32510 63870 32562 63922
rect 32562 63870 32564 63922
rect 32508 63868 32564 63870
rect 32396 63810 32452 63812
rect 32396 63758 32398 63810
rect 32398 63758 32450 63810
rect 32450 63758 32452 63810
rect 32396 63756 32452 63758
rect 32060 62914 32116 62916
rect 32060 62862 32062 62914
rect 32062 62862 32114 62914
rect 32114 62862 32116 62914
rect 32060 62860 32116 62862
rect 32620 63980 32676 64036
rect 33180 63868 33236 63924
rect 32844 62860 32900 62916
rect 32060 62412 32116 62468
rect 29596 61068 29652 61124
rect 28924 60786 28980 60788
rect 28924 60734 28926 60786
rect 28926 60734 28978 60786
rect 28978 60734 28980 60786
rect 28924 60732 28980 60734
rect 28700 60674 28756 60676
rect 28700 60622 28702 60674
rect 28702 60622 28754 60674
rect 28754 60622 28756 60674
rect 28700 60620 28756 60622
rect 29260 60172 29316 60228
rect 29372 60002 29428 60004
rect 29372 59950 29374 60002
rect 29374 59950 29426 60002
rect 29426 59950 29428 60002
rect 29372 59948 29428 59950
rect 32956 62412 33012 62468
rect 29932 60562 29988 60564
rect 29932 60510 29934 60562
rect 29934 60510 29986 60562
rect 29986 60510 29988 60562
rect 29932 60508 29988 60510
rect 30380 59948 30436 60004
rect 29820 58322 29876 58324
rect 29820 58270 29822 58322
rect 29822 58270 29874 58322
rect 29874 58270 29876 58322
rect 29820 58268 29876 58270
rect 31164 59724 31220 59780
rect 32060 60508 32116 60564
rect 32396 60732 32452 60788
rect 32396 60002 32452 60004
rect 32396 59950 32398 60002
rect 32398 59950 32450 60002
rect 32450 59950 32452 60002
rect 32396 59948 32452 59950
rect 31612 59052 31668 59108
rect 30380 58044 30436 58100
rect 30492 58322 30548 58324
rect 30492 58270 30494 58322
rect 30494 58270 30546 58322
rect 30546 58270 30548 58322
rect 30492 58268 30548 58270
rect 30044 57260 30100 57316
rect 30156 57596 30212 57652
rect 27020 55020 27076 55076
rect 27580 54514 27636 54516
rect 27580 54462 27582 54514
rect 27582 54462 27634 54514
rect 27634 54462 27636 54514
rect 27580 54460 27636 54462
rect 27916 55074 27972 55076
rect 27916 55022 27918 55074
rect 27918 55022 27970 55074
rect 27970 55022 27972 55074
rect 27916 55020 27972 55022
rect 28140 53842 28196 53844
rect 28140 53790 28142 53842
rect 28142 53790 28194 53842
rect 28194 53790 28196 53842
rect 28140 53788 28196 53790
rect 28476 54402 28532 54404
rect 28476 54350 28478 54402
rect 28478 54350 28530 54402
rect 28530 54350 28532 54402
rect 28476 54348 28532 54350
rect 29148 54402 29204 54404
rect 29148 54350 29150 54402
rect 29150 54350 29202 54402
rect 29202 54350 29204 54402
rect 29148 54348 29204 54350
rect 29372 55020 29428 55076
rect 30604 57260 30660 57316
rect 30940 57650 30996 57652
rect 30940 57598 30942 57650
rect 30942 57598 30994 57650
rect 30994 57598 30996 57650
rect 30940 57596 30996 57598
rect 30716 55186 30772 55188
rect 30716 55134 30718 55186
rect 30718 55134 30770 55186
rect 30770 55134 30772 55186
rect 30716 55132 30772 55134
rect 29372 53954 29428 53956
rect 29372 53902 29374 53954
rect 29374 53902 29426 53954
rect 29426 53902 29428 53954
rect 29372 53900 29428 53902
rect 28924 53788 28980 53844
rect 28924 53452 28980 53508
rect 28476 51378 28532 51380
rect 28476 51326 28478 51378
rect 28478 51326 28530 51378
rect 28530 51326 28532 51378
rect 28476 51324 28532 51326
rect 25788 49138 25844 49140
rect 25788 49086 25790 49138
rect 25790 49086 25842 49138
rect 25842 49086 25844 49138
rect 25788 49084 25844 49086
rect 26124 48188 26180 48244
rect 26908 47740 26964 47796
rect 26012 46508 26068 46564
rect 26236 46562 26292 46564
rect 26236 46510 26238 46562
rect 26238 46510 26290 46562
rect 26290 46510 26292 46562
rect 26236 46508 26292 46510
rect 26236 45724 26292 45780
rect 27020 45836 27076 45892
rect 26012 42754 26068 42756
rect 26012 42702 26014 42754
rect 26014 42702 26066 42754
rect 26066 42702 26068 42754
rect 26012 42700 26068 42702
rect 25564 41132 25620 41188
rect 25564 40908 25620 40964
rect 24444 40572 24500 40628
rect 23660 39564 23716 39620
rect 23884 40402 23940 40404
rect 23884 40350 23886 40402
rect 23886 40350 23938 40402
rect 23938 40350 23940 40402
rect 23884 40348 23940 40350
rect 23548 37548 23604 37604
rect 23324 35922 23380 35924
rect 23324 35870 23326 35922
rect 23326 35870 23378 35922
rect 23378 35870 23380 35922
rect 23324 35868 23380 35870
rect 23660 35644 23716 35700
rect 23324 35308 23380 35364
rect 25004 39676 25060 39732
rect 24668 39564 24724 39620
rect 24220 39340 24276 39396
rect 23884 38834 23940 38836
rect 23884 38782 23886 38834
rect 23886 38782 23938 38834
rect 23938 38782 23940 38834
rect 23884 38780 23940 38782
rect 24332 38892 24388 38948
rect 23996 37938 24052 37940
rect 23996 37886 23998 37938
rect 23998 37886 24050 37938
rect 24050 37886 24052 37938
rect 23996 37884 24052 37886
rect 24556 38668 24612 38724
rect 24668 38108 24724 38164
rect 23996 37548 24052 37604
rect 23884 37436 23940 37492
rect 23996 36876 24052 36932
rect 26012 41132 26068 41188
rect 26572 41692 26628 41748
rect 28364 50540 28420 50596
rect 27356 49420 27412 49476
rect 27244 47740 27300 47796
rect 27468 48242 27524 48244
rect 27468 48190 27470 48242
rect 27470 48190 27522 48242
rect 27522 48190 27524 48242
rect 27468 48188 27524 48190
rect 27244 47292 27300 47348
rect 27356 46508 27412 46564
rect 27468 45948 27524 46004
rect 27244 45890 27300 45892
rect 27244 45838 27246 45890
rect 27246 45838 27298 45890
rect 27298 45838 27300 45890
rect 27244 45836 27300 45838
rect 27132 42754 27188 42756
rect 27132 42702 27134 42754
rect 27134 42702 27186 42754
rect 27186 42702 27188 42754
rect 27132 42700 27188 42702
rect 27244 42082 27300 42084
rect 27244 42030 27246 42082
rect 27246 42030 27298 42082
rect 27298 42030 27300 42082
rect 27244 42028 27300 42030
rect 27468 41244 27524 41300
rect 27692 42588 27748 42644
rect 26908 41132 26964 41188
rect 26460 41074 26516 41076
rect 26460 41022 26462 41074
rect 26462 41022 26514 41074
rect 26514 41022 26516 41074
rect 26460 41020 26516 41022
rect 26348 40124 26404 40180
rect 26124 39730 26180 39732
rect 26124 39678 26126 39730
rect 26126 39678 26178 39730
rect 26178 39678 26180 39730
rect 26124 39676 26180 39678
rect 25564 39452 25620 39508
rect 25340 37490 25396 37492
rect 25340 37438 25342 37490
rect 25342 37438 25394 37490
rect 25394 37438 25396 37490
rect 25340 37436 25396 37438
rect 25228 37154 25284 37156
rect 25228 37102 25230 37154
rect 25230 37102 25282 37154
rect 25282 37102 25284 37154
rect 25228 37100 25284 37102
rect 24332 36482 24388 36484
rect 24332 36430 24334 36482
rect 24334 36430 24386 36482
rect 24386 36430 24388 36482
rect 24332 36428 24388 36430
rect 24220 35980 24276 36036
rect 23548 33516 23604 33572
rect 25228 36876 25284 36932
rect 23884 33068 23940 33124
rect 25228 35980 25284 36036
rect 25452 35532 25508 35588
rect 26236 39618 26292 39620
rect 26236 39566 26238 39618
rect 26238 39566 26290 39618
rect 26290 39566 26292 39618
rect 26236 39564 26292 39566
rect 26572 39452 26628 39508
rect 27356 41020 27412 41076
rect 26684 39004 26740 39060
rect 27132 38892 27188 38948
rect 26348 38834 26404 38836
rect 26348 38782 26350 38834
rect 26350 38782 26402 38834
rect 26402 38782 26404 38834
rect 26348 38780 26404 38782
rect 27244 40348 27300 40404
rect 25676 38668 25732 38724
rect 26012 38668 26068 38724
rect 26124 38444 26180 38500
rect 26796 38332 26852 38388
rect 26908 38444 26964 38500
rect 26572 37996 26628 38052
rect 26012 37826 26068 37828
rect 26012 37774 26014 37826
rect 26014 37774 26066 37826
rect 26066 37774 26068 37826
rect 26012 37772 26068 37774
rect 26124 37378 26180 37380
rect 26124 37326 26126 37378
rect 26126 37326 26178 37378
rect 26178 37326 26180 37378
rect 26124 37324 26180 37326
rect 26796 37212 26852 37268
rect 26012 36876 26068 36932
rect 27020 38162 27076 38164
rect 27020 38110 27022 38162
rect 27022 38110 27074 38162
rect 27074 38110 27076 38162
rect 27020 38108 27076 38110
rect 27132 37324 27188 37380
rect 27468 40962 27524 40964
rect 27468 40910 27470 40962
rect 27470 40910 27522 40962
rect 27522 40910 27524 40962
rect 27468 40908 27524 40910
rect 29148 51378 29204 51380
rect 29148 51326 29150 51378
rect 29150 51326 29202 51378
rect 29202 51326 29204 51378
rect 29148 51324 29204 51326
rect 29036 50764 29092 50820
rect 29372 50652 29428 50708
rect 29260 50594 29316 50596
rect 29260 50542 29262 50594
rect 29262 50542 29314 50594
rect 29314 50542 29316 50594
rect 29260 50540 29316 50542
rect 28700 50034 28756 50036
rect 28700 49982 28702 50034
rect 28702 49982 28754 50034
rect 28754 49982 28756 50034
rect 28700 49980 28756 49982
rect 29036 49756 29092 49812
rect 27916 47458 27972 47460
rect 27916 47406 27918 47458
rect 27918 47406 27970 47458
rect 27970 47406 27972 47458
rect 27916 47404 27972 47406
rect 28252 47346 28308 47348
rect 28252 47294 28254 47346
rect 28254 47294 28306 47346
rect 28306 47294 28308 47346
rect 28252 47292 28308 47294
rect 28364 47068 28420 47124
rect 30380 53788 30436 53844
rect 30044 53506 30100 53508
rect 30044 53454 30046 53506
rect 30046 53454 30098 53506
rect 30098 53454 30100 53506
rect 30044 53452 30100 53454
rect 30604 53452 30660 53508
rect 30716 53676 30772 53732
rect 32284 59106 32340 59108
rect 32284 59054 32286 59106
rect 32286 59054 32338 59106
rect 32338 59054 32340 59106
rect 32284 59052 32340 59054
rect 32284 57484 32340 57540
rect 32844 57484 32900 57540
rect 31612 57260 31668 57316
rect 32396 56924 32452 56980
rect 31612 55244 31668 55300
rect 31052 54348 31108 54404
rect 30828 52892 30884 52948
rect 30716 52780 30772 52836
rect 30940 52162 30996 52164
rect 30940 52110 30942 52162
rect 30942 52110 30994 52162
rect 30994 52110 30996 52162
rect 30940 52108 30996 52110
rect 29596 50540 29652 50596
rect 30156 50594 30212 50596
rect 30156 50542 30158 50594
rect 30158 50542 30210 50594
rect 30210 50542 30212 50594
rect 30156 50540 30212 50542
rect 30604 50482 30660 50484
rect 30604 50430 30606 50482
rect 30606 50430 30658 50482
rect 30658 50430 30660 50482
rect 30604 50428 30660 50430
rect 29932 50316 29988 50372
rect 29820 49980 29876 50036
rect 30492 49756 30548 49812
rect 28588 47068 28644 47124
rect 27916 45052 27972 45108
rect 28028 42364 28084 42420
rect 27916 42028 27972 42084
rect 28028 41916 28084 41972
rect 28140 41804 28196 41860
rect 27692 41132 27748 41188
rect 27580 40348 27636 40404
rect 27804 40460 27860 40516
rect 27916 41074 27972 41076
rect 27916 41022 27918 41074
rect 27918 41022 27970 41074
rect 27970 41022 27972 41074
rect 27916 41020 27972 41022
rect 28028 40908 28084 40964
rect 27468 39394 27524 39396
rect 27468 39342 27470 39394
rect 27470 39342 27522 39394
rect 27522 39342 27524 39394
rect 27468 39340 27524 39342
rect 27692 39058 27748 39060
rect 27692 39006 27694 39058
rect 27694 39006 27746 39058
rect 27746 39006 27748 39058
rect 27692 39004 27748 39006
rect 28028 38834 28084 38836
rect 28028 38782 28030 38834
rect 28030 38782 28082 38834
rect 28082 38782 28084 38834
rect 28028 38780 28084 38782
rect 28700 46786 28756 46788
rect 28700 46734 28702 46786
rect 28702 46734 28754 46786
rect 28754 46734 28756 46786
rect 28700 46732 28756 46734
rect 30492 48748 30548 48804
rect 29372 47068 29428 47124
rect 29820 46786 29876 46788
rect 29820 46734 29822 46786
rect 29822 46734 29874 46786
rect 29874 46734 29876 46786
rect 29820 46732 29876 46734
rect 29820 45948 29876 46004
rect 30940 50652 30996 50708
rect 30828 50482 30884 50484
rect 30828 50430 30830 50482
rect 30830 50430 30882 50482
rect 30882 50430 30884 50482
rect 30828 50428 30884 50430
rect 31052 49698 31108 49700
rect 31052 49646 31054 49698
rect 31054 49646 31106 49698
rect 31106 49646 31108 49698
rect 31052 49644 31108 49646
rect 30940 48972 30996 49028
rect 30156 46172 30212 46228
rect 28476 45106 28532 45108
rect 28476 45054 28478 45106
rect 28478 45054 28530 45106
rect 28530 45054 28532 45106
rect 28476 45052 28532 45054
rect 29148 45052 29204 45108
rect 28364 42812 28420 42868
rect 28476 42530 28532 42532
rect 28476 42478 28478 42530
rect 28478 42478 28530 42530
rect 28530 42478 28532 42530
rect 28476 42476 28532 42478
rect 28364 42364 28420 42420
rect 29148 42754 29204 42756
rect 29148 42702 29150 42754
rect 29150 42702 29202 42754
rect 29202 42702 29204 42754
rect 29148 42700 29204 42702
rect 28924 42252 28980 42308
rect 29820 43650 29876 43652
rect 29820 43598 29822 43650
rect 29822 43598 29874 43650
rect 29874 43598 29876 43650
rect 29820 43596 29876 43598
rect 29932 42812 29988 42868
rect 29708 42588 29764 42644
rect 28476 42028 28532 42084
rect 28812 42140 28868 42196
rect 29484 41970 29540 41972
rect 29484 41918 29486 41970
rect 29486 41918 29538 41970
rect 29538 41918 29540 41970
rect 29484 41916 29540 41918
rect 28924 40572 28980 40628
rect 28588 40124 28644 40180
rect 28364 38556 28420 38612
rect 27468 38050 27524 38052
rect 27468 37998 27470 38050
rect 27470 37998 27522 38050
rect 27522 37998 27524 38050
rect 27468 37996 27524 37998
rect 28252 37996 28308 38052
rect 27580 37884 27636 37940
rect 28140 37938 28196 37940
rect 28140 37886 28142 37938
rect 28142 37886 28194 37938
rect 28194 37886 28196 37938
rect 28140 37884 28196 37886
rect 27580 37436 27636 37492
rect 28364 37826 28420 37828
rect 28364 37774 28366 37826
rect 28366 37774 28418 37826
rect 28418 37774 28420 37826
rect 28364 37772 28420 37774
rect 26908 36482 26964 36484
rect 26908 36430 26910 36482
rect 26910 36430 26962 36482
rect 26962 36430 26964 36482
rect 26908 36428 26964 36430
rect 27244 35922 27300 35924
rect 27244 35870 27246 35922
rect 27246 35870 27298 35922
rect 27298 35870 27300 35922
rect 27244 35868 27300 35870
rect 28588 38050 28644 38052
rect 28588 37998 28590 38050
rect 28590 37998 28642 38050
rect 28642 37998 28644 38050
rect 28588 37996 28644 37998
rect 29484 40348 29540 40404
rect 30044 42140 30100 42196
rect 29708 40572 29764 40628
rect 30156 41468 30212 41524
rect 31052 46172 31108 46228
rect 31052 46002 31108 46004
rect 31052 45950 31054 46002
rect 31054 45950 31106 46002
rect 31106 45950 31108 46002
rect 31052 45948 31108 45950
rect 31276 53900 31332 53956
rect 31500 55186 31556 55188
rect 31500 55134 31502 55186
rect 31502 55134 31554 55186
rect 31554 55134 31556 55186
rect 31500 55132 31556 55134
rect 32508 56194 32564 56196
rect 32508 56142 32510 56194
rect 32510 56142 32562 56194
rect 32562 56142 32564 56194
rect 32508 56140 32564 56142
rect 32284 55244 32340 55300
rect 31948 54402 32004 54404
rect 31948 54350 31950 54402
rect 31950 54350 32002 54402
rect 32002 54350 32004 54402
rect 31948 54348 32004 54350
rect 32508 54236 32564 54292
rect 31388 53788 31444 53844
rect 31276 53170 31332 53172
rect 31276 53118 31278 53170
rect 31278 53118 31330 53170
rect 31330 53118 31332 53170
rect 31276 53116 31332 53118
rect 30940 43596 30996 43652
rect 31276 52892 31332 52948
rect 31164 44322 31220 44324
rect 31164 44270 31166 44322
rect 31166 44270 31218 44322
rect 31218 44270 31220 44322
rect 31164 44268 31220 44270
rect 32172 53116 32228 53172
rect 31948 52834 32004 52836
rect 31948 52782 31950 52834
rect 31950 52782 32002 52834
rect 32002 52782 32004 52834
rect 31948 52780 32004 52782
rect 32508 52332 32564 52388
rect 32396 52274 32452 52276
rect 32396 52222 32398 52274
rect 32398 52222 32450 52274
rect 32450 52222 32452 52274
rect 32396 52220 32452 52222
rect 31836 52162 31892 52164
rect 31836 52110 31838 52162
rect 31838 52110 31890 52162
rect 31890 52110 31892 52162
rect 31836 52108 31892 52110
rect 32284 50764 32340 50820
rect 31724 49026 31780 49028
rect 31724 48974 31726 49026
rect 31726 48974 31778 49026
rect 31778 48974 31780 49026
rect 31724 48972 31780 48974
rect 31500 46732 31556 46788
rect 31388 46562 31444 46564
rect 31388 46510 31390 46562
rect 31390 46510 31442 46562
rect 31442 46510 31444 46562
rect 31388 46508 31444 46510
rect 31724 46562 31780 46564
rect 31724 46510 31726 46562
rect 31726 46510 31778 46562
rect 31778 46510 31780 46562
rect 31724 46508 31780 46510
rect 31500 45218 31556 45220
rect 31500 45166 31502 45218
rect 31502 45166 31554 45218
rect 31554 45166 31556 45218
rect 31500 45164 31556 45166
rect 31388 44434 31444 44436
rect 31388 44382 31390 44434
rect 31390 44382 31442 44434
rect 31442 44382 31444 44434
rect 31388 44380 31444 44382
rect 32508 49644 32564 49700
rect 32732 49756 32788 49812
rect 32284 49196 32340 49252
rect 31948 46508 32004 46564
rect 31948 46172 32004 46228
rect 32060 45724 32116 45780
rect 32060 44380 32116 44436
rect 31948 44268 32004 44324
rect 30940 42476 30996 42532
rect 30492 41804 30548 41860
rect 31276 42642 31332 42644
rect 31276 42590 31278 42642
rect 31278 42590 31330 42642
rect 31330 42590 31332 42642
rect 31276 42588 31332 42590
rect 30268 40460 30324 40516
rect 30156 39228 30212 39284
rect 30380 39004 30436 39060
rect 30044 38834 30100 38836
rect 30044 38782 30046 38834
rect 30046 38782 30098 38834
rect 30098 38782 30100 38834
rect 30044 38780 30100 38782
rect 29260 38444 29316 38500
rect 29932 38722 29988 38724
rect 29932 38670 29934 38722
rect 29934 38670 29986 38722
rect 29986 38670 29988 38722
rect 29932 38668 29988 38670
rect 28700 37772 28756 37828
rect 29148 37996 29204 38052
rect 29260 37938 29316 37940
rect 29260 37886 29262 37938
rect 29262 37886 29314 37938
rect 29314 37886 29316 37938
rect 29260 37884 29316 37886
rect 29372 37212 29428 37268
rect 27356 35532 27412 35588
rect 25676 35308 25732 35364
rect 27916 35026 27972 35028
rect 27916 34974 27918 35026
rect 27918 34974 27970 35026
rect 27970 34974 27972 35026
rect 27916 34972 27972 34974
rect 29148 34972 29204 35028
rect 28364 34412 28420 34468
rect 25116 33404 25172 33460
rect 24668 33122 24724 33124
rect 24668 33070 24670 33122
rect 24670 33070 24722 33122
rect 24722 33070 24724 33122
rect 24668 33068 24724 33070
rect 28140 33346 28196 33348
rect 28140 33294 28142 33346
rect 28142 33294 28194 33346
rect 28194 33294 28196 33346
rect 28140 33292 28196 33294
rect 25788 33234 25844 33236
rect 25788 33182 25790 33234
rect 25790 33182 25842 33234
rect 25842 33182 25844 33234
rect 25788 33180 25844 33182
rect 24108 31836 24164 31892
rect 22988 30380 23044 30436
rect 23436 30994 23492 30996
rect 23436 30942 23438 30994
rect 23438 30942 23490 30994
rect 23490 30942 23492 30994
rect 23436 30940 23492 30942
rect 22764 29932 22820 29988
rect 21532 29538 21588 29540
rect 21532 29486 21534 29538
rect 21534 29486 21586 29538
rect 21586 29486 21588 29538
rect 21532 29484 21588 29486
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 18956 24892 19012 24948
rect 19404 24892 19460 24948
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 18732 23660 18788 23716
rect 18956 23772 19012 23828
rect 18956 22540 19012 22596
rect 18620 21810 18676 21812
rect 18620 21758 18622 21810
rect 18622 21758 18674 21810
rect 18674 21758 18676 21810
rect 18620 21756 18676 21758
rect 15820 20690 15876 20692
rect 15820 20638 15822 20690
rect 15822 20638 15874 20690
rect 15874 20638 15876 20690
rect 15820 20636 15876 20638
rect 15036 20076 15092 20132
rect 19292 21810 19348 21812
rect 19292 21758 19294 21810
rect 19294 21758 19346 21810
rect 19346 21758 19348 21810
rect 19292 21756 19348 21758
rect 16716 20076 16772 20132
rect 18956 21698 19012 21700
rect 18956 21646 18958 21698
rect 18958 21646 19010 21698
rect 19010 21646 19012 21698
rect 18956 21644 19012 21646
rect 17724 19964 17780 20020
rect 18060 20130 18116 20132
rect 18060 20078 18062 20130
rect 18062 20078 18114 20130
rect 18114 20078 18116 20130
rect 18060 20076 18116 20078
rect 15148 18396 15204 18452
rect 18620 20860 18676 20916
rect 18396 20690 18452 20692
rect 18396 20638 18398 20690
rect 18398 20638 18450 20690
rect 18450 20638 18452 20690
rect 18396 20636 18452 20638
rect 18508 20524 18564 20580
rect 18620 20018 18676 20020
rect 18620 19966 18622 20018
rect 18622 19966 18674 20018
rect 18674 19966 18676 20018
rect 18620 19964 18676 19966
rect 17276 18956 17332 19012
rect 14700 17388 14756 17444
rect 16828 17052 16884 17108
rect 16604 16940 16660 16996
rect 11004 16268 11060 16324
rect 5852 11676 5908 11732
rect 14028 16044 14084 16100
rect 15820 16716 15876 16772
rect 15820 16098 15876 16100
rect 15820 16046 15822 16098
rect 15822 16046 15874 16098
rect 15874 16046 15876 16098
rect 15820 16044 15876 16046
rect 18508 19010 18564 19012
rect 18508 18958 18510 19010
rect 18510 18958 18562 19010
rect 18562 18958 18564 19010
rect 18508 18956 18564 18958
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 18284 18450 18340 18452
rect 18284 18398 18286 18450
rect 18286 18398 18338 18450
rect 18338 18398 18340 18450
rect 18284 18396 18340 18398
rect 17500 17442 17556 17444
rect 17500 17390 17502 17442
rect 17502 17390 17554 17442
rect 17554 17390 17556 17442
rect 17500 17388 17556 17390
rect 17388 17276 17444 17332
rect 18284 17442 18340 17444
rect 18284 17390 18286 17442
rect 18286 17390 18338 17442
rect 18338 17390 18340 17442
rect 18284 17388 18340 17390
rect 18396 17276 18452 17332
rect 17724 17164 17780 17220
rect 18284 17164 18340 17220
rect 18060 17052 18116 17108
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 17276 14588 17332 14644
rect 14700 13916 14756 13972
rect 16828 13804 16884 13860
rect 14028 13580 14084 13636
rect 17500 13634 17556 13636
rect 17500 13582 17502 13634
rect 17502 13582 17554 13634
rect 17554 13582 17556 13634
rect 17500 13580 17556 13582
rect 17836 13186 17892 13188
rect 17836 13134 17838 13186
rect 17838 13134 17890 13186
rect 17890 13134 17892 13186
rect 17836 13132 17892 13134
rect 17948 12850 18004 12852
rect 17948 12798 17950 12850
rect 17950 12798 18002 12850
rect 18002 12798 18004 12850
rect 17948 12796 18004 12798
rect 17836 12738 17892 12740
rect 17836 12686 17838 12738
rect 17838 12686 17890 12738
rect 17890 12686 17892 12738
rect 17836 12684 17892 12686
rect 17276 11506 17332 11508
rect 17276 11454 17278 11506
rect 17278 11454 17330 11506
rect 17330 11454 17332 11506
rect 17276 11452 17332 11454
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 15932 11116 15988 11172
rect 14364 10108 14420 10164
rect 17500 10108 17556 10164
rect 15932 9938 15988 9940
rect 15932 9886 15934 9938
rect 15934 9886 15986 9938
rect 15986 9886 15988 9938
rect 15932 9884 15988 9886
rect 16828 9660 16884 9716
rect 14700 9548 14756 9604
rect 15820 9602 15876 9604
rect 15820 9550 15822 9602
rect 15822 9550 15874 9602
rect 15874 9550 15876 9602
rect 15820 9548 15876 9550
rect 17724 11340 17780 11396
rect 18508 17052 18564 17108
rect 18620 16994 18676 16996
rect 18620 16942 18622 16994
rect 18622 16942 18674 16994
rect 18674 16942 18676 16994
rect 18620 16940 18676 16942
rect 19068 18620 19124 18676
rect 19068 18450 19124 18452
rect 19068 18398 19070 18450
rect 19070 18398 19122 18450
rect 19122 18398 19124 18450
rect 19068 18396 19124 18398
rect 18956 17500 19012 17556
rect 19292 20914 19348 20916
rect 19292 20862 19294 20914
rect 19294 20862 19346 20914
rect 19346 20862 19348 20914
rect 19292 20860 19348 20862
rect 19852 23660 19908 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 22540 19796 22596
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19964 21810 20020 21812
rect 19964 21758 19966 21810
rect 19966 21758 20018 21810
rect 20018 21758 20020 21810
rect 19964 21756 20020 21758
rect 20076 21644 20132 21700
rect 20300 20860 20356 20916
rect 21532 29314 21588 29316
rect 21532 29262 21534 29314
rect 21534 29262 21586 29314
rect 21586 29262 21588 29314
rect 21532 29260 21588 29262
rect 20748 29148 20804 29204
rect 19628 20524 19684 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19404 20076 19460 20132
rect 19292 19292 19348 19348
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19292 18620 19348 18676
rect 19852 17666 19908 17668
rect 19852 17614 19854 17666
rect 19854 17614 19906 17666
rect 19906 17614 19908 17666
rect 19852 17612 19908 17614
rect 19180 17388 19236 17444
rect 18284 14642 18340 14644
rect 18284 14590 18286 14642
rect 18286 14590 18338 14642
rect 18338 14590 18340 14642
rect 18284 14588 18340 14590
rect 18508 14530 18564 14532
rect 18508 14478 18510 14530
rect 18510 14478 18562 14530
rect 18562 14478 18564 14530
rect 18508 14476 18564 14478
rect 18508 13804 18564 13860
rect 18284 13132 18340 13188
rect 18284 11900 18340 11956
rect 18284 11452 18340 11508
rect 17724 10108 17780 10164
rect 17612 9772 17668 9828
rect 18732 16210 18788 16212
rect 18732 16158 18734 16210
rect 18734 16158 18786 16210
rect 18786 16158 18788 16210
rect 18732 16156 18788 16158
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16882 19684 16884
rect 19628 16830 19630 16882
rect 19630 16830 19682 16882
rect 19682 16830 19684 16882
rect 19628 16828 19684 16830
rect 19404 16156 19460 16212
rect 22092 29538 22148 29540
rect 22092 29486 22094 29538
rect 22094 29486 22146 29538
rect 22146 29486 22148 29538
rect 22092 29484 22148 29486
rect 21644 29148 21700 29204
rect 22428 29538 22484 29540
rect 22428 29486 22430 29538
rect 22430 29486 22482 29538
rect 22482 29486 22484 29538
rect 22428 29484 22484 29486
rect 22316 26514 22372 26516
rect 22316 26462 22318 26514
rect 22318 26462 22370 26514
rect 22370 26462 22372 26514
rect 22316 26460 22372 26462
rect 20748 25116 20804 25172
rect 21756 25228 21812 25284
rect 22540 25282 22596 25284
rect 22540 25230 22542 25282
rect 22542 25230 22594 25282
rect 22594 25230 22596 25282
rect 22540 25228 22596 25230
rect 21644 23884 21700 23940
rect 22204 23938 22260 23940
rect 22204 23886 22206 23938
rect 22206 23886 22258 23938
rect 22258 23886 22260 23938
rect 22204 23884 22260 23886
rect 20748 23714 20804 23716
rect 20748 23662 20750 23714
rect 20750 23662 20802 23714
rect 20802 23662 20804 23714
rect 20748 23660 20804 23662
rect 21980 23436 22036 23492
rect 22428 23548 22484 23604
rect 22876 29650 22932 29652
rect 22876 29598 22878 29650
rect 22878 29598 22930 29650
rect 22930 29598 22932 29650
rect 22876 29596 22932 29598
rect 22876 27858 22932 27860
rect 22876 27806 22878 27858
rect 22878 27806 22930 27858
rect 22930 27806 22932 27858
rect 22876 27804 22932 27806
rect 22876 26908 22932 26964
rect 22764 24780 22820 24836
rect 22652 24668 22708 24724
rect 22764 23548 22820 23604
rect 22652 23436 22708 23492
rect 20748 22652 20804 22708
rect 20524 21644 20580 21700
rect 21756 21586 21812 21588
rect 21756 21534 21758 21586
rect 21758 21534 21810 21586
rect 21810 21534 21812 21586
rect 21756 21532 21812 21534
rect 20748 20690 20804 20692
rect 20748 20638 20750 20690
rect 20750 20638 20802 20690
rect 20802 20638 20804 20690
rect 20748 20636 20804 20638
rect 21980 20690 22036 20692
rect 21980 20638 21982 20690
rect 21982 20638 22034 20690
rect 22034 20638 22036 20690
rect 21980 20636 22036 20638
rect 21868 20578 21924 20580
rect 21868 20526 21870 20578
rect 21870 20526 21922 20578
rect 21922 20526 21924 20578
rect 21868 20524 21924 20526
rect 22764 23266 22820 23268
rect 22764 23214 22766 23266
rect 22766 23214 22818 23266
rect 22818 23214 22820 23266
rect 22764 23212 22820 23214
rect 22988 23154 23044 23156
rect 22988 23102 22990 23154
rect 22990 23102 23042 23154
rect 23042 23102 23044 23154
rect 22988 23100 23044 23102
rect 22764 21644 22820 21700
rect 23212 29650 23268 29652
rect 23212 29598 23214 29650
rect 23214 29598 23266 29650
rect 23266 29598 23268 29650
rect 23212 29596 23268 29598
rect 23996 30994 24052 30996
rect 23996 30942 23998 30994
rect 23998 30942 24050 30994
rect 24050 30942 24052 30994
rect 23996 30940 24052 30942
rect 23996 30156 24052 30212
rect 24220 30098 24276 30100
rect 24220 30046 24222 30098
rect 24222 30046 24274 30098
rect 24274 30046 24276 30098
rect 24220 30044 24276 30046
rect 24444 29986 24500 29988
rect 24444 29934 24446 29986
rect 24446 29934 24498 29986
rect 24498 29934 24500 29986
rect 24444 29932 24500 29934
rect 23660 29538 23716 29540
rect 23660 29486 23662 29538
rect 23662 29486 23714 29538
rect 23714 29486 23716 29538
rect 23660 29484 23716 29486
rect 24780 29372 24836 29428
rect 23436 27692 23492 27748
rect 23324 26460 23380 26516
rect 23996 26908 24052 26964
rect 23772 26460 23828 26516
rect 23436 25900 23492 25956
rect 23884 25506 23940 25508
rect 23884 25454 23886 25506
rect 23886 25454 23938 25506
rect 23938 25454 23940 25506
rect 23884 25452 23940 25454
rect 23212 25340 23268 25396
rect 23436 25228 23492 25284
rect 21644 17724 21700 17780
rect 21196 17388 21252 17444
rect 23212 24780 23268 24836
rect 22540 18284 22596 18340
rect 22316 17778 22372 17780
rect 22316 17726 22318 17778
rect 22318 17726 22370 17778
rect 22370 17726 22372 17778
rect 22316 17724 22372 17726
rect 23436 24722 23492 24724
rect 23436 24670 23438 24722
rect 23438 24670 23490 24722
rect 23490 24670 23492 24722
rect 23436 24668 23492 24670
rect 23324 23436 23380 23492
rect 24556 26850 24612 26852
rect 24556 26798 24558 26850
rect 24558 26798 24610 26850
rect 24610 26798 24612 26850
rect 24556 26796 24612 26798
rect 24220 26124 24276 26180
rect 24444 25900 24500 25956
rect 24108 25676 24164 25732
rect 24220 25506 24276 25508
rect 24220 25454 24222 25506
rect 24222 25454 24274 25506
rect 24274 25454 24276 25506
rect 24220 25452 24276 25454
rect 24332 23436 24388 23492
rect 23996 23324 24052 23380
rect 23884 22258 23940 22260
rect 23884 22206 23886 22258
rect 23886 22206 23938 22258
rect 23938 22206 23940 22258
rect 23884 22204 23940 22206
rect 28364 33628 28420 33684
rect 28252 33180 28308 33236
rect 27804 33068 27860 33124
rect 29372 34690 29428 34692
rect 29372 34638 29374 34690
rect 29374 34638 29426 34690
rect 29426 34638 29428 34690
rect 29372 34636 29428 34638
rect 28812 33628 28868 33684
rect 30604 37938 30660 37940
rect 30604 37886 30606 37938
rect 30606 37886 30658 37938
rect 30658 37886 30660 37938
rect 30604 37884 30660 37886
rect 30268 37324 30324 37380
rect 31164 40460 31220 40516
rect 30940 39340 30996 39396
rect 31276 39004 31332 39060
rect 30940 38780 30996 38836
rect 30828 38610 30884 38612
rect 30828 38558 30830 38610
rect 30830 38558 30882 38610
rect 30882 38558 30884 38610
rect 30828 38556 30884 38558
rect 30828 37826 30884 37828
rect 30828 37774 30830 37826
rect 30830 37774 30882 37826
rect 30882 37774 30884 37826
rect 30828 37772 30884 37774
rect 29708 35644 29764 35700
rect 31276 37436 31332 37492
rect 31500 37884 31556 37940
rect 31388 37324 31444 37380
rect 30492 35698 30548 35700
rect 30492 35646 30494 35698
rect 30494 35646 30546 35698
rect 30546 35646 30548 35698
rect 30492 35644 30548 35646
rect 29820 34914 29876 34916
rect 29820 34862 29822 34914
rect 29822 34862 29874 34914
rect 29874 34862 29876 34914
rect 29820 34860 29876 34862
rect 29596 34188 29652 34244
rect 30044 34636 30100 34692
rect 30940 34972 30996 35028
rect 30716 34860 30772 34916
rect 29820 33964 29876 34020
rect 29484 33404 29540 33460
rect 28924 33292 28980 33348
rect 28700 33068 28756 33124
rect 29372 33068 29428 33124
rect 26796 31890 26852 31892
rect 26796 31838 26798 31890
rect 26798 31838 26850 31890
rect 26850 31838 26852 31890
rect 26796 31836 26852 31838
rect 25900 30156 25956 30212
rect 25452 29932 25508 29988
rect 25228 29372 25284 29428
rect 25452 29036 25508 29092
rect 25564 29650 25620 29652
rect 25564 29598 25566 29650
rect 25566 29598 25618 29650
rect 25618 29598 25620 29650
rect 25564 29596 25620 29598
rect 25564 28812 25620 28868
rect 25788 27692 25844 27748
rect 28140 30156 28196 30212
rect 26460 29260 26516 29316
rect 26908 29650 26964 29652
rect 26908 29598 26910 29650
rect 26910 29598 26962 29650
rect 26962 29598 26964 29650
rect 26908 29596 26964 29598
rect 27804 29650 27860 29652
rect 27804 29598 27806 29650
rect 27806 29598 27858 29650
rect 27858 29598 27860 29650
rect 27804 29596 27860 29598
rect 27692 29538 27748 29540
rect 27692 29486 27694 29538
rect 27694 29486 27746 29538
rect 27746 29486 27748 29538
rect 27692 29484 27748 29486
rect 27580 29372 27636 29428
rect 27692 29314 27748 29316
rect 27692 29262 27694 29314
rect 27694 29262 27746 29314
rect 27746 29262 27748 29314
rect 27692 29260 27748 29262
rect 26908 29148 26964 29204
rect 28588 30716 28644 30772
rect 29932 31052 29988 31108
rect 29708 30828 29764 30884
rect 29596 30268 29652 30324
rect 28476 29538 28532 29540
rect 28476 29486 28478 29538
rect 28478 29486 28530 29538
rect 28530 29486 28532 29538
rect 28476 29484 28532 29486
rect 28140 29260 28196 29316
rect 28700 29148 28756 29204
rect 28476 28812 28532 28868
rect 28364 28588 28420 28644
rect 28812 28588 28868 28644
rect 28700 28028 28756 28084
rect 28924 28082 28980 28084
rect 28924 28030 28926 28082
rect 28926 28030 28978 28082
rect 28978 28030 28980 28082
rect 28924 28028 28980 28030
rect 24668 26012 24724 26068
rect 24556 25676 24612 25732
rect 24556 25394 24612 25396
rect 24556 25342 24558 25394
rect 24558 25342 24610 25394
rect 24610 25342 24612 25394
rect 24556 25340 24612 25342
rect 24892 23548 24948 23604
rect 24220 23154 24276 23156
rect 24220 23102 24222 23154
rect 24222 23102 24274 23154
rect 24274 23102 24276 23154
rect 24220 23100 24276 23102
rect 24444 22370 24500 22372
rect 24444 22318 24446 22370
rect 24446 22318 24498 22370
rect 24498 22318 24500 22370
rect 24444 22316 24500 22318
rect 24108 22204 24164 22260
rect 23996 21532 24052 21588
rect 24892 21532 24948 21588
rect 23212 19404 23268 19460
rect 23212 19180 23268 19236
rect 23660 19234 23716 19236
rect 23660 19182 23662 19234
rect 23662 19182 23714 19234
rect 23714 19182 23716 19234
rect 23660 19180 23716 19182
rect 24332 19234 24388 19236
rect 24332 19182 24334 19234
rect 24334 19182 24386 19234
rect 24386 19182 24388 19234
rect 24332 19180 24388 19182
rect 25340 26796 25396 26852
rect 25564 26572 25620 26628
rect 25116 26402 25172 26404
rect 25116 26350 25118 26402
rect 25118 26350 25170 26402
rect 25170 26350 25172 26402
rect 25116 26348 25172 26350
rect 25900 26684 25956 26740
rect 26012 26348 26068 26404
rect 26684 27298 26740 27300
rect 26684 27246 26686 27298
rect 26686 27246 26738 27298
rect 26738 27246 26740 27298
rect 26684 27244 26740 27246
rect 28140 27244 28196 27300
rect 26348 26908 26404 26964
rect 29484 29484 29540 29540
rect 29708 29314 29764 29316
rect 29708 29262 29710 29314
rect 29710 29262 29762 29314
rect 29762 29262 29764 29314
rect 29708 29260 29764 29262
rect 29708 28588 29764 28644
rect 30268 34242 30324 34244
rect 30268 34190 30270 34242
rect 30270 34190 30322 34242
rect 30322 34190 30324 34242
rect 30268 34188 30324 34190
rect 31500 37100 31556 37156
rect 31164 36258 31220 36260
rect 31164 36206 31166 36258
rect 31166 36206 31218 36258
rect 31218 36206 31220 36258
rect 31164 36204 31220 36206
rect 32508 46562 32564 46564
rect 32508 46510 32510 46562
rect 32510 46510 32562 46562
rect 32562 46510 32564 46562
rect 32508 46508 32564 46510
rect 33068 60508 33124 60564
rect 33180 60284 33236 60340
rect 33628 59778 33684 59780
rect 33628 59726 33630 59778
rect 33630 59726 33682 59778
rect 33682 59726 33684 59778
rect 33628 59724 33684 59726
rect 33404 59052 33460 59108
rect 33180 57538 33236 57540
rect 33180 57486 33182 57538
rect 33182 57486 33234 57538
rect 33234 57486 33236 57538
rect 33180 57484 33236 57486
rect 32956 55298 33012 55300
rect 32956 55246 32958 55298
rect 32958 55246 33010 55298
rect 33010 55246 33012 55298
rect 32956 55244 33012 55246
rect 32956 49250 33012 49252
rect 32956 49198 32958 49250
rect 32958 49198 33010 49250
rect 33010 49198 33012 49250
rect 32956 49196 33012 49198
rect 32844 46508 32900 46564
rect 33180 54236 33236 54292
rect 33292 52780 33348 52836
rect 34860 65436 34916 65492
rect 35532 65490 35588 65492
rect 35532 65438 35534 65490
rect 35534 65438 35586 65490
rect 35586 65438 35588 65490
rect 35532 65436 35588 65438
rect 34972 65378 35028 65380
rect 34972 65326 34974 65378
rect 34974 65326 35026 65378
rect 35026 65326 35028 65378
rect 34972 65324 35028 65326
rect 35644 65324 35700 65380
rect 34636 64428 34692 64484
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 37436 65212 37492 65268
rect 38556 65324 38612 65380
rect 36652 64652 36708 64708
rect 37100 64706 37156 64708
rect 37100 64654 37102 64706
rect 37102 64654 37154 64706
rect 37154 64654 37156 64706
rect 37100 64652 37156 64654
rect 38556 64706 38612 64708
rect 38556 64654 38558 64706
rect 38558 64654 38610 64706
rect 38610 64654 38612 64706
rect 38556 64652 38612 64654
rect 39228 64092 39284 64148
rect 45052 66444 45108 66500
rect 43036 66162 43092 66164
rect 43036 66110 43038 66162
rect 43038 66110 43090 66162
rect 43090 66110 43092 66162
rect 43036 66108 43092 66110
rect 46172 66108 46228 66164
rect 41020 65436 41076 65492
rect 42700 65436 42756 65492
rect 41132 65378 41188 65380
rect 41132 65326 41134 65378
rect 41134 65326 41186 65378
rect 41186 65326 41188 65378
rect 41132 65324 41188 65326
rect 40124 65212 40180 65268
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 37884 62466 37940 62468
rect 37884 62414 37886 62466
rect 37886 62414 37938 62466
rect 37938 62414 37940 62466
rect 37884 62412 37940 62414
rect 36316 62300 36372 62356
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 34748 61180 34804 61236
rect 34636 61068 34692 61124
rect 33852 60844 33908 60900
rect 34748 60844 34804 60900
rect 34748 60508 34804 60564
rect 35644 61404 35700 61460
rect 35420 61180 35476 61236
rect 35196 61068 35252 61124
rect 35420 60898 35476 60900
rect 35420 60846 35422 60898
rect 35422 60846 35474 60898
rect 35474 60846 35476 60898
rect 35420 60844 35476 60846
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 36764 62188 36820 62244
rect 36092 61180 36148 61236
rect 35868 61068 35924 61124
rect 36204 59276 36260 59332
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 37212 61458 37268 61460
rect 37212 61406 37214 61458
rect 37214 61406 37266 61458
rect 37266 61406 37268 61458
rect 37212 61404 37268 61406
rect 38332 60956 38388 61012
rect 37548 60844 37604 60900
rect 37772 60786 37828 60788
rect 37772 60734 37774 60786
rect 37774 60734 37826 60786
rect 37826 60734 37828 60786
rect 37772 60732 37828 60734
rect 36988 60508 37044 60564
rect 37324 60674 37380 60676
rect 37324 60622 37326 60674
rect 37326 60622 37378 60674
rect 37378 60622 37380 60674
rect 37324 60620 37380 60622
rect 37212 59330 37268 59332
rect 37212 59278 37214 59330
rect 37214 59278 37266 59330
rect 37266 59278 37268 59330
rect 37212 59276 37268 59278
rect 37996 60674 38052 60676
rect 37996 60622 37998 60674
rect 37998 60622 38050 60674
rect 38050 60622 38052 60674
rect 37996 60620 38052 60622
rect 39116 60898 39172 60900
rect 39116 60846 39118 60898
rect 39118 60846 39170 60898
rect 39170 60846 39172 60898
rect 39116 60844 39172 60846
rect 38668 60620 38724 60676
rect 39004 60620 39060 60676
rect 37324 58940 37380 58996
rect 38108 59724 38164 59780
rect 33740 57484 33796 57540
rect 35980 57708 36036 57764
rect 34972 57372 35028 57428
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 33740 56978 33796 56980
rect 33740 56926 33742 56978
rect 33742 56926 33794 56978
rect 33794 56926 33796 56978
rect 33740 56924 33796 56926
rect 35196 56700 35252 56756
rect 35644 56194 35700 56196
rect 35644 56142 35646 56194
rect 35646 56142 35698 56194
rect 35698 56142 35700 56194
rect 35644 56140 35700 56142
rect 33740 55356 33796 55412
rect 36092 56754 36148 56756
rect 36092 56702 36094 56754
rect 36094 56702 36146 56754
rect 36146 56702 36148 56754
rect 36092 56700 36148 56702
rect 36428 56812 36484 56868
rect 36204 56140 36260 56196
rect 35980 56028 36036 56084
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 55522 35252 55524
rect 35196 55470 35198 55522
rect 35198 55470 35250 55522
rect 35250 55470 35252 55522
rect 35196 55468 35252 55470
rect 35980 55468 36036 55524
rect 37772 58492 37828 58548
rect 37660 57708 37716 57764
rect 37772 57372 37828 57428
rect 37100 56866 37156 56868
rect 37100 56814 37102 56866
rect 37102 56814 37154 56866
rect 37154 56814 37156 56866
rect 37100 56812 37156 56814
rect 37324 56700 37380 56756
rect 37212 56082 37268 56084
rect 37212 56030 37214 56082
rect 37214 56030 37266 56082
rect 37266 56030 37268 56082
rect 37212 56028 37268 56030
rect 36316 55916 36372 55972
rect 34860 55410 34916 55412
rect 34860 55358 34862 55410
rect 34862 55358 34914 55410
rect 34914 55358 34916 55410
rect 34860 55356 34916 55358
rect 33516 52834 33572 52836
rect 33516 52782 33518 52834
rect 33518 52782 33570 52834
rect 33570 52782 33572 52834
rect 33516 52780 33572 52782
rect 33292 52332 33348 52388
rect 33404 52108 33460 52164
rect 33180 49196 33236 49252
rect 33404 49810 33460 49812
rect 33404 49758 33406 49810
rect 33406 49758 33458 49810
rect 33458 49758 33460 49810
rect 33404 49756 33460 49758
rect 33180 45778 33236 45780
rect 33180 45726 33182 45778
rect 33182 45726 33234 45778
rect 33234 45726 33236 45778
rect 33180 45724 33236 45726
rect 32396 44940 32452 44996
rect 32284 44434 32340 44436
rect 32284 44382 32286 44434
rect 32286 44382 32338 44434
rect 32338 44382 32340 44434
rect 32284 44380 32340 44382
rect 32396 44322 32452 44324
rect 32396 44270 32398 44322
rect 32398 44270 32450 44322
rect 32450 44270 32452 44322
rect 32396 44268 32452 44270
rect 33292 44994 33348 44996
rect 33292 44942 33294 44994
rect 33294 44942 33346 44994
rect 33346 44942 33348 44994
rect 33292 44940 33348 44942
rect 33068 44322 33124 44324
rect 33068 44270 33070 44322
rect 33070 44270 33122 44322
rect 33122 44270 33124 44322
rect 33068 44268 33124 44270
rect 33180 43036 33236 43092
rect 32508 41468 32564 41524
rect 32508 41132 32564 41188
rect 33180 41020 33236 41076
rect 32172 39730 32228 39732
rect 32172 39678 32174 39730
rect 32174 39678 32226 39730
rect 32226 39678 32228 39730
rect 32172 39676 32228 39678
rect 32060 39340 32116 39396
rect 31948 38444 32004 38500
rect 31052 34748 31108 34804
rect 30940 34242 30996 34244
rect 30940 34190 30942 34242
rect 30942 34190 30994 34242
rect 30994 34190 30996 34242
rect 30940 34188 30996 34190
rect 30492 31724 30548 31780
rect 31612 34972 31668 35028
rect 31836 34130 31892 34132
rect 31836 34078 31838 34130
rect 31838 34078 31890 34130
rect 31890 34078 31892 34130
rect 31836 34076 31892 34078
rect 31836 33628 31892 33684
rect 31500 33404 31556 33460
rect 31276 33346 31332 33348
rect 31276 33294 31278 33346
rect 31278 33294 31330 33346
rect 31330 33294 31332 33346
rect 31276 33292 31332 33294
rect 31612 33292 31668 33348
rect 31500 31836 31556 31892
rect 31836 32620 31892 32676
rect 31724 32396 31780 32452
rect 30156 30716 30212 30772
rect 30156 30268 30212 30324
rect 31052 31218 31108 31220
rect 31052 31166 31054 31218
rect 31054 31166 31106 31218
rect 31106 31166 31108 31218
rect 31052 31164 31108 31166
rect 33404 41468 33460 41524
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 37996 56866 38052 56868
rect 37996 56814 37998 56866
rect 37998 56814 38050 56866
rect 38050 56814 38052 56866
rect 37996 56812 38052 56814
rect 34524 53730 34580 53732
rect 34524 53678 34526 53730
rect 34526 53678 34578 53730
rect 34578 53678 34580 53730
rect 34524 53676 34580 53678
rect 35980 53116 36036 53172
rect 35644 53004 35700 53060
rect 34412 52946 34468 52948
rect 34412 52894 34414 52946
rect 34414 52894 34466 52946
rect 34466 52894 34468 52946
rect 34412 52892 34468 52894
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 33740 52220 33796 52276
rect 35980 52946 36036 52948
rect 35980 52894 35982 52946
rect 35982 52894 36034 52946
rect 36034 52894 36036 52946
rect 35980 52892 36036 52894
rect 36204 53788 36260 53844
rect 37100 53842 37156 53844
rect 37100 53790 37102 53842
rect 37102 53790 37154 53842
rect 37154 53790 37156 53842
rect 37100 53788 37156 53790
rect 37996 53788 38052 53844
rect 36428 53676 36484 53732
rect 36316 53116 36372 53172
rect 35644 52162 35700 52164
rect 35644 52110 35646 52162
rect 35646 52110 35698 52162
rect 35698 52110 35700 52162
rect 35644 52108 35700 52110
rect 37324 53116 37380 53172
rect 36652 53058 36708 53060
rect 36652 53006 36654 53058
rect 36654 53006 36706 53058
rect 36706 53006 36708 53058
rect 36652 53004 36708 53006
rect 36764 52946 36820 52948
rect 36764 52894 36766 52946
rect 36766 52894 36818 52946
rect 36818 52894 36820 52946
rect 36764 52892 36820 52894
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 34188 49756 34244 49812
rect 36764 51212 36820 51268
rect 37772 51266 37828 51268
rect 37772 51214 37774 51266
rect 37774 51214 37826 51266
rect 37826 51214 37828 51266
rect 37772 51212 37828 51214
rect 39228 59052 39284 59108
rect 39004 58940 39060 58996
rect 38556 58492 38612 58548
rect 38220 56700 38276 56756
rect 39004 56082 39060 56084
rect 39004 56030 39006 56082
rect 39006 56030 39058 56082
rect 39058 56030 39060 56082
rect 39004 56028 39060 56030
rect 38332 55186 38388 55188
rect 38332 55134 38334 55186
rect 38334 55134 38386 55186
rect 38386 55134 38388 55186
rect 38332 55132 38388 55134
rect 38556 53452 38612 53508
rect 38556 51212 38612 51268
rect 35084 49810 35140 49812
rect 35084 49758 35086 49810
rect 35086 49758 35138 49810
rect 35138 49758 35140 49810
rect 35084 49756 35140 49758
rect 34860 49420 34916 49476
rect 37660 49922 37716 49924
rect 37660 49870 37662 49922
rect 37662 49870 37714 49922
rect 37714 49870 37716 49922
rect 37660 49868 37716 49870
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 33740 49196 33796 49252
rect 35084 48748 35140 48804
rect 34636 47404 34692 47460
rect 34748 46844 34804 46900
rect 34972 47404 35028 47460
rect 34412 45276 34468 45332
rect 34076 45164 34132 45220
rect 33964 44940 34020 44996
rect 33740 44322 33796 44324
rect 33740 44270 33742 44322
rect 33742 44270 33794 44322
rect 33794 44270 33796 44322
rect 33740 44268 33796 44270
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35420 47682 35476 47684
rect 35420 47630 35422 47682
rect 35422 47630 35474 47682
rect 35474 47630 35476 47682
rect 35420 47628 35476 47630
rect 36652 47628 36708 47684
rect 36428 47404 36484 47460
rect 36092 47068 36148 47124
rect 37436 47628 37492 47684
rect 37996 47570 38052 47572
rect 37996 47518 37998 47570
rect 37998 47518 38050 47570
rect 38050 47518 38052 47570
rect 37996 47516 38052 47518
rect 37100 47180 37156 47236
rect 37660 47180 37716 47236
rect 35868 46620 35924 46676
rect 36652 46674 36708 46676
rect 36652 46622 36654 46674
rect 36654 46622 36706 46674
rect 36706 46622 36708 46674
rect 36652 46620 36708 46622
rect 37436 46620 37492 46676
rect 35756 46396 35812 46452
rect 36316 46450 36372 46452
rect 36316 46398 36318 46450
rect 36318 46398 36370 46450
rect 36370 46398 36372 46450
rect 36316 46396 36372 46398
rect 37100 46396 37156 46452
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 36204 45276 36260 45332
rect 36652 45330 36708 45332
rect 36652 45278 36654 45330
rect 36654 45278 36706 45330
rect 36706 45278 36708 45330
rect 36652 45276 36708 45278
rect 35420 44994 35476 44996
rect 35420 44942 35422 44994
rect 35422 44942 35474 44994
rect 35474 44942 35476 44994
rect 35420 44940 35476 44942
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34076 44210 34132 44212
rect 34076 44158 34078 44210
rect 34078 44158 34130 44210
rect 34130 44158 34132 44210
rect 34076 44156 34132 44158
rect 34636 44098 34692 44100
rect 34636 44046 34638 44098
rect 34638 44046 34690 44098
rect 34690 44046 34692 44098
rect 34636 44044 34692 44046
rect 34860 44098 34916 44100
rect 34860 44046 34862 44098
rect 34862 44046 34914 44098
rect 34914 44046 34916 44098
rect 34860 44044 34916 44046
rect 35644 43820 35700 43876
rect 36764 43932 36820 43988
rect 33740 43484 33796 43540
rect 33740 42028 33796 42084
rect 33740 41746 33796 41748
rect 33740 41694 33742 41746
rect 33742 41694 33794 41746
rect 33794 41694 33796 41746
rect 33740 41692 33796 41694
rect 33628 41468 33684 41524
rect 33516 41186 33572 41188
rect 33516 41134 33518 41186
rect 33518 41134 33570 41186
rect 33570 41134 33572 41186
rect 33516 41132 33572 41134
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36428 42140 36484 42196
rect 34076 42082 34132 42084
rect 34076 42030 34078 42082
rect 34078 42030 34130 42082
rect 34130 42030 34132 42082
rect 34076 42028 34132 42030
rect 35532 42082 35588 42084
rect 35532 42030 35534 42082
rect 35534 42030 35586 42082
rect 35586 42030 35588 42082
rect 35532 42028 35588 42030
rect 34412 41468 34468 41524
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 32060 36204 32116 36260
rect 33068 36988 33124 37044
rect 32172 35532 32228 35588
rect 32060 31778 32116 31780
rect 32060 31726 32062 31778
rect 32062 31726 32114 31778
rect 32114 31726 32116 31778
rect 32060 31724 32116 31726
rect 32508 35698 32564 35700
rect 32508 35646 32510 35698
rect 32510 35646 32562 35698
rect 32562 35646 32564 35698
rect 32508 35644 32564 35646
rect 32956 33628 33012 33684
rect 32284 32620 32340 32676
rect 32284 32060 32340 32116
rect 33068 31836 33124 31892
rect 32060 31218 32116 31220
rect 32060 31166 32062 31218
rect 32062 31166 32114 31218
rect 32114 31166 32116 31218
rect 32060 31164 32116 31166
rect 32284 30156 32340 30212
rect 30492 30098 30548 30100
rect 30492 30046 30494 30098
rect 30494 30046 30546 30098
rect 30546 30046 30548 30098
rect 30492 30044 30548 30046
rect 29932 29986 29988 29988
rect 29932 29934 29934 29986
rect 29934 29934 29986 29986
rect 29986 29934 29988 29986
rect 29932 29932 29988 29934
rect 31276 30098 31332 30100
rect 31276 30046 31278 30098
rect 31278 30046 31330 30098
rect 31330 30046 31332 30098
rect 31276 30044 31332 30046
rect 30604 29932 30660 29988
rect 31388 29986 31444 29988
rect 31388 29934 31390 29986
rect 31390 29934 31442 29986
rect 31442 29934 31444 29986
rect 31388 29932 31444 29934
rect 30828 29650 30884 29652
rect 30828 29598 30830 29650
rect 30830 29598 30882 29650
rect 30882 29598 30884 29650
rect 30828 29596 30884 29598
rect 31836 29650 31892 29652
rect 31836 29598 31838 29650
rect 31838 29598 31890 29650
rect 31890 29598 31892 29650
rect 31836 29596 31892 29598
rect 31164 29538 31220 29540
rect 31164 29486 31166 29538
rect 31166 29486 31218 29538
rect 31218 29486 31220 29538
rect 31164 29484 31220 29486
rect 31276 29036 31332 29092
rect 30604 28812 30660 28868
rect 30380 28700 30436 28756
rect 30268 28642 30324 28644
rect 30268 28590 30270 28642
rect 30270 28590 30322 28642
rect 30322 28590 30324 28642
rect 30268 28588 30324 28590
rect 30716 28530 30772 28532
rect 30716 28478 30718 28530
rect 30718 28478 30770 28530
rect 30770 28478 30772 28530
rect 30716 28476 30772 28478
rect 26684 26850 26740 26852
rect 26684 26798 26686 26850
rect 26686 26798 26738 26850
rect 26738 26798 26740 26850
rect 26684 26796 26740 26798
rect 27020 26796 27076 26852
rect 26124 25900 26180 25956
rect 26236 26012 26292 26068
rect 25900 25676 25956 25732
rect 26012 25564 26068 25620
rect 26348 25900 26404 25956
rect 26572 26290 26628 26292
rect 26572 26238 26574 26290
rect 26574 26238 26626 26290
rect 26626 26238 26628 26290
rect 26572 26236 26628 26238
rect 26460 25564 26516 25620
rect 26908 26124 26964 26180
rect 26908 25676 26964 25732
rect 26236 25282 26292 25284
rect 26236 25230 26238 25282
rect 26238 25230 26290 25282
rect 26290 25230 26292 25282
rect 26236 25228 26292 25230
rect 25452 25004 25508 25060
rect 25228 24722 25284 24724
rect 25228 24670 25230 24722
rect 25230 24670 25282 24722
rect 25282 24670 25284 24722
rect 25228 24668 25284 24670
rect 25116 23660 25172 23716
rect 25340 23772 25396 23828
rect 25340 23436 25396 23492
rect 25228 22204 25284 22260
rect 26684 25004 26740 25060
rect 25564 24946 25620 24948
rect 25564 24894 25566 24946
rect 25566 24894 25618 24946
rect 25618 24894 25620 24946
rect 25564 24892 25620 24894
rect 26348 24892 26404 24948
rect 26348 24444 26404 24500
rect 25788 23436 25844 23492
rect 25900 22316 25956 22372
rect 25340 21810 25396 21812
rect 25340 21758 25342 21810
rect 25342 21758 25394 21810
rect 25394 21758 25396 21810
rect 25340 21756 25396 21758
rect 28588 26460 28644 26516
rect 29708 28028 29764 28084
rect 27468 26348 27524 26404
rect 28812 26402 28868 26404
rect 28812 26350 28814 26402
rect 28814 26350 28866 26402
rect 28866 26350 28868 26402
rect 28812 26348 28868 26350
rect 28252 26290 28308 26292
rect 28252 26238 28254 26290
rect 28254 26238 28306 26290
rect 28306 26238 28308 26290
rect 28252 26236 28308 26238
rect 28588 26290 28644 26292
rect 28588 26238 28590 26290
rect 28590 26238 28642 26290
rect 28642 26238 28644 26290
rect 28588 26236 28644 26238
rect 27132 25564 27188 25620
rect 27244 25452 27300 25508
rect 27580 25788 27636 25844
rect 27692 25730 27748 25732
rect 27692 25678 27694 25730
rect 27694 25678 27746 25730
rect 27746 25678 27748 25730
rect 27692 25676 27748 25678
rect 27804 25618 27860 25620
rect 27804 25566 27806 25618
rect 27806 25566 27858 25618
rect 27858 25566 27860 25618
rect 27804 25564 27860 25566
rect 27692 25452 27748 25508
rect 28140 25564 28196 25620
rect 28028 25340 28084 25396
rect 27692 24834 27748 24836
rect 27692 24782 27694 24834
rect 27694 24782 27746 24834
rect 27746 24782 27748 24834
rect 27692 24780 27748 24782
rect 27468 24722 27524 24724
rect 27468 24670 27470 24722
rect 27470 24670 27522 24722
rect 27522 24670 27524 24722
rect 27468 24668 27524 24670
rect 27132 24498 27188 24500
rect 27132 24446 27134 24498
rect 27134 24446 27186 24498
rect 27186 24446 27188 24498
rect 27132 24444 27188 24446
rect 26796 23436 26852 23492
rect 26908 23548 26964 23604
rect 27580 23378 27636 23380
rect 27580 23326 27582 23378
rect 27582 23326 27634 23378
rect 27634 23326 27636 23378
rect 27580 23324 27636 23326
rect 29148 26290 29204 26292
rect 29148 26238 29150 26290
rect 29150 26238 29202 26290
rect 29202 26238 29204 26290
rect 29148 26236 29204 26238
rect 28588 25618 28644 25620
rect 28588 25566 28590 25618
rect 28590 25566 28642 25618
rect 28642 25566 28644 25618
rect 28588 25564 28644 25566
rect 28140 24668 28196 24724
rect 28252 23884 28308 23940
rect 27916 23436 27972 23492
rect 27804 22204 27860 22260
rect 29596 26460 29652 26516
rect 29372 26236 29428 26292
rect 31164 28642 31220 28644
rect 31164 28590 31166 28642
rect 31166 28590 31218 28642
rect 31218 28590 31220 28642
rect 31164 28588 31220 28590
rect 31052 27970 31108 27972
rect 31052 27918 31054 27970
rect 31054 27918 31106 27970
rect 31106 27918 31108 27970
rect 31052 27916 31108 27918
rect 30268 26514 30324 26516
rect 30268 26462 30270 26514
rect 30270 26462 30322 26514
rect 30322 26462 30324 26514
rect 30268 26460 30324 26462
rect 30828 26514 30884 26516
rect 30828 26462 30830 26514
rect 30830 26462 30882 26514
rect 30882 26462 30884 26514
rect 30828 26460 30884 26462
rect 28924 25564 28980 25620
rect 29148 25506 29204 25508
rect 29148 25454 29150 25506
rect 29150 25454 29202 25506
rect 29202 25454 29204 25506
rect 29148 25452 29204 25454
rect 28924 25228 28980 25284
rect 29484 25116 29540 25172
rect 28924 24834 28980 24836
rect 28924 24782 28926 24834
rect 28926 24782 28978 24834
rect 28978 24782 28980 24834
rect 28924 24780 28980 24782
rect 29148 24556 29204 24612
rect 29260 23714 29316 23716
rect 29260 23662 29262 23714
rect 29262 23662 29314 23714
rect 29314 23662 29316 23714
rect 29260 23660 29316 23662
rect 28812 23100 28868 23156
rect 28476 21756 28532 21812
rect 29372 20860 29428 20916
rect 26796 20130 26852 20132
rect 26796 20078 26798 20130
rect 26798 20078 26850 20130
rect 26850 20078 26852 20130
rect 26796 20076 26852 20078
rect 26572 20018 26628 20020
rect 26572 19966 26574 20018
rect 26574 19966 26626 20018
rect 26626 19966 26628 20018
rect 26572 19964 26628 19966
rect 26236 19346 26292 19348
rect 26236 19294 26238 19346
rect 26238 19294 26290 19346
rect 26290 19294 26292 19346
rect 26236 19292 26292 19294
rect 25004 19180 25060 19236
rect 27244 20018 27300 20020
rect 27244 19966 27246 20018
rect 27246 19966 27298 20018
rect 27298 19966 27300 20018
rect 27244 19964 27300 19966
rect 26796 19292 26852 19348
rect 23100 18396 23156 18452
rect 22764 17554 22820 17556
rect 22764 17502 22766 17554
rect 22766 17502 22818 17554
rect 22818 17502 22820 17554
rect 22764 17500 22820 17502
rect 24220 18508 24276 18564
rect 23772 18338 23828 18340
rect 23772 18286 23774 18338
rect 23774 18286 23826 18338
rect 23826 18286 23828 18338
rect 23772 18284 23828 18286
rect 24444 18284 24500 18340
rect 24444 17612 24500 17668
rect 25004 18060 25060 18116
rect 20412 16156 20468 16212
rect 21868 16156 21924 16212
rect 19292 15986 19348 15988
rect 19292 15934 19294 15986
rect 19294 15934 19346 15986
rect 19346 15934 19348 15986
rect 19292 15932 19348 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 22428 16210 22484 16212
rect 22428 16158 22430 16210
rect 22430 16158 22482 16210
rect 22482 16158 22484 16210
rect 22428 16156 22484 16158
rect 19068 14476 19124 14532
rect 18732 13858 18788 13860
rect 18732 13806 18734 13858
rect 18734 13806 18786 13858
rect 18786 13806 18788 13858
rect 18732 13804 18788 13806
rect 18844 13746 18900 13748
rect 18844 13694 18846 13746
rect 18846 13694 18898 13746
rect 18898 13694 18900 13746
rect 18844 13692 18900 13694
rect 18956 13468 19012 13524
rect 18732 12850 18788 12852
rect 18732 12798 18734 12850
rect 18734 12798 18786 12850
rect 18786 12798 18788 12850
rect 18732 12796 18788 12798
rect 18732 11452 18788 11508
rect 19180 12850 19236 12852
rect 19180 12798 19182 12850
rect 19182 12798 19234 12850
rect 19234 12798 19236 12850
rect 19180 12796 19236 12798
rect 18956 11676 19012 11732
rect 18844 11340 18900 11396
rect 18956 11282 19012 11284
rect 18956 11230 18958 11282
rect 18958 11230 19010 11282
rect 19010 11230 19012 11282
rect 18956 11228 19012 11230
rect 18844 11170 18900 11172
rect 18844 11118 18846 11170
rect 18846 11118 18898 11170
rect 18898 11118 18900 11170
rect 18844 11116 18900 11118
rect 18396 10722 18452 10724
rect 18396 10670 18398 10722
rect 18398 10670 18450 10722
rect 18450 10670 18452 10722
rect 18396 10668 18452 10670
rect 22764 16156 22820 16212
rect 22988 15874 23044 15876
rect 22988 15822 22990 15874
rect 22990 15822 23042 15874
rect 23042 15822 23044 15874
rect 22988 15820 23044 15822
rect 22652 14812 22708 14868
rect 22428 14476 22484 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20748 13970 20804 13972
rect 20748 13918 20750 13970
rect 20750 13918 20802 13970
rect 20802 13918 20804 13970
rect 20748 13916 20804 13918
rect 19852 13804 19908 13860
rect 21084 13804 21140 13860
rect 19404 13468 19460 13524
rect 19852 13356 19908 13412
rect 19404 12738 19460 12740
rect 19404 12686 19406 12738
rect 19406 12686 19458 12738
rect 19458 12686 19460 12738
rect 19404 12684 19460 12686
rect 20412 13522 20468 13524
rect 20412 13470 20414 13522
rect 20414 13470 20466 13522
rect 20466 13470 20468 13522
rect 20412 13468 20468 13470
rect 20076 13132 20132 13188
rect 20300 13356 20356 13412
rect 20188 13020 20244 13076
rect 21196 13468 21252 13524
rect 20860 13020 20916 13076
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 22092 13804 22148 13860
rect 21756 13746 21812 13748
rect 21756 13694 21758 13746
rect 21758 13694 21810 13746
rect 21810 13694 21812 13746
rect 21756 13692 21812 13694
rect 21644 12796 21700 12852
rect 21196 11900 21252 11956
rect 21308 11676 21364 11732
rect 20188 11170 20244 11172
rect 20188 11118 20190 11170
rect 20190 11118 20242 11170
rect 20242 11118 20244 11170
rect 20188 11116 20244 11118
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19292 10780 19348 10836
rect 19180 10556 19236 10612
rect 22204 13692 22260 13748
rect 22652 13858 22708 13860
rect 22652 13806 22654 13858
rect 22654 13806 22706 13858
rect 22706 13806 22708 13858
rect 22652 13804 22708 13806
rect 23660 15820 23716 15876
rect 23212 14588 23268 14644
rect 23100 13692 23156 13748
rect 23212 13580 23268 13636
rect 23324 13804 23380 13860
rect 22540 12962 22596 12964
rect 22540 12910 22542 12962
rect 22542 12910 22594 12962
rect 22594 12910 22596 12962
rect 22540 12908 22596 12910
rect 22428 12850 22484 12852
rect 22428 12798 22430 12850
rect 22430 12798 22482 12850
rect 22482 12798 22484 12850
rect 22428 12796 22484 12798
rect 22652 11676 22708 11732
rect 24780 15708 24836 15764
rect 24332 14252 24388 14308
rect 23548 13468 23604 13524
rect 23772 13186 23828 13188
rect 23772 13134 23774 13186
rect 23774 13134 23826 13186
rect 23826 13134 23828 13186
rect 23772 13132 23828 13134
rect 24220 12962 24276 12964
rect 24220 12910 24222 12962
rect 24222 12910 24274 12962
rect 24274 12910 24276 12962
rect 24220 12908 24276 12910
rect 24668 13468 24724 13524
rect 24556 13132 24612 13188
rect 21980 11228 22036 11284
rect 21532 10668 21588 10724
rect 17948 9660 18004 9716
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 15484 6690 15540 6692
rect 15484 6638 15486 6690
rect 15486 6638 15538 6690
rect 15538 6638 15540 6690
rect 15484 6636 15540 6638
rect 18844 9996 18900 10052
rect 18620 9938 18676 9940
rect 18620 9886 18622 9938
rect 18622 9886 18674 9938
rect 18674 9886 18676 9938
rect 18620 9884 18676 9886
rect 19404 9826 19460 9828
rect 19404 9774 19406 9826
rect 19406 9774 19458 9826
rect 19458 9774 19460 9826
rect 19404 9772 19460 9774
rect 18620 9714 18676 9716
rect 18620 9662 18622 9714
rect 18622 9662 18674 9714
rect 18674 9662 18676 9714
rect 18620 9660 18676 9662
rect 18956 9660 19012 9716
rect 19068 9602 19124 9604
rect 19068 9550 19070 9602
rect 19070 9550 19122 9602
rect 19122 9550 19124 9602
rect 19068 9548 19124 9550
rect 19068 9324 19124 9380
rect 19516 9324 19572 9380
rect 18172 9100 18228 9156
rect 18956 9154 19012 9156
rect 18956 9102 18958 9154
rect 18958 9102 19010 9154
rect 19010 9102 19012 9154
rect 18956 9100 19012 9102
rect 19404 9100 19460 9156
rect 18844 7868 18900 7924
rect 17500 6636 17556 6692
rect 17724 6748 17780 6804
rect 16156 6578 16212 6580
rect 16156 6526 16158 6578
rect 16158 6526 16210 6578
rect 16210 6526 16212 6578
rect 16156 6524 16212 6526
rect 17388 6524 17444 6580
rect 18620 6802 18676 6804
rect 18620 6750 18622 6802
rect 18622 6750 18674 6802
rect 18674 6750 18676 6802
rect 18620 6748 18676 6750
rect 18508 6636 18564 6692
rect 19292 7586 19348 7588
rect 19292 7534 19294 7586
rect 19294 7534 19346 7586
rect 19346 7534 19348 7586
rect 19292 7532 19348 7534
rect 18956 7474 19012 7476
rect 18956 7422 18958 7474
rect 18958 7422 19010 7474
rect 19010 7422 19012 7474
rect 18956 7420 19012 7422
rect 18844 7196 18900 7252
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19068 6972 19124 7028
rect 18956 6578 19012 6580
rect 18956 6526 18958 6578
rect 18958 6526 19010 6578
rect 19010 6526 19012 6578
rect 18956 6524 19012 6526
rect 19964 10108 20020 10164
rect 19852 9660 19908 9716
rect 21420 9602 21476 9604
rect 21420 9550 21422 9602
rect 21422 9550 21474 9602
rect 21474 9550 21476 9602
rect 21420 9548 21476 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 7868 19684 7924
rect 21644 10332 21700 10388
rect 23324 12460 23380 12516
rect 24780 12962 24836 12964
rect 24780 12910 24782 12962
rect 24782 12910 24834 12962
rect 24834 12910 24836 12962
rect 24780 12908 24836 12910
rect 22764 10332 22820 10388
rect 21756 9884 21812 9940
rect 22204 9938 22260 9940
rect 22204 9886 22206 9938
rect 22206 9886 22258 9938
rect 22258 9886 22260 9938
rect 22204 9884 22260 9886
rect 23436 9714 23492 9716
rect 23436 9662 23438 9714
rect 23438 9662 23490 9714
rect 23490 9662 23492 9714
rect 23436 9660 23492 9662
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19964 7250 20020 7252
rect 19964 7198 19966 7250
rect 19966 7198 20018 7250
rect 20018 7198 20020 7250
rect 19964 7196 20020 7198
rect 21084 7362 21140 7364
rect 21084 7310 21086 7362
rect 21086 7310 21138 7362
rect 21138 7310 21140 7362
rect 21084 7308 21140 7310
rect 20748 7250 20804 7252
rect 20748 7198 20750 7250
rect 20750 7198 20802 7250
rect 20802 7198 20804 7250
rect 20748 7196 20804 7198
rect 20188 6972 20244 7028
rect 20524 6972 20580 7028
rect 20188 6748 20244 6804
rect 19404 6636 19460 6692
rect 19292 6412 19348 6468
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18508 5180 18564 5236
rect 20300 6636 20356 6692
rect 20636 6690 20692 6692
rect 20636 6638 20638 6690
rect 20638 6638 20690 6690
rect 20690 6638 20692 6690
rect 20636 6636 20692 6638
rect 20300 6300 20356 6356
rect 22428 8428 22484 8484
rect 21532 7532 21588 7588
rect 21308 7084 21364 7140
rect 21420 7196 21476 7252
rect 21308 6690 21364 6692
rect 21308 6638 21310 6690
rect 21310 6638 21362 6690
rect 21362 6638 21364 6690
rect 21308 6636 21364 6638
rect 21196 6412 21252 6468
rect 20748 6076 20804 6132
rect 21644 7308 21700 7364
rect 22764 7084 22820 7140
rect 23548 7084 23604 7140
rect 22204 6802 22260 6804
rect 22204 6750 22206 6802
rect 22206 6750 22258 6802
rect 22258 6750 22260 6802
rect 22204 6748 22260 6750
rect 23212 6748 23268 6804
rect 21980 6578 22036 6580
rect 21980 6526 21982 6578
rect 21982 6526 22034 6578
rect 22034 6526 22036 6578
rect 21980 6524 22036 6526
rect 21756 6466 21812 6468
rect 21756 6414 21758 6466
rect 21758 6414 21810 6466
rect 21810 6414 21812 6466
rect 21756 6412 21812 6414
rect 22316 6412 22372 6468
rect 21644 6130 21700 6132
rect 21644 6078 21646 6130
rect 21646 6078 21698 6130
rect 21698 6078 21700 6130
rect 21644 6076 21700 6078
rect 21756 5906 21812 5908
rect 21756 5854 21758 5906
rect 21758 5854 21810 5906
rect 21810 5854 21812 5906
rect 21756 5852 21812 5854
rect 21308 5740 21364 5796
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22092 5740 22148 5796
rect 21420 5234 21476 5236
rect 21420 5182 21422 5234
rect 21422 5182 21474 5234
rect 21474 5182 21476 5234
rect 21420 5180 21476 5182
rect 23324 6636 23380 6692
rect 23660 6412 23716 6468
rect 23772 7308 23828 7364
rect 23884 6972 23940 7028
rect 23884 6466 23940 6468
rect 23884 6414 23886 6466
rect 23886 6414 23938 6466
rect 23938 6414 23940 6466
rect 23884 6412 23940 6414
rect 24556 10610 24612 10612
rect 24556 10558 24558 10610
rect 24558 10558 24610 10610
rect 24610 10558 24612 10610
rect 24556 10556 24612 10558
rect 24668 10108 24724 10164
rect 27468 18620 27524 18676
rect 27692 20076 27748 20132
rect 27132 18396 27188 18452
rect 25340 17388 25396 17444
rect 27580 17106 27636 17108
rect 27580 17054 27582 17106
rect 27582 17054 27634 17106
rect 27634 17054 27636 17106
rect 27580 17052 27636 17054
rect 30268 26066 30324 26068
rect 30268 26014 30270 26066
rect 30270 26014 30322 26066
rect 30322 26014 30324 26066
rect 30268 26012 30324 26014
rect 30156 25452 30212 25508
rect 31388 27916 31444 27972
rect 31836 28476 31892 28532
rect 31500 27858 31556 27860
rect 31500 27806 31502 27858
rect 31502 27806 31554 27858
rect 31554 27806 31556 27858
rect 31500 27804 31556 27806
rect 32060 27970 32116 27972
rect 32060 27918 32062 27970
rect 32062 27918 32114 27970
rect 32114 27918 32116 27970
rect 32060 27916 32116 27918
rect 31836 26460 31892 26516
rect 29932 25116 29988 25172
rect 33516 37266 33572 37268
rect 33516 37214 33518 37266
rect 33518 37214 33570 37266
rect 33570 37214 33572 37266
rect 33516 37212 33572 37214
rect 33292 36092 33348 36148
rect 33628 34076 33684 34132
rect 34188 41020 34244 41076
rect 34748 41074 34804 41076
rect 34748 41022 34750 41074
rect 34750 41022 34802 41074
rect 34802 41022 34804 41074
rect 34748 41020 34804 41022
rect 34076 38444 34132 38500
rect 33964 37884 34020 37940
rect 34300 37212 34356 37268
rect 34412 37324 34468 37380
rect 34076 37154 34132 37156
rect 34076 37102 34078 37154
rect 34078 37102 34130 37154
rect 34130 37102 34132 37154
rect 34076 37100 34132 37102
rect 33964 35644 34020 35700
rect 33852 33292 33908 33348
rect 34188 35586 34244 35588
rect 34188 35534 34190 35586
rect 34190 35534 34242 35586
rect 34242 35534 34244 35586
rect 34188 35532 34244 35534
rect 34412 33964 34468 34020
rect 34524 37772 34580 37828
rect 35084 40962 35140 40964
rect 35084 40910 35086 40962
rect 35086 40910 35138 40962
rect 35138 40910 35140 40962
rect 35084 40908 35140 40910
rect 34972 40460 35028 40516
rect 35644 40908 35700 40964
rect 36092 41186 36148 41188
rect 36092 41134 36094 41186
rect 36094 41134 36146 41186
rect 36146 41134 36148 41186
rect 36092 41132 36148 41134
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 39730 35252 39732
rect 35196 39678 35198 39730
rect 35198 39678 35250 39730
rect 35250 39678 35252 39730
rect 35196 39676 35252 39678
rect 34636 37324 34692 37380
rect 34748 38668 34804 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 37660 46620 37716 46676
rect 37548 46508 37604 46564
rect 37548 45890 37604 45892
rect 37548 45838 37550 45890
rect 37550 45838 37602 45890
rect 37602 45838 37604 45890
rect 37548 45836 37604 45838
rect 38556 49868 38612 49924
rect 39452 62524 39508 62580
rect 41580 64146 41636 64148
rect 41580 64094 41582 64146
rect 41582 64094 41634 64146
rect 41634 64094 41636 64146
rect 41580 64092 41636 64094
rect 41020 63026 41076 63028
rect 41020 62974 41022 63026
rect 41022 62974 41074 63026
rect 41074 62974 41076 63026
rect 41020 62972 41076 62974
rect 42028 65324 42084 65380
rect 41804 62972 41860 63028
rect 41916 62860 41972 62916
rect 41244 62354 41300 62356
rect 41244 62302 41246 62354
rect 41246 62302 41298 62354
rect 41298 62302 41300 62354
rect 41244 62300 41300 62302
rect 41020 62242 41076 62244
rect 41020 62190 41022 62242
rect 41022 62190 41074 62242
rect 41074 62190 41076 62242
rect 41020 62188 41076 62190
rect 39452 58940 39508 58996
rect 39564 55132 39620 55188
rect 42028 61404 42084 61460
rect 41020 61292 41076 61348
rect 39900 60786 39956 60788
rect 39900 60734 39902 60786
rect 39902 60734 39954 60786
rect 39954 60734 39956 60786
rect 39900 60732 39956 60734
rect 40236 60732 40292 60788
rect 39900 60508 39956 60564
rect 40236 60002 40292 60004
rect 40236 59950 40238 60002
rect 40238 59950 40290 60002
rect 40290 59950 40292 60002
rect 40236 59948 40292 59950
rect 39452 54626 39508 54628
rect 39452 54574 39454 54626
rect 39454 54574 39506 54626
rect 39506 54574 39508 54626
rect 39452 54572 39508 54574
rect 39564 53676 39620 53732
rect 39452 53564 39508 53620
rect 40012 53340 40068 53396
rect 40796 59778 40852 59780
rect 40796 59726 40798 59778
rect 40798 59726 40850 59778
rect 40850 59726 40852 59778
rect 40796 59724 40852 59726
rect 40684 59500 40740 59556
rect 41020 59106 41076 59108
rect 41020 59054 41022 59106
rect 41022 59054 41074 59106
rect 41074 59054 41076 59106
rect 41020 59052 41076 59054
rect 41020 58492 41076 58548
rect 40460 55020 40516 55076
rect 40796 54572 40852 54628
rect 41020 54012 41076 54068
rect 41244 59500 41300 59556
rect 41244 59218 41300 59220
rect 41244 59166 41246 59218
rect 41246 59166 41298 59218
rect 41298 59166 41300 59218
rect 41244 59164 41300 59166
rect 41468 60562 41524 60564
rect 41468 60510 41470 60562
rect 41470 60510 41522 60562
rect 41522 60510 41524 60562
rect 41468 60508 41524 60510
rect 41916 60508 41972 60564
rect 41468 59724 41524 59780
rect 41804 59388 41860 59444
rect 43372 63922 43428 63924
rect 43372 63870 43374 63922
rect 43374 63870 43426 63922
rect 43426 63870 43428 63922
rect 43372 63868 43428 63870
rect 44380 65324 44436 65380
rect 44940 64092 44996 64148
rect 44828 63980 44884 64036
rect 42252 62188 42308 62244
rect 42924 62914 42980 62916
rect 42924 62862 42926 62914
rect 42926 62862 42978 62914
rect 42978 62862 42980 62914
rect 42924 62860 42980 62862
rect 43820 63922 43876 63924
rect 43820 63870 43822 63922
rect 43822 63870 43874 63922
rect 43874 63870 43876 63922
rect 43820 63868 43876 63870
rect 43484 63138 43540 63140
rect 43484 63086 43486 63138
rect 43486 63086 43538 63138
rect 43538 63086 43540 63138
rect 43484 63084 43540 63086
rect 42700 62300 42756 62356
rect 43484 62354 43540 62356
rect 43484 62302 43486 62354
rect 43486 62302 43538 62354
rect 43538 62302 43540 62354
rect 43484 62300 43540 62302
rect 43596 62188 43652 62244
rect 43708 61458 43764 61460
rect 43708 61406 43710 61458
rect 43710 61406 43762 61458
rect 43762 61406 43764 61458
rect 43708 61404 43764 61406
rect 42476 60508 42532 60564
rect 42364 59330 42420 59332
rect 42364 59278 42366 59330
rect 42366 59278 42418 59330
rect 42418 59278 42420 59330
rect 42364 59276 42420 59278
rect 41916 58940 41972 58996
rect 41804 58546 41860 58548
rect 41804 58494 41806 58546
rect 41806 58494 41858 58546
rect 41858 58494 41860 58546
rect 41804 58492 41860 58494
rect 42812 59388 42868 59444
rect 43036 59330 43092 59332
rect 43036 59278 43038 59330
rect 43038 59278 43090 59330
rect 43090 59278 43092 59330
rect 43036 59276 43092 59278
rect 42364 58492 42420 58548
rect 43260 59218 43316 59220
rect 43260 59166 43262 59218
rect 43262 59166 43314 59218
rect 43314 59166 43316 59218
rect 43260 59164 43316 59166
rect 44044 63138 44100 63140
rect 44044 63086 44046 63138
rect 44046 63086 44098 63138
rect 44098 63086 44100 63138
rect 44044 63084 44100 63086
rect 44156 63026 44212 63028
rect 44156 62974 44158 63026
rect 44158 62974 44210 63026
rect 44210 62974 44212 63026
rect 44156 62972 44212 62974
rect 43932 62354 43988 62356
rect 43932 62302 43934 62354
rect 43934 62302 43986 62354
rect 43986 62302 43988 62354
rect 43932 62300 43988 62302
rect 45164 63868 45220 63924
rect 45612 64204 45668 64260
rect 44940 63138 44996 63140
rect 44940 63086 44942 63138
rect 44942 63086 44994 63138
rect 44994 63086 44996 63138
rect 44940 63084 44996 63086
rect 45052 63026 45108 63028
rect 45052 62974 45054 63026
rect 45054 62974 45106 63026
rect 45106 62974 45108 63026
rect 45052 62972 45108 62974
rect 45276 62914 45332 62916
rect 45276 62862 45278 62914
rect 45278 62862 45330 62914
rect 45330 62862 45332 62914
rect 45276 62860 45332 62862
rect 45276 62412 45332 62468
rect 44940 62354 44996 62356
rect 44940 62302 44942 62354
rect 44942 62302 44994 62354
rect 44994 62302 44996 62354
rect 44940 62300 44996 62302
rect 46060 64034 46116 64036
rect 46060 63982 46062 64034
rect 46062 63982 46114 64034
rect 46114 63982 46116 64034
rect 46060 63980 46116 63982
rect 45948 63922 46004 63924
rect 45948 63870 45950 63922
rect 45950 63870 46002 63922
rect 46002 63870 46004 63922
rect 45948 63868 46004 63870
rect 46508 65324 46564 65380
rect 46508 64204 46564 64260
rect 46060 63138 46116 63140
rect 46060 63086 46062 63138
rect 46062 63086 46114 63138
rect 46114 63086 46116 63138
rect 46060 63084 46116 63086
rect 46060 62412 46116 62468
rect 44156 61404 44212 61460
rect 45724 62354 45780 62356
rect 45724 62302 45726 62354
rect 45726 62302 45778 62354
rect 45778 62302 45780 62354
rect 45724 62300 45780 62302
rect 46956 64204 47012 64260
rect 46508 62412 46564 62468
rect 47292 63084 47348 63140
rect 47180 62914 47236 62916
rect 47180 62862 47182 62914
rect 47182 62862 47234 62914
rect 47234 62862 47236 62914
rect 47180 62860 47236 62862
rect 48412 66498 48468 66500
rect 48412 66446 48414 66498
rect 48414 66446 48466 66498
rect 48466 66446 48468 66498
rect 48412 66444 48468 66446
rect 49084 66444 49140 66500
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 52220 66498 52276 66500
rect 52220 66446 52222 66498
rect 52222 66446 52274 66498
rect 52274 66446 52276 66498
rect 52220 66444 52276 66446
rect 53116 66444 53172 66500
rect 51100 65548 51156 65604
rect 47740 65378 47796 65380
rect 47740 65326 47742 65378
rect 47742 65326 47794 65378
rect 47794 65326 47796 65378
rect 47740 65324 47796 65326
rect 47516 64316 47572 64372
rect 44268 60226 44324 60228
rect 44268 60174 44270 60226
rect 44270 60174 44322 60226
rect 44322 60174 44324 60226
rect 44268 60172 44324 60174
rect 44940 59948 44996 60004
rect 44156 59388 44212 59444
rect 43820 59164 43876 59220
rect 45276 59218 45332 59220
rect 45276 59166 45278 59218
rect 45278 59166 45330 59218
rect 45330 59166 45332 59218
rect 45276 59164 45332 59166
rect 45724 59218 45780 59220
rect 45724 59166 45726 59218
rect 45726 59166 45778 59218
rect 45778 59166 45780 59218
rect 45724 59164 45780 59166
rect 43260 58716 43316 58772
rect 41132 58268 41188 58324
rect 40236 53676 40292 53732
rect 40908 53618 40964 53620
rect 40908 53566 40910 53618
rect 40910 53566 40962 53618
rect 40962 53566 40964 53618
rect 40908 53564 40964 53566
rect 41020 53506 41076 53508
rect 41020 53454 41022 53506
rect 41022 53454 41074 53506
rect 41074 53454 41076 53506
rect 41020 53452 41076 53454
rect 40124 51996 40180 52052
rect 41020 50764 41076 50820
rect 39228 49868 39284 49924
rect 39340 49980 39396 50036
rect 38444 47458 38500 47460
rect 38444 47406 38446 47458
rect 38446 47406 38498 47458
rect 38498 47406 38500 47458
rect 38444 47404 38500 47406
rect 38556 47234 38612 47236
rect 38556 47182 38558 47234
rect 38558 47182 38610 47234
rect 38610 47182 38612 47234
rect 38556 47180 38612 47182
rect 39004 47068 39060 47124
rect 38892 46674 38948 46676
rect 38892 46622 38894 46674
rect 38894 46622 38946 46674
rect 38946 46622 38948 46674
rect 38892 46620 38948 46622
rect 38220 46284 38276 46340
rect 37996 45612 38052 45668
rect 38444 45612 38500 45668
rect 38892 45276 38948 45332
rect 38892 44268 38948 44324
rect 36876 41692 36932 41748
rect 36764 38892 36820 38948
rect 37100 39676 37156 39732
rect 35532 37548 35588 37604
rect 35756 37378 35812 37380
rect 35756 37326 35758 37378
rect 35758 37326 35810 37378
rect 35810 37326 35812 37378
rect 35756 37324 35812 37326
rect 35644 37212 35700 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35980 36988 36036 37044
rect 35420 36482 35476 36484
rect 35420 36430 35422 36482
rect 35422 36430 35474 36482
rect 35474 36430 35476 36482
rect 35420 36428 35476 36430
rect 35084 36092 35140 36148
rect 34748 34972 34804 35028
rect 34188 33516 34244 33572
rect 33180 30156 33236 30212
rect 33628 32396 33684 32452
rect 33516 28588 33572 28644
rect 34300 33346 34356 33348
rect 34300 33294 34302 33346
rect 34302 33294 34354 33346
rect 34354 33294 34356 33346
rect 34300 33292 34356 33294
rect 34076 32060 34132 32116
rect 34300 31948 34356 32004
rect 34300 31778 34356 31780
rect 34300 31726 34302 31778
rect 34302 31726 34354 31778
rect 34354 31726 34356 31778
rect 34300 31724 34356 31726
rect 36092 36316 36148 36372
rect 35980 36092 36036 36148
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35868 35308 35924 35364
rect 35404 35252 35460 35254
rect 35756 35026 35812 35028
rect 35756 34974 35758 35026
rect 35758 34974 35810 35026
rect 35810 34974 35812 35026
rect 35756 34972 35812 34974
rect 34972 34076 35028 34132
rect 34972 33516 35028 33572
rect 35084 34748 35140 34804
rect 37100 38780 37156 38836
rect 41020 50034 41076 50036
rect 41020 49982 41022 50034
rect 41022 49982 41074 50034
rect 41074 49982 41076 50034
rect 41020 49980 41076 49982
rect 43148 58380 43204 58436
rect 42588 57538 42644 57540
rect 42588 57486 42590 57538
rect 42590 57486 42642 57538
rect 42642 57486 42644 57538
rect 42588 57484 42644 57486
rect 44828 58380 44884 58436
rect 45276 58492 45332 58548
rect 43148 57538 43204 57540
rect 43148 57486 43150 57538
rect 43150 57486 43202 57538
rect 43202 57486 43204 57538
rect 43148 57484 43204 57486
rect 43596 57596 43652 57652
rect 42252 56866 42308 56868
rect 42252 56814 42254 56866
rect 42254 56814 42306 56866
rect 42306 56814 42308 56866
rect 42252 56812 42308 56814
rect 42924 56700 42980 56756
rect 41692 55916 41748 55972
rect 41580 55410 41636 55412
rect 41580 55358 41582 55410
rect 41582 55358 41634 55410
rect 41634 55358 41636 55410
rect 41580 55356 41636 55358
rect 41468 55020 41524 55076
rect 42924 55916 42980 55972
rect 43260 56754 43316 56756
rect 43260 56702 43262 56754
rect 43262 56702 43314 56754
rect 43314 56702 43316 56754
rect 43260 56700 43316 56702
rect 44492 57650 44548 57652
rect 44492 57598 44494 57650
rect 44494 57598 44546 57650
rect 44546 57598 44548 57650
rect 44492 57596 44548 57598
rect 45500 55970 45556 55972
rect 45500 55918 45502 55970
rect 45502 55918 45554 55970
rect 45554 55918 45556 55970
rect 45500 55916 45556 55918
rect 42140 55410 42196 55412
rect 42140 55358 42142 55410
rect 42142 55358 42194 55410
rect 42194 55358 42196 55410
rect 42140 55356 42196 55358
rect 41804 54738 41860 54740
rect 41804 54686 41806 54738
rect 41806 54686 41858 54738
rect 41858 54686 41860 54738
rect 41804 54684 41860 54686
rect 44268 55244 44324 55300
rect 42364 55020 42420 55076
rect 44940 55298 44996 55300
rect 44940 55246 44942 55298
rect 44942 55246 44994 55298
rect 44994 55246 44996 55298
rect 44940 55244 44996 55246
rect 42476 54738 42532 54740
rect 42476 54686 42478 54738
rect 42478 54686 42530 54738
rect 42530 54686 42532 54738
rect 42476 54684 42532 54686
rect 42028 53788 42084 53844
rect 42476 54012 42532 54068
rect 41356 53340 41412 53396
rect 47068 59388 47124 59444
rect 46956 58546 47012 58548
rect 46956 58494 46958 58546
rect 46958 58494 47010 58546
rect 47010 58494 47012 58546
rect 46956 58492 47012 58494
rect 47068 57372 47124 57428
rect 47740 63420 47796 63476
rect 47740 63084 47796 63140
rect 48860 62524 48916 62580
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 52332 65436 52388 65492
rect 49532 63922 49588 63924
rect 49532 63870 49534 63922
rect 49534 63870 49586 63922
rect 49586 63870 49588 63922
rect 49532 63868 49588 63870
rect 49980 63196 50036 63252
rect 49644 63084 49700 63140
rect 48860 61852 48916 61908
rect 48860 60172 48916 60228
rect 50092 62188 50148 62244
rect 49084 61010 49140 61012
rect 49084 60958 49086 61010
rect 49086 60958 49138 61010
rect 49138 60958 49140 61010
rect 49084 60956 49140 60958
rect 48300 59388 48356 59444
rect 48188 59330 48244 59332
rect 48188 59278 48190 59330
rect 48190 59278 48242 59330
rect 48242 59278 48244 59330
rect 48188 59276 48244 59278
rect 48636 59164 48692 59220
rect 48188 57372 48244 57428
rect 47628 56252 47684 56308
rect 46396 55916 46452 55972
rect 44268 54012 44324 54068
rect 44268 53676 44324 53732
rect 47964 56252 48020 56308
rect 46732 55356 46788 55412
rect 46060 54572 46116 54628
rect 46844 54572 46900 54628
rect 46956 55132 47012 55188
rect 45500 53564 45556 53620
rect 45836 53676 45892 53732
rect 43820 52780 43876 52836
rect 45500 52220 45556 52276
rect 43148 52050 43204 52052
rect 43148 51998 43150 52050
rect 43150 51998 43202 52050
rect 43202 51998 43204 52050
rect 43148 51996 43204 51998
rect 44156 52050 44212 52052
rect 44156 51998 44158 52050
rect 44158 51998 44210 52050
rect 44210 51998 44212 52050
rect 44156 51996 44212 51998
rect 42476 51548 42532 51604
rect 43260 51602 43316 51604
rect 43260 51550 43262 51602
rect 43262 51550 43314 51602
rect 43314 51550 43316 51602
rect 43260 51548 43316 51550
rect 41244 51154 41300 51156
rect 41244 51102 41246 51154
rect 41246 51102 41298 51154
rect 41298 51102 41300 51154
rect 41244 51100 41300 51102
rect 41468 50594 41524 50596
rect 41468 50542 41470 50594
rect 41470 50542 41522 50594
rect 41522 50542 41524 50594
rect 41468 50540 41524 50542
rect 43260 51324 43316 51380
rect 41804 51212 41860 51268
rect 42252 51266 42308 51268
rect 42252 51214 42254 51266
rect 42254 51214 42306 51266
rect 42306 51214 42308 51266
rect 42252 51212 42308 51214
rect 41692 51154 41748 51156
rect 41692 51102 41694 51154
rect 41694 51102 41746 51154
rect 41746 51102 41748 51154
rect 41692 51100 41748 51102
rect 41804 50818 41860 50820
rect 41804 50766 41806 50818
rect 41806 50766 41858 50818
rect 41858 50766 41860 50818
rect 41804 50764 41860 50766
rect 41468 49810 41524 49812
rect 41468 49758 41470 49810
rect 41470 49758 41522 49810
rect 41522 49758 41524 49810
rect 41468 49756 41524 49758
rect 42140 49980 42196 50036
rect 39900 46786 39956 46788
rect 39900 46734 39902 46786
rect 39902 46734 39954 46786
rect 39954 46734 39956 46786
rect 39900 46732 39956 46734
rect 41020 46508 41076 46564
rect 39564 46396 39620 46452
rect 40908 46450 40964 46452
rect 40908 46398 40910 46450
rect 40910 46398 40962 46450
rect 40962 46398 40964 46450
rect 40908 46396 40964 46398
rect 40796 44322 40852 44324
rect 40796 44270 40798 44322
rect 40798 44270 40850 44322
rect 40850 44270 40852 44322
rect 40796 44268 40852 44270
rect 37772 42700 37828 42756
rect 38108 42140 38164 42196
rect 39452 42754 39508 42756
rect 39452 42702 39454 42754
rect 39454 42702 39506 42754
rect 39506 42702 39508 42754
rect 39452 42700 39508 42702
rect 39228 42028 39284 42084
rect 38220 41916 38276 41972
rect 38108 41858 38164 41860
rect 38108 41806 38110 41858
rect 38110 41806 38162 41858
rect 38162 41806 38164 41858
rect 38108 41804 38164 41806
rect 37660 41186 37716 41188
rect 37660 41134 37662 41186
rect 37662 41134 37714 41186
rect 37714 41134 37716 41186
rect 37660 41132 37716 41134
rect 38108 40460 38164 40516
rect 38892 41916 38948 41972
rect 36876 37772 36932 37828
rect 37548 38668 37604 38724
rect 39004 38946 39060 38948
rect 39004 38894 39006 38946
rect 39006 38894 39058 38946
rect 39058 38894 39060 38946
rect 39004 38892 39060 38894
rect 37884 38108 37940 38164
rect 37212 37938 37268 37940
rect 37212 37886 37214 37938
rect 37214 37886 37266 37938
rect 37266 37886 37268 37938
rect 37212 37884 37268 37886
rect 37100 37490 37156 37492
rect 37100 37438 37102 37490
rect 37102 37438 37154 37490
rect 37154 37438 37156 37490
rect 37100 37436 37156 37438
rect 37436 37826 37492 37828
rect 37436 37774 37438 37826
rect 37438 37774 37490 37826
rect 37490 37774 37492 37826
rect 37436 37772 37492 37774
rect 37772 37378 37828 37380
rect 37772 37326 37774 37378
rect 37774 37326 37826 37378
rect 37826 37326 37828 37378
rect 37772 37324 37828 37326
rect 37324 36876 37380 36932
rect 37212 36428 37268 36484
rect 36204 34972 36260 35028
rect 36540 36092 36596 36148
rect 36540 35532 36596 35588
rect 36988 35308 37044 35364
rect 36764 34130 36820 34132
rect 36764 34078 36766 34130
rect 36766 34078 36818 34130
rect 36818 34078 36820 34130
rect 36764 34076 36820 34078
rect 36876 33964 36932 34020
rect 37772 36988 37828 37044
rect 37660 36876 37716 36932
rect 37548 35084 37604 35140
rect 37100 34748 37156 34804
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34972 33068 35028 33124
rect 34748 32396 34804 32452
rect 34860 32620 34916 32676
rect 36204 32396 36260 32452
rect 37100 33122 37156 33124
rect 37100 33070 37102 33122
rect 37102 33070 37154 33122
rect 37154 33070 37156 33122
rect 37100 33068 37156 33070
rect 36988 32620 37044 32676
rect 37212 32732 37268 32788
rect 34860 32060 34916 32116
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 36204 32172 36260 32228
rect 35404 32116 35460 32118
rect 34748 31890 34804 31892
rect 34748 31838 34750 31890
rect 34750 31838 34802 31890
rect 34802 31838 34804 31890
rect 34748 31836 34804 31838
rect 35308 31948 35364 32004
rect 35196 31666 35252 31668
rect 35196 31614 35198 31666
rect 35198 31614 35250 31666
rect 35250 31614 35252 31666
rect 35196 31612 35252 31614
rect 35756 32002 35812 32004
rect 35756 31950 35758 32002
rect 35758 31950 35810 32002
rect 35810 31950 35812 32002
rect 35756 31948 35812 31950
rect 37436 33964 37492 34020
rect 38780 38162 38836 38164
rect 38780 38110 38782 38162
rect 38782 38110 38834 38162
rect 38834 38110 38836 38162
rect 38780 38108 38836 38110
rect 37996 37436 38052 37492
rect 37996 36316 38052 36372
rect 38668 37884 38724 37940
rect 38780 37324 38836 37380
rect 39676 38556 39732 38612
rect 39564 37378 39620 37380
rect 39564 37326 39566 37378
rect 39566 37326 39618 37378
rect 39618 37326 39620 37378
rect 39564 37324 39620 37326
rect 39228 37100 39284 37156
rect 39676 37100 39732 37156
rect 38556 36482 38612 36484
rect 38556 36430 38558 36482
rect 38558 36430 38610 36482
rect 38610 36430 38612 36482
rect 38556 36428 38612 36430
rect 38220 36092 38276 36148
rect 39228 36428 39284 36484
rect 37436 32508 37492 32564
rect 38332 35308 38388 35364
rect 38332 35084 38388 35140
rect 38220 35026 38276 35028
rect 38220 34974 38222 35026
rect 38222 34974 38274 35026
rect 38274 34974 38276 35026
rect 38220 34972 38276 34974
rect 37996 34076 38052 34132
rect 38332 34076 38388 34132
rect 38108 33234 38164 33236
rect 38108 33182 38110 33234
rect 38110 33182 38162 33234
rect 38162 33182 38164 33234
rect 38108 33180 38164 33182
rect 38108 32786 38164 32788
rect 38108 32734 38110 32786
rect 38110 32734 38162 32786
rect 38162 32734 38164 32786
rect 38108 32732 38164 32734
rect 37660 32508 37716 32564
rect 37212 31948 37268 32004
rect 37884 31890 37940 31892
rect 37884 31838 37886 31890
rect 37886 31838 37938 31890
rect 37938 31838 37940 31890
rect 37884 31836 37940 31838
rect 35420 31778 35476 31780
rect 35420 31726 35422 31778
rect 35422 31726 35474 31778
rect 35474 31726 35476 31778
rect 35420 31724 35476 31726
rect 35868 31724 35924 31780
rect 37996 31778 38052 31780
rect 37996 31726 37998 31778
rect 37998 31726 38050 31778
rect 38050 31726 38052 31778
rect 37996 31724 38052 31726
rect 34860 30716 34916 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35420 30098 35476 30100
rect 35420 30046 35422 30098
rect 35422 30046 35474 30098
rect 35474 30046 35476 30098
rect 35420 30044 35476 30046
rect 34524 29932 34580 29988
rect 35084 29708 35140 29764
rect 35196 29034 35252 29036
rect 34524 28924 34580 28980
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 33852 28028 33908 28084
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 34860 28588 34916 28644
rect 34524 28140 34580 28196
rect 34972 27804 35028 27860
rect 35308 27580 35364 27636
rect 36428 29596 36484 29652
rect 35868 29148 35924 29204
rect 35868 28700 35924 28756
rect 36988 29596 37044 29652
rect 36876 29426 36932 29428
rect 36876 29374 36878 29426
rect 36878 29374 36930 29426
rect 36930 29374 36932 29426
rect 36876 29372 36932 29374
rect 36092 28140 36148 28196
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34412 26796 34468 26852
rect 33292 26348 33348 26404
rect 32396 25900 32452 25956
rect 32620 25452 32676 25508
rect 33852 25676 33908 25732
rect 32956 25394 33012 25396
rect 32956 25342 32958 25394
rect 32958 25342 33010 25394
rect 33010 25342 33012 25394
rect 32956 25340 33012 25342
rect 33180 25282 33236 25284
rect 33180 25230 33182 25282
rect 33182 25230 33234 25282
rect 33234 25230 33236 25282
rect 33180 25228 33236 25230
rect 32284 25116 32340 25172
rect 29708 24556 29764 24612
rect 31724 24444 31780 24500
rect 31612 23826 31668 23828
rect 31612 23774 31614 23826
rect 31614 23774 31666 23826
rect 31666 23774 31668 23826
rect 31612 23772 31668 23774
rect 29932 23660 29988 23716
rect 30716 23324 30772 23380
rect 30716 22988 30772 23044
rect 30156 20914 30212 20916
rect 30156 20862 30158 20914
rect 30158 20862 30210 20914
rect 30210 20862 30212 20914
rect 30156 20860 30212 20862
rect 30940 20748 30996 20804
rect 29036 20132 29092 20188
rect 28252 19964 28308 20020
rect 28476 18674 28532 18676
rect 28476 18622 28478 18674
rect 28478 18622 28530 18674
rect 28530 18622 28532 18674
rect 28476 18620 28532 18622
rect 29372 18620 29428 18676
rect 28588 18450 28644 18452
rect 28588 18398 28590 18450
rect 28590 18398 28642 18450
rect 28642 18398 28644 18450
rect 28588 18396 28644 18398
rect 28924 18284 28980 18340
rect 27916 17388 27972 17444
rect 28364 17442 28420 17444
rect 28364 17390 28366 17442
rect 28366 17390 28418 17442
rect 28418 17390 28420 17442
rect 28364 17388 28420 17390
rect 28700 17164 28756 17220
rect 28812 17612 28868 17668
rect 27468 15986 27524 15988
rect 27468 15934 27470 15986
rect 27470 15934 27522 15986
rect 27522 15934 27524 15986
rect 27468 15932 27524 15934
rect 25228 15708 25284 15764
rect 26796 14812 26852 14868
rect 26460 14642 26516 14644
rect 26460 14590 26462 14642
rect 26462 14590 26514 14642
rect 26514 14590 26516 14642
rect 26460 14588 26516 14590
rect 25228 12962 25284 12964
rect 25228 12910 25230 12962
rect 25230 12910 25282 12962
rect 25282 12910 25284 12962
rect 25228 12908 25284 12910
rect 25228 12684 25284 12740
rect 25340 10610 25396 10612
rect 25340 10558 25342 10610
rect 25342 10558 25394 10610
rect 25394 10558 25396 10610
rect 25340 10556 25396 10558
rect 25004 9884 25060 9940
rect 25340 10332 25396 10388
rect 27580 14642 27636 14644
rect 27580 14590 27582 14642
rect 27582 14590 27634 14642
rect 27634 14590 27636 14642
rect 27580 14588 27636 14590
rect 27132 14306 27188 14308
rect 27132 14254 27134 14306
rect 27134 14254 27186 14306
rect 27186 14254 27188 14306
rect 27132 14252 27188 14254
rect 28140 17052 28196 17108
rect 28252 16716 28308 16772
rect 28812 16770 28868 16772
rect 28812 16718 28814 16770
rect 28814 16718 28866 16770
rect 28866 16718 28868 16770
rect 28812 16716 28868 16718
rect 28140 15986 28196 15988
rect 28140 15934 28142 15986
rect 28142 15934 28194 15986
rect 28194 15934 28196 15986
rect 28140 15932 28196 15934
rect 28364 15986 28420 15988
rect 28364 15934 28366 15986
rect 28366 15934 28418 15986
rect 28418 15934 28420 15986
rect 28364 15932 28420 15934
rect 28476 14700 28532 14756
rect 28140 14252 28196 14308
rect 26684 12684 26740 12740
rect 27020 12012 27076 12068
rect 27468 12738 27524 12740
rect 27468 12686 27470 12738
rect 27470 12686 27522 12738
rect 27522 12686 27524 12738
rect 27468 12684 27524 12686
rect 27132 11452 27188 11508
rect 26684 9772 26740 9828
rect 25452 8428 25508 8484
rect 24108 7250 24164 7252
rect 24108 7198 24110 7250
rect 24110 7198 24162 7250
rect 24162 7198 24164 7250
rect 24108 7196 24164 7198
rect 24444 6972 24500 7028
rect 24332 6802 24388 6804
rect 24332 6750 24334 6802
rect 24334 6750 24386 6802
rect 24386 6750 24388 6802
rect 24332 6748 24388 6750
rect 23996 6300 24052 6356
rect 24108 6578 24164 6580
rect 24108 6526 24110 6578
rect 24110 6526 24162 6578
rect 24162 6526 24164 6578
rect 24108 6524 24164 6526
rect 24108 6188 24164 6244
rect 25116 6636 25172 6692
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 25004 6578 25060 6580
rect 25004 6526 25006 6578
rect 25006 6526 25058 6578
rect 25058 6526 25060 6578
rect 25004 6524 25060 6526
rect 26572 8428 26628 8484
rect 26348 7474 26404 7476
rect 26348 7422 26350 7474
rect 26350 7422 26402 7474
rect 26402 7422 26404 7474
rect 26348 7420 26404 7422
rect 27468 12012 27524 12068
rect 27468 11452 27524 11508
rect 27132 10556 27188 10612
rect 27020 10220 27076 10276
rect 27468 9884 27524 9940
rect 27804 12012 27860 12068
rect 29708 17388 29764 17444
rect 30492 19964 30548 20020
rect 30268 18956 30324 19012
rect 29932 18732 29988 18788
rect 29372 15986 29428 15988
rect 29372 15934 29374 15986
rect 29374 15934 29426 15986
rect 29426 15934 29428 15986
rect 29372 15932 29428 15934
rect 28924 13804 28980 13860
rect 28476 13020 28532 13076
rect 29484 12962 29540 12964
rect 29484 12910 29486 12962
rect 29486 12910 29538 12962
rect 29538 12910 29540 12962
rect 29484 12908 29540 12910
rect 28252 12066 28308 12068
rect 28252 12014 28254 12066
rect 28254 12014 28306 12066
rect 28306 12014 28308 12066
rect 28252 12012 28308 12014
rect 28252 11564 28308 11620
rect 29260 11506 29316 11508
rect 29260 11454 29262 11506
rect 29262 11454 29314 11506
rect 29314 11454 29316 11506
rect 29260 11452 29316 11454
rect 29932 13580 29988 13636
rect 30044 13804 30100 13860
rect 29932 12908 29988 12964
rect 30380 18620 30436 18676
rect 31052 20018 31108 20020
rect 31052 19966 31054 20018
rect 31054 19966 31106 20018
rect 31106 19966 31108 20018
rect 31052 19964 31108 19966
rect 30716 18956 30772 19012
rect 30492 17666 30548 17668
rect 30492 17614 30494 17666
rect 30494 17614 30546 17666
rect 30546 17614 30548 17666
rect 30492 17612 30548 17614
rect 31612 20130 31668 20132
rect 31612 20078 31614 20130
rect 31614 20078 31666 20130
rect 31666 20078 31668 20130
rect 31612 20076 31668 20078
rect 31388 20018 31444 20020
rect 31388 19966 31390 20018
rect 31390 19966 31442 20018
rect 31442 19966 31444 20018
rect 31388 19964 31444 19966
rect 32060 23826 32116 23828
rect 32060 23774 32062 23826
rect 32062 23774 32114 23826
rect 32114 23774 32116 23826
rect 32060 23772 32116 23774
rect 31948 23436 32004 23492
rect 31948 21644 32004 21700
rect 33516 25452 33572 25508
rect 33628 25228 33684 25284
rect 33404 23436 33460 23492
rect 34188 25676 34244 25732
rect 34972 25676 35028 25732
rect 34636 25452 34692 25508
rect 34076 25282 34132 25284
rect 34076 25230 34078 25282
rect 34078 25230 34130 25282
rect 34130 25230 34132 25282
rect 34076 25228 34132 25230
rect 34188 24780 34244 24836
rect 32060 20130 32116 20132
rect 32060 20078 32062 20130
rect 32062 20078 32114 20130
rect 32114 20078 32116 20130
rect 32060 20076 32116 20078
rect 31836 19964 31892 20020
rect 31500 19068 31556 19124
rect 31388 18338 31444 18340
rect 31388 18286 31390 18338
rect 31390 18286 31442 18338
rect 31442 18286 31444 18338
rect 31388 18284 31444 18286
rect 30940 17724 30996 17780
rect 30828 17388 30884 17444
rect 31388 17724 31444 17780
rect 31164 17666 31220 17668
rect 31164 17614 31166 17666
rect 31166 17614 31218 17666
rect 31218 17614 31220 17666
rect 31164 17612 31220 17614
rect 31612 17666 31668 17668
rect 31612 17614 31614 17666
rect 31614 17614 31666 17666
rect 31666 17614 31668 17666
rect 31612 17612 31668 17614
rect 31500 17164 31556 17220
rect 30492 13634 30548 13636
rect 30492 13582 30494 13634
rect 30494 13582 30546 13634
rect 30546 13582 30548 13634
rect 30492 13580 30548 13582
rect 30156 12178 30212 12180
rect 30156 12126 30158 12178
rect 30158 12126 30210 12178
rect 30210 12126 30212 12178
rect 30156 12124 30212 12126
rect 30604 11788 30660 11844
rect 29708 11564 29764 11620
rect 30156 11452 30212 11508
rect 27580 10108 27636 10164
rect 27356 8258 27412 8260
rect 27356 8206 27358 8258
rect 27358 8206 27410 8258
rect 27410 8206 27412 8258
rect 27356 8204 27412 8206
rect 29596 9884 29652 9940
rect 28028 9826 28084 9828
rect 28028 9774 28030 9826
rect 28030 9774 28082 9826
rect 28082 9774 28084 9826
rect 28028 9772 28084 9774
rect 28588 9714 28644 9716
rect 28588 9662 28590 9714
rect 28590 9662 28642 9714
rect 28642 9662 28644 9714
rect 28588 9660 28644 9662
rect 29932 9714 29988 9716
rect 29932 9662 29934 9714
rect 29934 9662 29986 9714
rect 29986 9662 29988 9714
rect 29932 9660 29988 9662
rect 30044 9602 30100 9604
rect 30044 9550 30046 9602
rect 30046 9550 30098 9602
rect 30098 9550 30100 9602
rect 30044 9548 30100 9550
rect 29708 9436 29764 9492
rect 28028 8092 28084 8148
rect 26908 7980 26964 8036
rect 25788 7362 25844 7364
rect 25788 7310 25790 7362
rect 25790 7310 25842 7362
rect 25842 7310 25844 7362
rect 25788 7308 25844 7310
rect 25900 7196 25956 7252
rect 26796 7308 26852 7364
rect 25900 6860 25956 6916
rect 27020 7308 27076 7364
rect 27244 7474 27300 7476
rect 27244 7422 27246 7474
rect 27246 7422 27298 7474
rect 27298 7422 27300 7474
rect 27244 7420 27300 7422
rect 27692 7362 27748 7364
rect 27692 7310 27694 7362
rect 27694 7310 27746 7362
rect 27746 7310 27748 7362
rect 27692 7308 27748 7310
rect 27244 6860 27300 6916
rect 26236 6636 26292 6692
rect 27244 6636 27300 6692
rect 29820 7980 29876 8036
rect 30492 9938 30548 9940
rect 30492 9886 30494 9938
rect 30494 9886 30546 9938
rect 30546 9886 30548 9938
rect 30492 9884 30548 9886
rect 31724 16268 31780 16324
rect 31948 19068 32004 19124
rect 31724 15820 31780 15876
rect 31948 18732 32004 18788
rect 31724 15202 31780 15204
rect 31724 15150 31726 15202
rect 31726 15150 31778 15202
rect 31778 15150 31780 15202
rect 31724 15148 31780 15150
rect 32172 18396 32228 18452
rect 32284 18172 32340 18228
rect 32508 16770 32564 16772
rect 32508 16718 32510 16770
rect 32510 16718 32562 16770
rect 32562 16718 32564 16770
rect 32508 16716 32564 16718
rect 32172 16210 32228 16212
rect 32172 16158 32174 16210
rect 32174 16158 32226 16210
rect 32226 16158 32228 16210
rect 32172 16156 32228 16158
rect 32508 15148 32564 15204
rect 32060 15090 32116 15092
rect 32060 15038 32062 15090
rect 32062 15038 32114 15090
rect 32114 15038 32116 15090
rect 32060 15036 32116 15038
rect 31612 12572 31668 12628
rect 31500 11788 31556 11844
rect 32172 13692 32228 13748
rect 31836 13580 31892 13636
rect 32060 12908 32116 12964
rect 32172 12796 32228 12852
rect 32396 12796 32452 12852
rect 33180 22988 33236 23044
rect 33628 22652 33684 22708
rect 33852 22876 33908 22932
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35420 25564 35476 25620
rect 35420 25394 35476 25396
rect 35420 25342 35422 25394
rect 35422 25342 35474 25394
rect 35474 25342 35476 25394
rect 35420 25340 35476 25342
rect 36204 25676 36260 25732
rect 36988 28700 37044 28756
rect 37772 29820 37828 29876
rect 37100 28588 37156 28644
rect 37100 28140 37156 28196
rect 37884 29372 37940 29428
rect 37436 28140 37492 28196
rect 37772 27580 37828 27636
rect 35420 24722 35476 24724
rect 35420 24670 35422 24722
rect 35422 24670 35474 24722
rect 35474 24670 35476 24722
rect 35420 24668 35476 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36092 25228 36148 25284
rect 35980 24556 36036 24612
rect 35084 22876 35140 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35532 22428 35588 22484
rect 33068 18732 33124 18788
rect 33180 17388 33236 17444
rect 32732 15820 32788 15876
rect 33180 15874 33236 15876
rect 33180 15822 33182 15874
rect 33182 15822 33234 15874
rect 33234 15822 33236 15874
rect 33180 15820 33236 15822
rect 32732 14588 32788 14644
rect 33068 13746 33124 13748
rect 33068 13694 33070 13746
rect 33070 13694 33122 13746
rect 33122 13694 33124 13746
rect 33068 13692 33124 13694
rect 32620 12908 32676 12964
rect 32508 12572 32564 12628
rect 33628 21810 33684 21812
rect 33628 21758 33630 21810
rect 33630 21758 33682 21810
rect 33682 21758 33684 21810
rect 33628 21756 33684 21758
rect 34524 21644 34580 21700
rect 33964 20802 34020 20804
rect 33964 20750 33966 20802
rect 33966 20750 34018 20802
rect 34018 20750 34020 20802
rect 33964 20748 34020 20750
rect 33740 19404 33796 19460
rect 34860 21586 34916 21588
rect 34860 21534 34862 21586
rect 34862 21534 34914 21586
rect 34914 21534 34916 21586
rect 34860 21532 34916 21534
rect 34188 19404 34244 19460
rect 34524 19292 34580 19348
rect 34188 19068 34244 19124
rect 33516 18396 33572 18452
rect 33628 18956 33684 19012
rect 33852 18674 33908 18676
rect 33852 18622 33854 18674
rect 33854 18622 33906 18674
rect 33906 18622 33908 18674
rect 33852 18620 33908 18622
rect 33628 18508 33684 18564
rect 33628 16156 33684 16212
rect 34188 16716 34244 16772
rect 33852 15148 33908 15204
rect 33404 15036 33460 15092
rect 33404 13356 33460 13412
rect 31836 11676 31892 11732
rect 32060 11228 32116 11284
rect 31164 10892 31220 10948
rect 31164 9884 31220 9940
rect 31388 9772 31444 9828
rect 31052 9660 31108 9716
rect 30604 9602 30660 9604
rect 30604 9550 30606 9602
rect 30606 9550 30658 9602
rect 30658 9550 30660 9602
rect 30604 9548 30660 9550
rect 28140 7420 28196 7476
rect 26460 6466 26516 6468
rect 26460 6414 26462 6466
rect 26462 6414 26514 6466
rect 26514 6414 26516 6466
rect 26460 6412 26516 6414
rect 27692 6412 27748 6468
rect 26236 6188 26292 6244
rect 25340 4338 25396 4340
rect 25340 4286 25342 4338
rect 25342 4286 25394 4338
rect 25394 4286 25396 4338
rect 25340 4284 25396 4286
rect 30492 6636 30548 6692
rect 29372 6524 29428 6580
rect 30156 6188 30212 6244
rect 29372 5852 29428 5908
rect 28588 4562 28644 4564
rect 28588 4510 28590 4562
rect 28590 4510 28642 4562
rect 28642 4510 28644 4562
rect 28588 4508 28644 4510
rect 30492 6188 30548 6244
rect 29708 5292 29764 5348
rect 30940 8316 30996 8372
rect 30716 8034 30772 8036
rect 30716 7982 30718 8034
rect 30718 7982 30770 8034
rect 30770 7982 30772 8034
rect 30716 7980 30772 7982
rect 31164 7980 31220 8036
rect 31724 10892 31780 10948
rect 31836 9826 31892 9828
rect 31836 9774 31838 9826
rect 31838 9774 31890 9826
rect 31890 9774 31892 9826
rect 31836 9772 31892 9774
rect 33740 14306 33796 14308
rect 33740 14254 33742 14306
rect 33742 14254 33794 14306
rect 33794 14254 33796 14306
rect 33740 14252 33796 14254
rect 33740 13692 33796 13748
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 32956 12908 33012 12964
rect 33292 12796 33348 12852
rect 32956 12124 33012 12180
rect 33516 11676 33572 11732
rect 33516 11340 33572 11396
rect 33292 11004 33348 11060
rect 32284 9938 32340 9940
rect 32284 9886 32286 9938
rect 32286 9886 32338 9938
rect 32338 9886 32340 9938
rect 32284 9884 32340 9886
rect 34188 13970 34244 13972
rect 34188 13918 34190 13970
rect 34190 13918 34242 13970
rect 34242 13918 34244 13970
rect 34188 13916 34244 13918
rect 34636 19010 34692 19012
rect 34636 18958 34638 19010
rect 34638 18958 34690 19010
rect 34690 18958 34692 19010
rect 34636 18956 34692 18958
rect 34972 19010 35028 19012
rect 34972 18958 34974 19010
rect 34974 18958 35026 19010
rect 35026 18958 35028 19010
rect 34972 18956 35028 18958
rect 35644 21586 35700 21588
rect 35644 21534 35646 21586
rect 35646 21534 35698 21586
rect 35698 21534 35700 21586
rect 35644 21532 35700 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35420 19122 35476 19124
rect 35420 19070 35422 19122
rect 35422 19070 35474 19122
rect 35474 19070 35476 19122
rect 35420 19068 35476 19070
rect 35084 18620 35140 18676
rect 34748 18450 34804 18452
rect 34748 18398 34750 18450
rect 34750 18398 34802 18450
rect 34802 18398 34804 18450
rect 34748 18396 34804 18398
rect 36092 18844 36148 18900
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35868 18396 35924 18452
rect 35980 18508 36036 18564
rect 35532 17836 35588 17892
rect 35084 17388 35140 17444
rect 38108 28140 38164 28196
rect 38108 27804 38164 27860
rect 38220 27244 38276 27300
rect 38444 31724 38500 31780
rect 38780 34412 38836 34468
rect 39116 33404 39172 33460
rect 38892 33346 38948 33348
rect 38892 33294 38894 33346
rect 38894 33294 38946 33346
rect 38946 33294 38948 33346
rect 38892 33292 38948 33294
rect 40124 43596 40180 43652
rect 41020 43538 41076 43540
rect 41020 43486 41022 43538
rect 41022 43486 41074 43538
rect 41074 43486 41076 43538
rect 41020 43484 41076 43486
rect 40348 43426 40404 43428
rect 40348 43374 40350 43426
rect 40350 43374 40402 43426
rect 40402 43374 40404 43426
rect 40348 43372 40404 43374
rect 42812 50594 42868 50596
rect 42812 50542 42814 50594
rect 42814 50542 42866 50594
rect 42866 50542 42868 50594
rect 42812 50540 42868 50542
rect 42252 49756 42308 49812
rect 42140 49698 42196 49700
rect 42140 49646 42142 49698
rect 42142 49646 42194 49698
rect 42194 49646 42196 49698
rect 42140 49644 42196 49646
rect 41580 48130 41636 48132
rect 41580 48078 41582 48130
rect 41582 48078 41634 48130
rect 41634 48078 41636 48130
rect 41580 48076 41636 48078
rect 41692 47516 41748 47572
rect 42364 48354 42420 48356
rect 42364 48302 42366 48354
rect 42366 48302 42418 48354
rect 42418 48302 42420 48354
rect 42364 48300 42420 48302
rect 42588 48076 42644 48132
rect 42140 47516 42196 47572
rect 41692 46562 41748 46564
rect 41692 46510 41694 46562
rect 41694 46510 41746 46562
rect 41746 46510 41748 46562
rect 41692 46508 41748 46510
rect 43708 51548 43764 51604
rect 43372 49644 43428 49700
rect 43596 51212 43652 51268
rect 43036 48188 43092 48244
rect 43372 48354 43428 48356
rect 43372 48302 43374 48354
rect 43374 48302 43426 48354
rect 43426 48302 43428 48354
rect 43372 48300 43428 48302
rect 42924 47516 42980 47572
rect 43484 48242 43540 48244
rect 43484 48190 43486 48242
rect 43486 48190 43538 48242
rect 43538 48190 43540 48242
rect 43484 48188 43540 48190
rect 44156 50540 44212 50596
rect 44828 50594 44884 50596
rect 44828 50542 44830 50594
rect 44830 50542 44882 50594
rect 44882 50542 44884 50594
rect 44828 50540 44884 50542
rect 45836 50594 45892 50596
rect 45836 50542 45838 50594
rect 45838 50542 45890 50594
rect 45890 50542 45892 50594
rect 45836 50540 45892 50542
rect 46396 54514 46452 54516
rect 46396 54462 46398 54514
rect 46398 54462 46450 54514
rect 46450 54462 46452 54514
rect 46396 54460 46452 54462
rect 46956 54460 47012 54516
rect 46844 54402 46900 54404
rect 46844 54350 46846 54402
rect 46846 54350 46898 54402
rect 46898 54350 46900 54402
rect 46844 54348 46900 54350
rect 47852 54348 47908 54404
rect 47852 53788 47908 53844
rect 47516 53228 47572 53284
rect 46844 53170 46900 53172
rect 46844 53118 46846 53170
rect 46846 53118 46898 53170
rect 46898 53118 46900 53170
rect 46844 53116 46900 53118
rect 46396 52946 46452 52948
rect 46396 52894 46398 52946
rect 46398 52894 46450 52946
rect 46450 52894 46452 52946
rect 46396 52892 46452 52894
rect 46732 52892 46788 52948
rect 46508 52834 46564 52836
rect 46508 52782 46510 52834
rect 46510 52782 46562 52834
rect 46562 52782 46564 52834
rect 46508 52780 46564 52782
rect 46732 52274 46788 52276
rect 46732 52222 46734 52274
rect 46734 52222 46786 52274
rect 46786 52222 46788 52274
rect 46732 52220 46788 52222
rect 47516 52892 47572 52948
rect 47180 52444 47236 52500
rect 47292 51378 47348 51380
rect 47292 51326 47294 51378
rect 47294 51326 47346 51378
rect 47346 51326 47348 51378
rect 47292 51324 47348 51326
rect 46060 50540 46116 50596
rect 46732 50594 46788 50596
rect 46732 50542 46734 50594
rect 46734 50542 46786 50594
rect 46786 50542 46788 50594
rect 46732 50540 46788 50542
rect 43596 47964 43652 48020
rect 43484 47180 43540 47236
rect 43596 47516 43652 47572
rect 43260 46732 43316 46788
rect 44268 47570 44324 47572
rect 44268 47518 44270 47570
rect 44270 47518 44322 47570
rect 44322 47518 44324 47570
rect 44268 47516 44324 47518
rect 44828 47516 44884 47572
rect 43932 46956 43988 47012
rect 44828 47180 44884 47236
rect 44492 46674 44548 46676
rect 44492 46622 44494 46674
rect 44494 46622 44546 46674
rect 44546 46622 44548 46674
rect 44492 46620 44548 46622
rect 48188 56140 48244 56196
rect 47964 53228 48020 53284
rect 48300 51602 48356 51604
rect 48300 51550 48302 51602
rect 48302 51550 48354 51602
rect 48354 51550 48356 51602
rect 48300 51548 48356 51550
rect 47628 50540 47684 50596
rect 45276 46956 45332 47012
rect 45052 46508 45108 46564
rect 42140 44268 42196 44324
rect 41468 43538 41524 43540
rect 41468 43486 41470 43538
rect 41470 43486 41522 43538
rect 41522 43486 41524 43538
rect 41468 43484 41524 43486
rect 42252 43372 42308 43428
rect 42476 43426 42532 43428
rect 42476 43374 42478 43426
rect 42478 43374 42530 43426
rect 42530 43374 42532 43426
rect 42476 43372 42532 43374
rect 43036 43372 43092 43428
rect 42252 42924 42308 42980
rect 40348 41970 40404 41972
rect 40348 41918 40350 41970
rect 40350 41918 40402 41970
rect 40402 41918 40404 41970
rect 40348 41916 40404 41918
rect 40236 40348 40292 40404
rect 40348 41132 40404 41188
rect 41132 41020 41188 41076
rect 41244 40402 41300 40404
rect 41244 40350 41246 40402
rect 41246 40350 41298 40402
rect 41298 40350 41300 40402
rect 41244 40348 41300 40350
rect 41468 40348 41524 40404
rect 41804 41970 41860 41972
rect 41804 41918 41806 41970
rect 41806 41918 41858 41970
rect 41858 41918 41860 41970
rect 41804 41916 41860 41918
rect 45388 46674 45444 46676
rect 45388 46622 45390 46674
rect 45390 46622 45442 46674
rect 45442 46622 45444 46674
rect 45388 46620 45444 46622
rect 45948 46956 46004 47012
rect 45724 46674 45780 46676
rect 45724 46622 45726 46674
rect 45726 46622 45778 46674
rect 45778 46622 45780 46674
rect 45724 46620 45780 46622
rect 45836 46562 45892 46564
rect 45836 46510 45838 46562
rect 45838 46510 45890 46562
rect 45890 46510 45892 46562
rect 45836 46508 45892 46510
rect 44156 43596 44212 43652
rect 44268 43932 44324 43988
rect 43596 42924 43652 42980
rect 44156 42924 44212 42980
rect 43708 42476 43764 42532
rect 42252 41074 42308 41076
rect 42252 41022 42254 41074
rect 42254 41022 42306 41074
rect 42306 41022 42308 41074
rect 42252 41020 42308 41022
rect 41804 40684 41860 40740
rect 40236 38556 40292 38612
rect 39676 34018 39732 34020
rect 39676 33966 39678 34018
rect 39678 33966 39730 34018
rect 39730 33966 39732 34018
rect 39676 33964 39732 33966
rect 40236 34412 40292 34468
rect 39452 32732 39508 32788
rect 38892 32172 38948 32228
rect 39564 32284 39620 32340
rect 38556 31612 38612 31668
rect 38892 29932 38948 29988
rect 39900 33292 39956 33348
rect 40348 34130 40404 34132
rect 40348 34078 40350 34130
rect 40350 34078 40402 34130
rect 40402 34078 40404 34130
rect 40348 34076 40404 34078
rect 39900 32396 39956 32452
rect 40348 29986 40404 29988
rect 40348 29934 40350 29986
rect 40350 29934 40402 29986
rect 40402 29934 40404 29986
rect 40348 29932 40404 29934
rect 39788 29820 39844 29876
rect 40236 29314 40292 29316
rect 40236 29262 40238 29314
rect 40238 29262 40290 29314
rect 40290 29262 40292 29314
rect 40236 29260 40292 29262
rect 38668 28642 38724 28644
rect 38668 28590 38670 28642
rect 38670 28590 38722 28642
rect 38722 28590 38724 28642
rect 38668 28588 38724 28590
rect 38444 27970 38500 27972
rect 38444 27918 38446 27970
rect 38446 27918 38498 27970
rect 38498 27918 38500 27970
rect 38444 27916 38500 27918
rect 39004 27970 39060 27972
rect 39004 27918 39006 27970
rect 39006 27918 39058 27970
rect 39058 27918 39060 27970
rect 39004 27916 39060 27918
rect 38668 27858 38724 27860
rect 38668 27806 38670 27858
rect 38670 27806 38722 27858
rect 38722 27806 38724 27858
rect 38668 27804 38724 27806
rect 40012 28028 40068 28084
rect 39116 27580 39172 27636
rect 40012 27074 40068 27076
rect 40012 27022 40014 27074
rect 40014 27022 40066 27074
rect 40066 27022 40068 27074
rect 40012 27020 40068 27022
rect 38668 26962 38724 26964
rect 38668 26910 38670 26962
rect 38670 26910 38722 26962
rect 38722 26910 38724 26962
rect 38668 26908 38724 26910
rect 39676 26908 39732 26964
rect 37996 26460 38052 26516
rect 38444 26460 38500 26516
rect 37212 25564 37268 25620
rect 37100 25282 37156 25284
rect 37100 25230 37102 25282
rect 37102 25230 37154 25282
rect 37154 25230 37156 25282
rect 37100 25228 37156 25230
rect 37436 25340 37492 25396
rect 37996 25282 38052 25284
rect 37996 25230 37998 25282
rect 37998 25230 38050 25282
rect 38050 25230 38052 25282
rect 37996 25228 38052 25230
rect 39228 26514 39284 26516
rect 39228 26462 39230 26514
rect 39230 26462 39282 26514
rect 39282 26462 39284 26514
rect 39228 26460 39284 26462
rect 39452 26290 39508 26292
rect 39452 26238 39454 26290
rect 39454 26238 39506 26290
rect 39506 26238 39508 26290
rect 39452 26236 39508 26238
rect 39340 26124 39396 26180
rect 39116 26066 39172 26068
rect 39116 26014 39118 26066
rect 39118 26014 39170 26066
rect 39170 26014 39172 26066
rect 39116 26012 39172 26014
rect 39788 26402 39844 26404
rect 39788 26350 39790 26402
rect 39790 26350 39842 26402
rect 39842 26350 39844 26402
rect 39788 26348 39844 26350
rect 39788 26012 39844 26068
rect 40124 26124 40180 26180
rect 40012 25564 40068 25620
rect 39228 25394 39284 25396
rect 39228 25342 39230 25394
rect 39230 25342 39282 25394
rect 39282 25342 39284 25394
rect 39228 25340 39284 25342
rect 36876 24444 36932 24500
rect 37884 24668 37940 24724
rect 38444 24668 38500 24724
rect 37884 23324 37940 23380
rect 36428 23100 36484 23156
rect 36428 22482 36484 22484
rect 36428 22430 36430 22482
rect 36430 22430 36482 22482
rect 36482 22430 36484 22482
rect 36428 22428 36484 22430
rect 37212 22316 37268 22372
rect 38108 23212 38164 23268
rect 36316 21756 36372 21812
rect 36764 21810 36820 21812
rect 36764 21758 36766 21810
rect 36766 21758 36818 21810
rect 36818 21758 36820 21810
rect 36764 21756 36820 21758
rect 36428 20188 36484 20244
rect 35420 17052 35476 17108
rect 35980 17442 36036 17444
rect 35980 17390 35982 17442
rect 35982 17390 36034 17442
rect 36034 17390 36036 17442
rect 35980 17388 36036 17390
rect 34636 15426 34692 15428
rect 34636 15374 34638 15426
rect 34638 15374 34690 15426
rect 34690 15374 34692 15426
rect 34636 15372 34692 15374
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35532 16156 35588 16212
rect 35532 15708 35588 15764
rect 35308 15372 35364 15428
rect 36092 16210 36148 16212
rect 36092 16158 36094 16210
rect 36094 16158 36146 16210
rect 36146 16158 36148 16210
rect 36092 16156 36148 16158
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34524 13916 34580 13972
rect 34076 13356 34132 13412
rect 33964 13132 34020 13188
rect 33964 11282 34020 11284
rect 33964 11230 33966 11282
rect 33966 11230 34018 11282
rect 34018 11230 34020 11282
rect 33964 11228 34020 11230
rect 32844 9996 32900 10052
rect 32172 9772 32228 9828
rect 33292 9826 33348 9828
rect 33292 9774 33294 9826
rect 33294 9774 33346 9826
rect 33346 9774 33348 9826
rect 33292 9772 33348 9774
rect 31612 8034 31668 8036
rect 31612 7982 31614 8034
rect 31614 7982 31666 8034
rect 31666 7982 31668 8034
rect 31612 7980 31668 7982
rect 30940 7644 30996 7700
rect 31500 7698 31556 7700
rect 31500 7646 31502 7698
rect 31502 7646 31554 7698
rect 31554 7646 31556 7698
rect 31500 7644 31556 7646
rect 31724 7308 31780 7364
rect 31836 6636 31892 6692
rect 31500 6578 31556 6580
rect 31500 6526 31502 6578
rect 31502 6526 31554 6578
rect 31554 6526 31556 6578
rect 31500 6524 31556 6526
rect 30716 6466 30772 6468
rect 30716 6414 30718 6466
rect 30718 6414 30770 6466
rect 30770 6414 30772 6466
rect 30716 6412 30772 6414
rect 30604 5740 30660 5796
rect 31388 5906 31444 5908
rect 31388 5854 31390 5906
rect 31390 5854 31442 5906
rect 31442 5854 31444 5906
rect 31388 5852 31444 5854
rect 30940 5740 30996 5796
rect 30940 5292 30996 5348
rect 30940 5122 30996 5124
rect 30940 5070 30942 5122
rect 30942 5070 30994 5122
rect 30994 5070 30996 5122
rect 30940 5068 30996 5070
rect 30380 4508 30436 4564
rect 31948 6188 32004 6244
rect 32508 7756 32564 7812
rect 33404 9660 33460 9716
rect 33852 9884 33908 9940
rect 33964 9660 34020 9716
rect 34972 13356 35028 13412
rect 35756 13858 35812 13860
rect 35756 13806 35758 13858
rect 35758 13806 35810 13858
rect 35810 13806 35812 13858
rect 35756 13804 35812 13806
rect 35308 13468 35364 13524
rect 34748 13186 34804 13188
rect 34748 13134 34750 13186
rect 34750 13134 34802 13186
rect 34802 13134 34804 13186
rect 34748 13132 34804 13134
rect 35532 13580 35588 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34972 13074 35028 13076
rect 34972 13022 34974 13074
rect 34974 13022 35026 13074
rect 35026 13022 35028 13074
rect 34972 13020 35028 13022
rect 34524 12796 34580 12852
rect 34300 12012 34356 12068
rect 35420 12850 35476 12852
rect 35420 12798 35422 12850
rect 35422 12798 35474 12850
rect 35474 12798 35476 12850
rect 35420 12796 35476 12798
rect 35644 13132 35700 13188
rect 35980 12850 36036 12852
rect 35980 12798 35982 12850
rect 35982 12798 36034 12850
rect 36034 12798 36036 12850
rect 35980 12796 36036 12798
rect 34636 11900 34692 11956
rect 35084 12012 35140 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35532 11452 35588 11508
rect 35532 11004 35588 11060
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34636 9772 34692 9828
rect 34188 9714 34244 9716
rect 34188 9662 34190 9714
rect 34190 9662 34242 9714
rect 34242 9662 34244 9714
rect 34188 9660 34244 9662
rect 34524 9100 34580 9156
rect 34076 8316 34132 8372
rect 32620 7420 32676 7476
rect 33628 7474 33684 7476
rect 33628 7422 33630 7474
rect 33630 7422 33682 7474
rect 33682 7422 33684 7474
rect 33628 7420 33684 7422
rect 33964 7980 34020 8036
rect 33964 7586 34020 7588
rect 33964 7534 33966 7586
rect 33966 7534 34018 7586
rect 34018 7534 34020 7586
rect 33964 7532 34020 7534
rect 34300 7474 34356 7476
rect 34300 7422 34302 7474
rect 34302 7422 34354 7474
rect 34354 7422 34356 7474
rect 34300 7420 34356 7422
rect 32508 6636 32564 6692
rect 32172 6412 32228 6468
rect 33628 6300 33684 6356
rect 35644 9826 35700 9828
rect 35644 9774 35646 9826
rect 35646 9774 35698 9826
rect 35698 9774 35700 9826
rect 35644 9772 35700 9774
rect 36988 19404 37044 19460
rect 37324 22258 37380 22260
rect 37324 22206 37326 22258
rect 37326 22206 37378 22258
rect 37378 22206 37380 22258
rect 37324 22204 37380 22206
rect 37772 19906 37828 19908
rect 37772 19854 37774 19906
rect 37774 19854 37826 19906
rect 37826 19854 37828 19906
rect 37772 19852 37828 19854
rect 37100 19180 37156 19236
rect 37100 18508 37156 18564
rect 37884 18844 37940 18900
rect 37212 18284 37268 18340
rect 37100 18060 37156 18116
rect 36428 13074 36484 13076
rect 36428 13022 36430 13074
rect 36430 13022 36482 13074
rect 36482 13022 36484 13074
rect 36428 13020 36484 13022
rect 37772 17836 37828 17892
rect 37772 15932 37828 15988
rect 37548 15708 37604 15764
rect 37212 13804 37268 13860
rect 37548 13858 37604 13860
rect 37548 13806 37550 13858
rect 37550 13806 37602 13858
rect 37602 13806 37604 13858
rect 37548 13804 37604 13806
rect 37100 12796 37156 12852
rect 36204 11676 36260 11732
rect 37660 11900 37716 11956
rect 35084 9042 35140 9044
rect 35084 8990 35086 9042
rect 35086 8990 35138 9042
rect 35138 8990 35140 9042
rect 35084 8988 35140 8990
rect 32172 5852 32228 5908
rect 32060 5628 32116 5684
rect 34972 8034 35028 8036
rect 34972 7982 34974 8034
rect 34974 7982 35026 8034
rect 35026 7982 35028 8034
rect 34972 7980 35028 7982
rect 34972 7196 35028 7252
rect 35532 9154 35588 9156
rect 35532 9102 35534 9154
rect 35534 9102 35586 9154
rect 35586 9102 35588 9154
rect 35532 9100 35588 9102
rect 36092 9826 36148 9828
rect 36092 9774 36094 9826
rect 36094 9774 36146 9826
rect 36146 9774 36148 9826
rect 36092 9772 36148 9774
rect 37100 9772 37156 9828
rect 36540 9714 36596 9716
rect 36540 9662 36542 9714
rect 36542 9662 36594 9714
rect 36594 9662 36596 9714
rect 36540 9660 36596 9662
rect 38444 23154 38500 23156
rect 38444 23102 38446 23154
rect 38446 23102 38498 23154
rect 38498 23102 38500 23154
rect 38444 23100 38500 23102
rect 38444 22204 38500 22260
rect 39228 23266 39284 23268
rect 39228 23214 39230 23266
rect 39230 23214 39282 23266
rect 39282 23214 39284 23266
rect 39228 23212 39284 23214
rect 38780 22428 38836 22484
rect 38668 19852 38724 19908
rect 38780 19740 38836 19796
rect 38780 19234 38836 19236
rect 38780 19182 38782 19234
rect 38782 19182 38834 19234
rect 38834 19182 38836 19234
rect 38780 19180 38836 19182
rect 38332 19010 38388 19012
rect 38332 18958 38334 19010
rect 38334 18958 38386 19010
rect 38386 18958 38388 19010
rect 38332 18956 38388 18958
rect 38556 17836 38612 17892
rect 38332 16322 38388 16324
rect 38332 16270 38334 16322
rect 38334 16270 38386 16322
rect 38386 16270 38388 16322
rect 38332 16268 38388 16270
rect 38108 15372 38164 15428
rect 38556 15314 38612 15316
rect 38556 15262 38558 15314
rect 38558 15262 38610 15314
rect 38610 15262 38612 15314
rect 38556 15260 38612 15262
rect 38332 14700 38388 14756
rect 37884 13804 37940 13860
rect 38444 13858 38500 13860
rect 38444 13806 38446 13858
rect 38446 13806 38498 13858
rect 38498 13806 38500 13858
rect 38444 13804 38500 13806
rect 38108 11900 38164 11956
rect 37884 11564 37940 11620
rect 39116 19292 39172 19348
rect 39788 19346 39844 19348
rect 39788 19294 39790 19346
rect 39790 19294 39842 19346
rect 39842 19294 39844 19346
rect 39788 19292 39844 19294
rect 39564 18732 39620 18788
rect 40124 25506 40180 25508
rect 40124 25454 40126 25506
rect 40126 25454 40178 25506
rect 40178 25454 40180 25506
rect 40124 25452 40180 25454
rect 40236 23996 40292 24052
rect 40348 21532 40404 21588
rect 40908 37154 40964 37156
rect 40908 37102 40910 37154
rect 40910 37102 40962 37154
rect 40962 37102 40964 37154
rect 40908 37100 40964 37102
rect 41244 37100 41300 37156
rect 41468 34354 41524 34356
rect 41468 34302 41470 34354
rect 41470 34302 41522 34354
rect 41522 34302 41524 34354
rect 41468 34300 41524 34302
rect 40684 26236 40740 26292
rect 40684 25452 40740 25508
rect 40572 25394 40628 25396
rect 40572 25342 40574 25394
rect 40574 25342 40626 25394
rect 40626 25342 40628 25394
rect 40572 25340 40628 25342
rect 41020 34130 41076 34132
rect 41020 34078 41022 34130
rect 41022 34078 41074 34130
rect 41074 34078 41076 34130
rect 41020 34076 41076 34078
rect 41244 34076 41300 34132
rect 41692 33516 41748 33572
rect 43372 40460 43428 40516
rect 42252 39228 42308 39284
rect 43036 37154 43092 37156
rect 43036 37102 43038 37154
rect 43038 37102 43090 37154
rect 43090 37102 43092 37154
rect 43036 37100 43092 37102
rect 42476 35698 42532 35700
rect 42476 35646 42478 35698
rect 42478 35646 42530 35698
rect 42530 35646 42532 35698
rect 42476 35644 42532 35646
rect 42364 34748 42420 34804
rect 42364 34354 42420 34356
rect 42364 34302 42366 34354
rect 42366 34302 42418 34354
rect 42418 34302 42420 34354
rect 42364 34300 42420 34302
rect 42028 34130 42084 34132
rect 42028 34078 42030 34130
rect 42030 34078 42082 34130
rect 42082 34078 42084 34130
rect 42028 34076 42084 34078
rect 41916 33964 41972 34020
rect 41132 27858 41188 27860
rect 41132 27806 41134 27858
rect 41134 27806 41186 27858
rect 41186 27806 41188 27858
rect 41132 27804 41188 27806
rect 40908 27074 40964 27076
rect 40908 27022 40910 27074
rect 40910 27022 40962 27074
rect 40962 27022 40964 27074
rect 40908 27020 40964 27022
rect 41132 26290 41188 26292
rect 41132 26238 41134 26290
rect 41134 26238 41186 26290
rect 41186 26238 41188 26290
rect 41132 26236 41188 26238
rect 41020 26066 41076 26068
rect 41020 26014 41022 26066
rect 41022 26014 41074 26066
rect 41074 26014 41076 26066
rect 41020 26012 41076 26014
rect 41132 24834 41188 24836
rect 41132 24782 41134 24834
rect 41134 24782 41186 24834
rect 41186 24782 41188 24834
rect 41132 24780 41188 24782
rect 42364 33516 42420 33572
rect 42364 33180 42420 33236
rect 42028 32284 42084 32340
rect 43932 42364 43988 42420
rect 44940 43426 44996 43428
rect 44940 43374 44942 43426
rect 44942 43374 44994 43426
rect 44994 43374 44996 43426
rect 44940 43372 44996 43374
rect 44268 41244 44324 41300
rect 44156 40962 44212 40964
rect 44156 40910 44158 40962
rect 44158 40910 44210 40962
rect 44210 40910 44212 40962
rect 44156 40908 44212 40910
rect 44492 40908 44548 40964
rect 45388 43372 45444 43428
rect 45164 42530 45220 42532
rect 45164 42478 45166 42530
rect 45166 42478 45218 42530
rect 45218 42478 45220 42530
rect 45164 42476 45220 42478
rect 45612 42978 45668 42980
rect 45612 42926 45614 42978
rect 45614 42926 45666 42978
rect 45666 42926 45668 42978
rect 45612 42924 45668 42926
rect 45612 42700 45668 42756
rect 45500 42364 45556 42420
rect 47404 49586 47460 49588
rect 47404 49534 47406 49586
rect 47406 49534 47458 49586
rect 47458 49534 47460 49586
rect 47404 49532 47460 49534
rect 47740 47180 47796 47236
rect 47628 46396 47684 46452
rect 48412 45890 48468 45892
rect 48412 45838 48414 45890
rect 48414 45838 48466 45890
rect 48466 45838 48468 45890
rect 48412 45836 48468 45838
rect 48076 45666 48132 45668
rect 48076 45614 48078 45666
rect 48078 45614 48130 45666
rect 48130 45614 48132 45666
rect 48076 45612 48132 45614
rect 48300 45330 48356 45332
rect 48300 45278 48302 45330
rect 48302 45278 48354 45330
rect 48354 45278 48356 45330
rect 48300 45276 48356 45278
rect 46620 43372 46676 43428
rect 46844 43372 46900 43428
rect 46620 42754 46676 42756
rect 46620 42702 46622 42754
rect 46622 42702 46674 42754
rect 46674 42702 46676 42754
rect 46620 42700 46676 42702
rect 45948 42476 46004 42532
rect 46396 42530 46452 42532
rect 46396 42478 46398 42530
rect 46398 42478 46450 42530
rect 46450 42478 46452 42530
rect 46396 42476 46452 42478
rect 48188 43426 48244 43428
rect 48188 43374 48190 43426
rect 48190 43374 48242 43426
rect 48242 43374 48244 43426
rect 48188 43372 48244 43374
rect 45724 41916 45780 41972
rect 46844 41916 46900 41972
rect 45164 41298 45220 41300
rect 45164 41246 45166 41298
rect 45166 41246 45218 41298
rect 45218 41246 45220 41298
rect 45164 41244 45220 41246
rect 44604 39788 44660 39844
rect 43820 39618 43876 39620
rect 43820 39566 43822 39618
rect 43822 39566 43874 39618
rect 43874 39566 43876 39618
rect 43820 39564 43876 39566
rect 44268 39506 44324 39508
rect 44268 39454 44270 39506
rect 44270 39454 44322 39506
rect 44322 39454 44324 39506
rect 44268 39452 44324 39454
rect 45164 40908 45220 40964
rect 49756 60956 49812 61012
rect 48860 58716 48916 58772
rect 49532 60620 49588 60676
rect 50652 63420 50708 63476
rect 50764 63138 50820 63140
rect 50764 63086 50766 63138
rect 50766 63086 50818 63138
rect 50818 63086 50820 63138
rect 50764 63084 50820 63086
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 51772 65324 51828 65380
rect 50988 61852 51044 61908
rect 51100 63196 51156 63252
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50428 60956 50484 61012
rect 50988 61010 51044 61012
rect 50988 60958 50990 61010
rect 50990 60958 51042 61010
rect 51042 60958 51044 61010
rect 50988 60956 51044 60958
rect 50204 60844 50260 60900
rect 49756 60674 49812 60676
rect 49756 60622 49758 60674
rect 49758 60622 49810 60674
rect 49810 60622 49812 60674
rect 49756 60620 49812 60622
rect 49532 59276 49588 59332
rect 48748 56194 48804 56196
rect 48748 56142 48750 56194
rect 48750 56142 48802 56194
rect 48802 56142 48804 56194
rect 48748 56140 48804 56142
rect 50988 60620 51044 60676
rect 51324 63922 51380 63924
rect 51324 63870 51326 63922
rect 51326 63870 51378 63922
rect 51378 63870 51380 63922
rect 51324 63868 51380 63870
rect 52108 64428 52164 64484
rect 51660 62242 51716 62244
rect 51660 62190 51662 62242
rect 51662 62190 51714 62242
rect 51714 62190 51716 62242
rect 51660 62188 51716 62190
rect 51436 60956 51492 61012
rect 51212 60172 51268 60228
rect 51660 60732 51716 60788
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50428 59442 50484 59444
rect 50428 59390 50430 59442
rect 50430 59390 50482 59442
rect 50482 59390 50484 59442
rect 50428 59388 50484 59390
rect 49420 57372 49476 57428
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 49980 56306 50036 56308
rect 49980 56254 49982 56306
rect 49982 56254 50034 56306
rect 50034 56254 50036 56306
rect 49980 56252 50036 56254
rect 50316 56252 50372 56308
rect 51100 57538 51156 57540
rect 51100 57486 51102 57538
rect 51102 57486 51154 57538
rect 51154 57486 51156 57538
rect 51100 57484 51156 57486
rect 50316 56082 50372 56084
rect 50316 56030 50318 56082
rect 50318 56030 50370 56082
rect 50370 56030 50372 56082
rect 50316 56028 50372 56030
rect 49308 55132 49364 55188
rect 49980 55186 50036 55188
rect 49980 55134 49982 55186
rect 49982 55134 50034 55186
rect 50034 55134 50036 55186
rect 49980 55132 50036 55134
rect 49532 55074 49588 55076
rect 49532 55022 49534 55074
rect 49534 55022 49586 55074
rect 49586 55022 49588 55074
rect 49532 55020 49588 55022
rect 49196 54572 49252 54628
rect 50316 54460 50372 54516
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50876 56252 50932 56308
rect 50428 55020 50484 55076
rect 48748 51548 48804 51604
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50876 54514 50932 54516
rect 50876 54462 50878 54514
rect 50878 54462 50930 54514
rect 50930 54462 50932 54514
rect 50876 54460 50932 54462
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50988 53004 51044 53060
rect 51436 59388 51492 59444
rect 54124 65378 54180 65380
rect 54124 65326 54126 65378
rect 54126 65326 54178 65378
rect 54178 65326 54180 65378
rect 54124 65324 54180 65326
rect 54908 65324 54964 65380
rect 52780 64482 52836 64484
rect 52780 64430 52782 64482
rect 52782 64430 52834 64482
rect 52834 64430 52836 64482
rect 52780 64428 52836 64430
rect 54908 64428 54964 64484
rect 54236 64092 54292 64148
rect 53004 63250 53060 63252
rect 53004 63198 53006 63250
rect 53006 63198 53058 63250
rect 53058 63198 53060 63250
rect 53004 63196 53060 63198
rect 52108 62578 52164 62580
rect 52108 62526 52110 62578
rect 52110 62526 52162 62578
rect 52162 62526 52164 62578
rect 52108 62524 52164 62526
rect 52444 62466 52500 62468
rect 52444 62414 52446 62466
rect 52446 62414 52498 62466
rect 52498 62414 52500 62466
rect 52444 62412 52500 62414
rect 52892 62242 52948 62244
rect 52892 62190 52894 62242
rect 52894 62190 52946 62242
rect 52946 62190 52948 62242
rect 52892 62188 52948 62190
rect 53900 63250 53956 63252
rect 53900 63198 53902 63250
rect 53902 63198 53954 63250
rect 53954 63198 53956 63250
rect 53900 63196 53956 63198
rect 53228 62412 53284 62468
rect 53004 60786 53060 60788
rect 53004 60734 53006 60786
rect 53006 60734 53058 60786
rect 53058 60734 53060 60786
rect 53004 60732 53060 60734
rect 52780 60620 52836 60676
rect 54124 62188 54180 62244
rect 54572 64146 54628 64148
rect 54572 64094 54574 64146
rect 54574 64094 54626 64146
rect 54626 64094 54628 64146
rect 54572 64092 54628 64094
rect 56028 66498 56084 66500
rect 56028 66446 56030 66498
rect 56030 66446 56082 66498
rect 56082 66446 56084 66498
rect 56028 66444 56084 66446
rect 55468 65378 55524 65380
rect 55468 65326 55470 65378
rect 55470 65326 55522 65378
rect 55522 65326 55524 65378
rect 55468 65324 55524 65326
rect 55356 65100 55412 65156
rect 55244 64876 55300 64932
rect 55244 64034 55300 64036
rect 55244 63982 55246 64034
rect 55246 63982 55298 64034
rect 55298 63982 55300 64034
rect 55244 63980 55300 63982
rect 55132 63756 55188 63812
rect 55020 63420 55076 63476
rect 54348 60844 54404 60900
rect 54460 60956 54516 61012
rect 53340 60508 53396 60564
rect 54684 60508 54740 60564
rect 51884 60172 51940 60228
rect 55244 63250 55300 63252
rect 55244 63198 55246 63250
rect 55246 63198 55298 63250
rect 55298 63198 55300 63250
rect 55244 63196 55300 63198
rect 55020 62524 55076 62580
rect 58156 66108 58212 66164
rect 57596 65490 57652 65492
rect 57596 65438 57598 65490
rect 57598 65438 57650 65490
rect 57650 65438 57652 65490
rect 57596 65436 57652 65438
rect 57148 65100 57204 65156
rect 55804 64034 55860 64036
rect 55804 63982 55806 64034
rect 55806 63982 55858 64034
rect 55858 63982 55860 64034
rect 55804 63980 55860 63982
rect 55580 62524 55636 62580
rect 55468 61570 55524 61572
rect 55468 61518 55470 61570
rect 55470 61518 55522 61570
rect 55522 61518 55524 61570
rect 55468 61516 55524 61518
rect 51436 57650 51492 57652
rect 51436 57598 51438 57650
rect 51438 57598 51490 57650
rect 51490 57598 51492 57650
rect 51436 57596 51492 57598
rect 51436 56028 51492 56084
rect 51324 54684 51380 54740
rect 52108 60002 52164 60004
rect 52108 59950 52110 60002
rect 52110 59950 52162 60002
rect 52162 59950 52164 60002
rect 52108 59948 52164 59950
rect 53340 59948 53396 60004
rect 52556 58268 52612 58324
rect 53004 58268 53060 58324
rect 51996 56476 52052 56532
rect 52780 56476 52836 56532
rect 51884 56028 51940 56084
rect 55244 60956 55300 61012
rect 54236 59948 54292 60004
rect 54908 59948 54964 60004
rect 54684 59442 54740 59444
rect 54684 59390 54686 59442
rect 54686 59390 54738 59442
rect 54738 59390 54740 59442
rect 54684 59388 54740 59390
rect 56364 63756 56420 63812
rect 55916 63698 55972 63700
rect 55916 63646 55918 63698
rect 55918 63646 55970 63698
rect 55970 63646 55972 63698
rect 55916 63644 55972 63646
rect 56700 60956 56756 61012
rect 55804 60898 55860 60900
rect 55804 60846 55806 60898
rect 55806 60846 55858 60898
rect 55858 60846 55860 60898
rect 55804 60844 55860 60846
rect 56588 60898 56644 60900
rect 56588 60846 56590 60898
rect 56590 60846 56642 60898
rect 56642 60846 56644 60898
rect 56588 60844 56644 60846
rect 57372 63644 57428 63700
rect 58156 65490 58212 65492
rect 58156 65438 58158 65490
rect 58158 65438 58210 65490
rect 58210 65438 58212 65490
rect 58156 65436 58212 65438
rect 56700 60508 56756 60564
rect 57148 60620 57204 60676
rect 56700 59442 56756 59444
rect 56700 59390 56702 59442
rect 56702 59390 56754 59442
rect 56754 59390 56756 59442
rect 56700 59388 56756 59390
rect 55692 59164 55748 59220
rect 56812 59164 56868 59220
rect 51884 54738 51940 54740
rect 51884 54686 51886 54738
rect 51886 54686 51938 54738
rect 51938 54686 51940 54738
rect 51884 54684 51940 54686
rect 51660 54514 51716 54516
rect 51660 54462 51662 54514
rect 51662 54462 51714 54514
rect 51714 54462 51716 54514
rect 51660 54460 51716 54462
rect 51660 53900 51716 53956
rect 52668 53954 52724 53956
rect 52668 53902 52670 53954
rect 52670 53902 52722 53954
rect 52722 53902 52724 53954
rect 52668 53900 52724 53902
rect 52892 55074 52948 55076
rect 52892 55022 52894 55074
rect 52894 55022 52946 55074
rect 52946 55022 52948 55074
rect 52892 55020 52948 55022
rect 53116 54684 53172 54740
rect 53788 55020 53844 55076
rect 52780 53788 52836 53844
rect 53004 53842 53060 53844
rect 53004 53790 53006 53842
rect 53006 53790 53058 53842
rect 53058 53790 53060 53842
rect 53004 53788 53060 53790
rect 51660 53506 51716 53508
rect 51660 53454 51662 53506
rect 51662 53454 51714 53506
rect 51714 53454 51716 53506
rect 51660 53452 51716 53454
rect 51548 53116 51604 53172
rect 51660 53004 51716 53060
rect 51324 52444 51380 52500
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50764 49810 50820 49812
rect 50764 49758 50766 49810
rect 50766 49758 50818 49810
rect 50818 49758 50820 49810
rect 50764 49756 50820 49758
rect 48860 49532 48916 49588
rect 49196 48300 49252 48356
rect 48860 47180 48916 47236
rect 48748 46786 48804 46788
rect 48748 46734 48750 46786
rect 48750 46734 48802 46786
rect 48802 46734 48804 46786
rect 48748 46732 48804 46734
rect 48748 45330 48804 45332
rect 48748 45278 48750 45330
rect 48750 45278 48802 45330
rect 48802 45278 48804 45330
rect 48748 45276 48804 45278
rect 45836 39842 45892 39844
rect 45836 39790 45838 39842
rect 45838 39790 45890 39842
rect 45890 39790 45892 39842
rect 45836 39788 45892 39790
rect 48748 39788 48804 39844
rect 45052 39506 45108 39508
rect 45052 39454 45054 39506
rect 45054 39454 45106 39506
rect 45106 39454 45108 39506
rect 45052 39452 45108 39454
rect 47404 39618 47460 39620
rect 47404 39566 47406 39618
rect 47406 39566 47458 39618
rect 47458 39566 47460 39618
rect 47404 39564 47460 39566
rect 45724 39506 45780 39508
rect 45724 39454 45726 39506
rect 45726 39454 45778 39506
rect 45778 39454 45780 39506
rect 45724 39452 45780 39454
rect 48748 39228 48804 39284
rect 42700 34412 42756 34468
rect 46172 38722 46228 38724
rect 46172 38670 46174 38722
rect 46174 38670 46226 38722
rect 46226 38670 46228 38722
rect 46172 38668 46228 38670
rect 49644 47964 49700 48020
rect 49308 46674 49364 46676
rect 49308 46622 49310 46674
rect 49310 46622 49362 46674
rect 49362 46622 49364 46674
rect 49308 46620 49364 46622
rect 49308 45724 49364 45780
rect 49084 45218 49140 45220
rect 49084 45166 49086 45218
rect 49086 45166 49138 45218
rect 49138 45166 49140 45218
rect 49084 45164 49140 45166
rect 49196 41970 49252 41972
rect 49196 41918 49198 41970
rect 49198 41918 49250 41970
rect 49250 41918 49252 41970
rect 49196 41916 49252 41918
rect 49084 39788 49140 39844
rect 48972 39228 49028 39284
rect 45724 38108 45780 38164
rect 45052 34972 45108 35028
rect 46396 38162 46452 38164
rect 46396 38110 46398 38162
rect 46398 38110 46450 38162
rect 46450 38110 46452 38162
rect 46396 38108 46452 38110
rect 46060 37996 46116 38052
rect 46620 37884 46676 37940
rect 43820 34802 43876 34804
rect 43820 34750 43822 34802
rect 43822 34750 43874 34802
rect 43874 34750 43876 34802
rect 43820 34748 43876 34750
rect 43596 34412 43652 34468
rect 44268 34748 44324 34804
rect 43260 33292 43316 33348
rect 44492 34412 44548 34468
rect 44604 34130 44660 34132
rect 44604 34078 44606 34130
rect 44606 34078 44658 34130
rect 44658 34078 44660 34130
rect 44604 34076 44660 34078
rect 45052 34076 45108 34132
rect 43372 33180 43428 33236
rect 43596 32450 43652 32452
rect 43596 32398 43598 32450
rect 43598 32398 43650 32450
rect 43650 32398 43652 32450
rect 43596 32396 43652 32398
rect 41468 29260 41524 29316
rect 44044 32450 44100 32452
rect 44044 32398 44046 32450
rect 44046 32398 44098 32450
rect 44098 32398 44100 32450
rect 44044 32396 44100 32398
rect 48524 37938 48580 37940
rect 48524 37886 48526 37938
rect 48526 37886 48578 37938
rect 48578 37886 48580 37938
rect 48524 37884 48580 37886
rect 45500 35698 45556 35700
rect 45500 35646 45502 35698
rect 45502 35646 45554 35698
rect 45554 35646 45556 35698
rect 45500 35644 45556 35646
rect 45500 35026 45556 35028
rect 45500 34974 45502 35026
rect 45502 34974 45554 35026
rect 45554 34974 45556 35026
rect 45500 34972 45556 34974
rect 45724 34130 45780 34132
rect 45724 34078 45726 34130
rect 45726 34078 45778 34130
rect 45778 34078 45780 34130
rect 45724 34076 45780 34078
rect 48860 34972 48916 35028
rect 47740 34300 47796 34356
rect 45948 33068 46004 33124
rect 46732 32562 46788 32564
rect 46732 32510 46734 32562
rect 46734 32510 46786 32562
rect 46786 32510 46788 32562
rect 46732 32508 46788 32510
rect 44268 31778 44324 31780
rect 44268 31726 44270 31778
rect 44270 31726 44322 31778
rect 44322 31726 44324 31778
rect 44268 31724 44324 31726
rect 42364 30156 42420 30212
rect 41916 29932 41972 29988
rect 41804 29148 41860 29204
rect 42812 29202 42868 29204
rect 42812 29150 42814 29202
rect 42814 29150 42866 29202
rect 42866 29150 42868 29202
rect 42812 29148 42868 29150
rect 43372 28418 43428 28420
rect 43372 28366 43374 28418
rect 43374 28366 43426 28418
rect 43426 28366 43428 28418
rect 43372 28364 43428 28366
rect 44044 28364 44100 28420
rect 41916 27804 41972 27860
rect 41916 26908 41972 26964
rect 44380 28700 44436 28756
rect 41468 26402 41524 26404
rect 41468 26350 41470 26402
rect 41470 26350 41522 26402
rect 41522 26350 41524 26402
rect 41468 26348 41524 26350
rect 41468 25394 41524 25396
rect 41468 25342 41470 25394
rect 41470 25342 41522 25394
rect 41522 25342 41524 25394
rect 41468 25340 41524 25342
rect 41356 25228 41412 25284
rect 41244 24668 41300 24724
rect 40460 20188 40516 20244
rect 40348 20130 40404 20132
rect 40348 20078 40350 20130
rect 40350 20078 40402 20130
rect 40402 20078 40404 20130
rect 40348 20076 40404 20078
rect 40236 18844 40292 18900
rect 40236 18284 40292 18340
rect 40684 22482 40740 22484
rect 40684 22430 40686 22482
rect 40686 22430 40738 22482
rect 40738 22430 40740 22482
rect 40684 22428 40740 22430
rect 41020 23378 41076 23380
rect 41020 23326 41022 23378
rect 41022 23326 41074 23378
rect 41074 23326 41076 23378
rect 41020 23324 41076 23326
rect 40908 21756 40964 21812
rect 41468 22204 41524 22260
rect 41468 21586 41524 21588
rect 41468 21534 41470 21586
rect 41470 21534 41522 21586
rect 41522 21534 41524 21586
rect 41468 21532 41524 21534
rect 42588 26852 42644 26908
rect 41916 26178 41972 26180
rect 41916 26126 41918 26178
rect 41918 26126 41970 26178
rect 41970 26126 41972 26178
rect 41916 26124 41972 26126
rect 41916 25340 41972 25396
rect 42476 25282 42532 25284
rect 42476 25230 42478 25282
rect 42478 25230 42530 25282
rect 42530 25230 42532 25282
rect 42476 25228 42532 25230
rect 43932 26850 43988 26852
rect 43932 26798 43934 26850
rect 43934 26798 43986 26850
rect 43986 26798 43988 26850
rect 43932 26796 43988 26798
rect 42140 25116 42196 25172
rect 41804 24610 41860 24612
rect 41804 24558 41806 24610
rect 41806 24558 41858 24610
rect 41858 24558 41860 24610
rect 41804 24556 41860 24558
rect 42700 24556 42756 24612
rect 42700 23548 42756 23604
rect 41916 23436 41972 23492
rect 42476 23436 42532 23492
rect 42252 22428 42308 22484
rect 42028 22258 42084 22260
rect 42028 22206 42030 22258
rect 42030 22206 42082 22258
rect 42082 22206 42084 22258
rect 42028 22204 42084 22206
rect 41020 19906 41076 19908
rect 41020 19854 41022 19906
rect 41022 19854 41074 19906
rect 41074 19854 41076 19906
rect 41020 19852 41076 19854
rect 40908 19740 40964 19796
rect 40572 18060 40628 18116
rect 40012 17948 40068 18004
rect 39788 17724 39844 17780
rect 40684 17778 40740 17780
rect 40684 17726 40686 17778
rect 40686 17726 40738 17778
rect 40738 17726 40740 17778
rect 40684 17724 40740 17726
rect 40572 17612 40628 17668
rect 39676 15820 39732 15876
rect 39228 15426 39284 15428
rect 39228 15374 39230 15426
rect 39230 15374 39282 15426
rect 39282 15374 39284 15426
rect 39228 15372 39284 15374
rect 39676 15314 39732 15316
rect 39676 15262 39678 15314
rect 39678 15262 39730 15314
rect 39730 15262 39732 15314
rect 39676 15260 39732 15262
rect 39116 13916 39172 13972
rect 39564 14418 39620 14420
rect 39564 14366 39566 14418
rect 39566 14366 39618 14418
rect 39618 14366 39620 14418
rect 39564 14364 39620 14366
rect 38780 12962 38836 12964
rect 38780 12910 38782 12962
rect 38782 12910 38834 12962
rect 38834 12910 38836 12962
rect 38780 12908 38836 12910
rect 38780 11900 38836 11956
rect 39116 13522 39172 13524
rect 39116 13470 39118 13522
rect 39118 13470 39170 13522
rect 39170 13470 39172 13522
rect 39116 13468 39172 13470
rect 40012 14700 40068 14756
rect 40012 13468 40068 13524
rect 39676 12962 39732 12964
rect 39676 12910 39678 12962
rect 39678 12910 39730 12962
rect 39730 12910 39732 12962
rect 39676 12908 39732 12910
rect 39116 12178 39172 12180
rect 39116 12126 39118 12178
rect 39118 12126 39170 12178
rect 39170 12126 39172 12178
rect 39116 12124 39172 12126
rect 38668 11564 38724 11620
rect 38332 11506 38388 11508
rect 38332 11454 38334 11506
rect 38334 11454 38386 11506
rect 38386 11454 38388 11506
rect 38332 11452 38388 11454
rect 39452 11452 39508 11508
rect 40236 12348 40292 12404
rect 40236 12012 40292 12068
rect 39004 10780 39060 10836
rect 37324 9436 37380 9492
rect 35868 8988 35924 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36316 8204 36372 8260
rect 35532 7980 35588 8036
rect 35644 7586 35700 7588
rect 35644 7534 35646 7586
rect 35646 7534 35698 7586
rect 35698 7534 35700 7586
rect 35644 7532 35700 7534
rect 34636 5180 34692 5236
rect 32060 5068 32116 5124
rect 35420 7474 35476 7476
rect 35420 7422 35422 7474
rect 35422 7422 35474 7474
rect 35474 7422 35476 7474
rect 35420 7420 35476 7422
rect 36092 8034 36148 8036
rect 36092 7982 36094 8034
rect 36094 7982 36146 8034
rect 36146 7982 36148 8034
rect 36092 7980 36148 7982
rect 36316 7868 36372 7924
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35980 7250 36036 7252
rect 35980 7198 35982 7250
rect 35982 7198 36034 7250
rect 36034 7198 36036 7250
rect 35980 7196 36036 7198
rect 36204 7196 36260 7252
rect 36428 7586 36484 7588
rect 36428 7534 36430 7586
rect 36430 7534 36482 7586
rect 36482 7534 36484 7586
rect 36428 7532 36484 7534
rect 36764 7196 36820 7252
rect 36428 7084 36484 7140
rect 39228 9266 39284 9268
rect 39228 9214 39230 9266
rect 39230 9214 39282 9266
rect 39282 9214 39284 9266
rect 39228 9212 39284 9214
rect 37660 9154 37716 9156
rect 37660 9102 37662 9154
rect 37662 9102 37714 9154
rect 37714 9102 37716 9154
rect 37660 9100 37716 9102
rect 40236 10780 40292 10836
rect 39788 9100 39844 9156
rect 39004 8146 39060 8148
rect 39004 8094 39006 8146
rect 39006 8094 39058 8146
rect 39058 8094 39060 8146
rect 39004 8092 39060 8094
rect 38892 7868 38948 7924
rect 38108 7474 38164 7476
rect 38108 7422 38110 7474
rect 38110 7422 38162 7474
rect 38162 7422 38164 7474
rect 38108 7420 38164 7422
rect 38668 7474 38724 7476
rect 38668 7422 38670 7474
rect 38670 7422 38722 7474
rect 38722 7422 38724 7474
rect 38668 7420 38724 7422
rect 38220 7308 38276 7364
rect 37548 7084 37604 7140
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5234 35700 5236
rect 35644 5182 35646 5234
rect 35646 5182 35698 5234
rect 35698 5182 35700 5234
rect 35644 5180 35700 5182
rect 39340 7308 39396 7364
rect 38780 6972 38836 7028
rect 38556 6636 38612 6692
rect 39340 6524 39396 6580
rect 37660 5292 37716 5348
rect 39676 8146 39732 8148
rect 39676 8094 39678 8146
rect 39678 8094 39730 8146
rect 39730 8094 39732 8146
rect 39676 8092 39732 8094
rect 40460 10332 40516 10388
rect 40348 9714 40404 9716
rect 40348 9662 40350 9714
rect 40350 9662 40402 9714
rect 40402 9662 40404 9714
rect 40348 9660 40404 9662
rect 41244 20130 41300 20132
rect 41244 20078 41246 20130
rect 41246 20078 41298 20130
rect 41298 20078 41300 20130
rect 41244 20076 41300 20078
rect 41468 20018 41524 20020
rect 41468 19966 41470 20018
rect 41470 19966 41522 20018
rect 41522 19966 41524 20018
rect 41468 19964 41524 19966
rect 42140 19964 42196 20020
rect 41916 19740 41972 19796
rect 41244 18732 41300 18788
rect 41356 18450 41412 18452
rect 41356 18398 41358 18450
rect 41358 18398 41410 18450
rect 41410 18398 41412 18450
rect 41356 18396 41412 18398
rect 41468 17836 41524 17892
rect 43260 25228 43316 25284
rect 42924 23324 42980 23380
rect 43036 24444 43092 24500
rect 43148 24556 43204 24612
rect 42588 19906 42644 19908
rect 42588 19854 42590 19906
rect 42590 19854 42642 19906
rect 42642 19854 42644 19906
rect 42588 19852 42644 19854
rect 42364 19404 42420 19460
rect 42028 19010 42084 19012
rect 42028 18958 42030 19010
rect 42030 18958 42082 19010
rect 42082 18958 42084 19010
rect 42028 18956 42084 18958
rect 42364 18620 42420 18676
rect 42588 18450 42644 18452
rect 42588 18398 42590 18450
rect 42590 18398 42642 18450
rect 42642 18398 42644 18450
rect 42588 18396 42644 18398
rect 41804 18284 41860 18340
rect 42364 18172 42420 18228
rect 41692 17612 41748 17668
rect 40908 15708 40964 15764
rect 41020 16268 41076 16324
rect 41020 15260 41076 15316
rect 40908 14418 40964 14420
rect 40908 14366 40910 14418
rect 40910 14366 40962 14418
rect 40962 14366 40964 14418
rect 40908 14364 40964 14366
rect 41132 15820 41188 15876
rect 41916 15314 41972 15316
rect 41916 15262 41918 15314
rect 41918 15262 41970 15314
rect 41970 15262 41972 15314
rect 41916 15260 41972 15262
rect 41468 14642 41524 14644
rect 41468 14590 41470 14642
rect 41470 14590 41522 14642
rect 41522 14590 41524 14642
rect 41468 14588 41524 14590
rect 41692 15036 41748 15092
rect 41916 14530 41972 14532
rect 41916 14478 41918 14530
rect 41918 14478 41970 14530
rect 41970 14478 41972 14530
rect 41916 14476 41972 14478
rect 41132 14252 41188 14308
rect 41468 14252 41524 14308
rect 41916 13916 41972 13972
rect 42812 15036 42868 15092
rect 42588 14588 42644 14644
rect 42700 14306 42756 14308
rect 42700 14254 42702 14306
rect 42702 14254 42754 14306
rect 42754 14254 42756 14306
rect 42700 14252 42756 14254
rect 42140 13634 42196 13636
rect 42140 13582 42142 13634
rect 42142 13582 42194 13634
rect 42194 13582 42196 13634
rect 42140 13580 42196 13582
rect 41132 12796 41188 12852
rect 42028 12850 42084 12852
rect 42028 12798 42030 12850
rect 42030 12798 42082 12850
rect 42082 12798 42084 12850
rect 42028 12796 42084 12798
rect 43148 18620 43204 18676
rect 43036 14700 43092 14756
rect 43036 14476 43092 14532
rect 43708 25228 43764 25284
rect 43484 24610 43540 24612
rect 43484 24558 43486 24610
rect 43486 24558 43538 24610
rect 43538 24558 43540 24610
rect 43484 24556 43540 24558
rect 43596 23548 43652 23604
rect 43372 23436 43428 23492
rect 43372 22540 43428 22596
rect 43260 13970 43316 13972
rect 43260 13918 43262 13970
rect 43262 13918 43314 13970
rect 43314 13918 43316 13970
rect 43260 13916 43316 13918
rect 43708 22204 43764 22260
rect 43596 18172 43652 18228
rect 44268 26962 44324 26964
rect 44268 26910 44270 26962
rect 44270 26910 44322 26962
rect 44322 26910 44324 26962
rect 44268 26908 44324 26910
rect 43932 26012 43988 26068
rect 44380 25788 44436 25844
rect 44380 25228 44436 25284
rect 44156 23436 44212 23492
rect 44156 22482 44212 22484
rect 44156 22430 44158 22482
rect 44158 22430 44210 22482
rect 44210 22430 44212 22482
rect 44156 22428 44212 22430
rect 43932 18172 43988 18228
rect 44380 19852 44436 19908
rect 44380 19292 44436 19348
rect 44268 17836 44324 17892
rect 44156 16716 44212 16772
rect 47404 32562 47460 32564
rect 47404 32510 47406 32562
rect 47406 32510 47458 32562
rect 47458 32510 47460 32562
rect 47404 32508 47460 32510
rect 45388 31890 45444 31892
rect 45388 31838 45390 31890
rect 45390 31838 45442 31890
rect 45442 31838 45444 31890
rect 45388 31836 45444 31838
rect 45164 31724 45220 31780
rect 45276 30156 45332 30212
rect 47516 31666 47572 31668
rect 47516 31614 47518 31666
rect 47518 31614 47570 31666
rect 47570 31614 47572 31666
rect 47516 31612 47572 31614
rect 45612 30156 45668 30212
rect 46956 30322 47012 30324
rect 46956 30270 46958 30322
rect 46958 30270 47010 30322
rect 47010 30270 47012 30322
rect 46956 30268 47012 30270
rect 46508 29260 46564 29316
rect 45276 28754 45332 28756
rect 45276 28702 45278 28754
rect 45278 28702 45330 28754
rect 45330 28702 45332 28754
rect 45276 28700 45332 28702
rect 45052 26908 45108 26964
rect 44828 26796 44884 26852
rect 44940 26012 44996 26068
rect 46396 26348 46452 26404
rect 45164 25452 45220 25508
rect 44828 25394 44884 25396
rect 44828 25342 44830 25394
rect 44830 25342 44882 25394
rect 44882 25342 44884 25394
rect 44828 25340 44884 25342
rect 45836 26236 45892 26292
rect 45164 24668 45220 24724
rect 44828 24444 44884 24500
rect 44604 23996 44660 24052
rect 45276 24610 45332 24612
rect 45276 24558 45278 24610
rect 45278 24558 45330 24610
rect 45330 24558 45332 24610
rect 45276 24556 45332 24558
rect 48972 33628 49028 33684
rect 49532 45836 49588 45892
rect 50876 49026 50932 49028
rect 50876 48974 50878 49026
rect 50878 48974 50930 49026
rect 50930 48974 50932 49026
rect 50876 48972 50932 48974
rect 49868 47404 49924 47460
rect 49756 47234 49812 47236
rect 49756 47182 49758 47234
rect 49758 47182 49810 47234
rect 49810 47182 49812 47234
rect 49756 47180 49812 47182
rect 49756 46674 49812 46676
rect 49756 46622 49758 46674
rect 49758 46622 49810 46674
rect 49810 46622 49812 46674
rect 49756 46620 49812 46622
rect 51100 51100 51156 51156
rect 52780 53506 52836 53508
rect 52780 53454 52782 53506
rect 52782 53454 52834 53506
rect 52834 53454 52836 53506
rect 52780 53452 52836 53454
rect 53676 53452 53732 53508
rect 53900 55468 53956 55524
rect 53340 52220 53396 52276
rect 53228 52108 53284 52164
rect 51772 51154 51828 51156
rect 51772 51102 51774 51154
rect 51774 51102 51826 51154
rect 51826 51102 51828 51154
rect 51772 51100 51828 51102
rect 52444 51378 52500 51380
rect 52444 51326 52446 51378
rect 52446 51326 52498 51378
rect 52498 51326 52500 51378
rect 52444 51324 52500 51326
rect 51212 50652 51268 50708
rect 51212 49868 51268 49924
rect 51100 49756 51156 49812
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 51660 49922 51716 49924
rect 51660 49870 51662 49922
rect 51662 49870 51714 49922
rect 51714 49870 51716 49922
rect 51660 49868 51716 49870
rect 53228 50764 53284 50820
rect 52668 49810 52724 49812
rect 52668 49758 52670 49810
rect 52670 49758 52722 49810
rect 52722 49758 52724 49810
rect 52668 49756 52724 49758
rect 51548 49026 51604 49028
rect 51548 48974 51550 49026
rect 51550 48974 51602 49026
rect 51602 48974 51604 49026
rect 51548 48972 51604 48974
rect 49980 47180 50036 47236
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50540 46674 50596 46676
rect 50540 46622 50542 46674
rect 50542 46622 50594 46674
rect 50594 46622 50596 46674
rect 50540 46620 50596 46622
rect 50316 46508 50372 46564
rect 49980 45778 50036 45780
rect 49980 45726 49982 45778
rect 49982 45726 50034 45778
rect 50034 45726 50036 45778
rect 49980 45724 50036 45726
rect 49980 45106 50036 45108
rect 49980 45054 49982 45106
rect 49982 45054 50034 45106
rect 50034 45054 50036 45106
rect 49980 45052 50036 45054
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50428 45164 50484 45220
rect 50988 45164 51044 45220
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50204 42642 50260 42644
rect 50204 42590 50206 42642
rect 50206 42590 50258 42642
rect 50258 42590 50260 42642
rect 50204 42588 50260 42590
rect 50204 41916 50260 41972
rect 49868 41356 49924 41412
rect 49644 40908 49700 40964
rect 49420 38722 49476 38724
rect 49420 38670 49422 38722
rect 49422 38670 49474 38722
rect 49474 38670 49476 38722
rect 49420 38668 49476 38670
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50540 41298 50596 41300
rect 50540 41246 50542 41298
rect 50542 41246 50594 41298
rect 50594 41246 50596 41298
rect 50540 41244 50596 41246
rect 50652 41186 50708 41188
rect 50652 41134 50654 41186
rect 50654 41134 50706 41186
rect 50706 41134 50708 41186
rect 50652 41132 50708 41134
rect 49084 33516 49140 33572
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 52668 47458 52724 47460
rect 52668 47406 52670 47458
rect 52670 47406 52722 47458
rect 52722 47406 52724 47458
rect 52668 47404 52724 47406
rect 53676 52108 53732 52164
rect 54124 52162 54180 52164
rect 54124 52110 54126 52162
rect 54126 52110 54178 52162
rect 54178 52110 54180 52162
rect 54124 52108 54180 52110
rect 54012 50764 54068 50820
rect 54908 55468 54964 55524
rect 55132 55468 55188 55524
rect 55020 55244 55076 55300
rect 54796 54124 54852 54180
rect 54908 54290 54964 54292
rect 54908 54238 54910 54290
rect 54910 54238 54962 54290
rect 54962 54238 54964 54290
rect 54908 54236 54964 54238
rect 55132 54572 55188 54628
rect 55132 54124 55188 54180
rect 56476 55356 56532 55412
rect 55804 53788 55860 53844
rect 56140 54348 56196 54404
rect 56812 54572 56868 54628
rect 56700 54402 56756 54404
rect 56700 54350 56702 54402
rect 56702 54350 56754 54402
rect 56754 54350 56756 54402
rect 56700 54348 56756 54350
rect 57148 54236 57204 54292
rect 56140 52386 56196 52388
rect 56140 52334 56142 52386
rect 56142 52334 56194 52386
rect 56194 52334 56196 52386
rect 56140 52332 56196 52334
rect 56588 52332 56644 52388
rect 55132 52108 55188 52164
rect 54684 51436 54740 51492
rect 54460 49756 54516 49812
rect 55468 51548 55524 51604
rect 55356 51212 55412 51268
rect 57036 51548 57092 51604
rect 56812 51436 56868 51492
rect 56476 51378 56532 51380
rect 56476 51326 56478 51378
rect 56478 51326 56530 51378
rect 56530 51326 56532 51378
rect 56476 51324 56532 51326
rect 57932 61010 57988 61012
rect 57932 60958 57934 61010
rect 57934 60958 57986 61010
rect 57986 60958 57988 61010
rect 57932 60956 57988 60958
rect 57372 59388 57428 59444
rect 57372 52834 57428 52836
rect 57372 52782 57374 52834
rect 57374 52782 57426 52834
rect 57426 52782 57428 52834
rect 57372 52780 57428 52782
rect 54908 49196 54964 49252
rect 55468 49196 55524 49252
rect 56028 49196 56084 49252
rect 54684 48636 54740 48692
rect 53900 48412 53956 48468
rect 54796 48300 54852 48356
rect 54236 48242 54292 48244
rect 54236 48190 54238 48242
rect 54238 48190 54290 48242
rect 54290 48190 54292 48242
rect 54236 48188 54292 48190
rect 55692 48636 55748 48692
rect 55468 48354 55524 48356
rect 55468 48302 55470 48354
rect 55470 48302 55522 48354
rect 55522 48302 55524 48354
rect 55468 48300 55524 48302
rect 54908 48242 54964 48244
rect 54908 48190 54910 48242
rect 54910 48190 54962 48242
rect 54962 48190 54964 48242
rect 54908 48188 54964 48190
rect 56252 48188 56308 48244
rect 53676 47404 53732 47460
rect 52108 46508 52164 46564
rect 51100 44828 51156 44884
rect 51884 44940 51940 44996
rect 51436 44828 51492 44884
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51772 43708 51828 43764
rect 51660 42588 51716 42644
rect 51660 41186 51716 41188
rect 51660 41134 51662 41186
rect 51662 41134 51714 41186
rect 51714 41134 51716 41186
rect 51660 41132 51716 41134
rect 51660 40402 51716 40404
rect 51660 40350 51662 40402
rect 51662 40350 51714 40402
rect 51714 40350 51716 40402
rect 51660 40348 51716 40350
rect 51884 41356 51940 41412
rect 51996 41244 52052 41300
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 49980 36370 50036 36372
rect 49980 36318 49982 36370
rect 49982 36318 50034 36370
rect 50034 36318 50036 36370
rect 49980 36316 50036 36318
rect 50092 35420 50148 35476
rect 49980 35026 50036 35028
rect 49980 34974 49982 35026
rect 49982 34974 50034 35026
rect 50034 34974 50036 35026
rect 49980 34972 50036 34974
rect 49420 33404 49476 33460
rect 48972 32562 49028 32564
rect 48972 32510 48974 32562
rect 48974 32510 49026 32562
rect 49026 32510 49028 32562
rect 48972 32508 49028 32510
rect 49084 32172 49140 32228
rect 49644 32562 49700 32564
rect 49644 32510 49646 32562
rect 49646 32510 49698 32562
rect 49698 32510 49700 32562
rect 49644 32508 49700 32510
rect 49532 32172 49588 32228
rect 49308 31778 49364 31780
rect 49308 31726 49310 31778
rect 49310 31726 49362 31778
rect 49362 31726 49364 31778
rect 49308 31724 49364 31726
rect 49420 31666 49476 31668
rect 49420 31614 49422 31666
rect 49422 31614 49474 31666
rect 49474 31614 49476 31666
rect 49420 31612 49476 31614
rect 48412 30604 48468 30660
rect 49084 29596 49140 29652
rect 50092 31836 50148 31892
rect 50316 36316 50372 36372
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50316 35474 50372 35476
rect 50316 35422 50318 35474
rect 50318 35422 50370 35474
rect 50370 35422 50372 35474
rect 50316 35420 50372 35422
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 52220 35644 52276 35700
rect 51772 35474 51828 35476
rect 51772 35422 51774 35474
rect 51774 35422 51826 35474
rect 51826 35422 51828 35474
rect 51772 35420 51828 35422
rect 51100 34300 51156 34356
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50428 32562 50484 32564
rect 50428 32510 50430 32562
rect 50430 32510 50482 32562
rect 50482 32510 50484 32562
rect 50428 32508 50484 32510
rect 49868 30604 49924 30660
rect 49980 30268 50036 30324
rect 51436 32060 51492 32116
rect 50876 31836 50932 31892
rect 51884 33346 51940 33348
rect 51884 33294 51886 33346
rect 51886 33294 51938 33346
rect 51938 33294 51940 33346
rect 51884 33292 51940 33294
rect 51996 33234 52052 33236
rect 51996 33182 51998 33234
rect 51998 33182 52050 33234
rect 52050 33182 52052 33234
rect 51996 33180 52052 33182
rect 52220 32620 52276 32676
rect 51772 31836 51828 31892
rect 50428 31724 50484 31780
rect 49868 30210 49924 30212
rect 49868 30158 49870 30210
rect 49870 30158 49922 30210
rect 49922 30158 49924 30210
rect 49868 30156 49924 30158
rect 50204 30882 50260 30884
rect 50204 30830 50206 30882
rect 50206 30830 50258 30882
rect 50258 30830 50260 30882
rect 50204 30828 50260 30830
rect 50764 31554 50820 31556
rect 50764 31502 50766 31554
rect 50766 31502 50818 31554
rect 50818 31502 50820 31554
rect 50764 31500 50820 31502
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50876 30828 50932 30884
rect 51548 30380 51604 30436
rect 50316 30268 50372 30324
rect 49532 28812 49588 28868
rect 48524 28754 48580 28756
rect 48524 28702 48526 28754
rect 48526 28702 48578 28754
rect 48578 28702 48580 28754
rect 48524 28700 48580 28702
rect 49756 28754 49812 28756
rect 49756 28702 49758 28754
rect 49758 28702 49810 28754
rect 49810 28702 49812 28754
rect 49756 28700 49812 28702
rect 46620 25618 46676 25620
rect 46620 25566 46622 25618
rect 46622 25566 46674 25618
rect 46674 25566 46676 25618
rect 46620 25564 46676 25566
rect 45948 25506 46004 25508
rect 45948 25454 45950 25506
rect 45950 25454 46002 25506
rect 46002 25454 46004 25506
rect 45948 25452 46004 25454
rect 47628 26066 47684 26068
rect 47628 26014 47630 26066
rect 47630 26014 47682 26066
rect 47682 26014 47684 26066
rect 47628 26012 47684 26014
rect 49084 26012 49140 26068
rect 47292 25564 47348 25620
rect 50876 30210 50932 30212
rect 50876 30158 50878 30210
rect 50878 30158 50930 30210
rect 50930 30158 50932 30210
rect 50876 30156 50932 30158
rect 54796 46562 54852 46564
rect 54796 46510 54798 46562
rect 54798 46510 54850 46562
rect 54850 46510 54852 46562
rect 54796 46508 54852 46510
rect 53004 46396 53060 46452
rect 54908 45890 54964 45892
rect 54908 45838 54910 45890
rect 54910 45838 54962 45890
rect 54962 45838 54964 45890
rect 54908 45836 54964 45838
rect 53340 45330 53396 45332
rect 53340 45278 53342 45330
rect 53342 45278 53394 45330
rect 53394 45278 53396 45330
rect 53340 45276 53396 45278
rect 54908 45276 54964 45332
rect 52892 44994 52948 44996
rect 52892 44942 52894 44994
rect 52894 44942 52946 44994
rect 52946 44942 52948 44994
rect 52892 44940 52948 44942
rect 54572 44546 54628 44548
rect 54572 44494 54574 44546
rect 54574 44494 54626 44546
rect 54626 44494 54628 44546
rect 54572 44492 54628 44494
rect 53564 43596 53620 43652
rect 52780 43538 52836 43540
rect 52780 43486 52782 43538
rect 52782 43486 52834 43538
rect 52834 43486 52836 43538
rect 52780 43484 52836 43486
rect 53228 43538 53284 43540
rect 53228 43486 53230 43538
rect 53230 43486 53282 43538
rect 53282 43486 53284 43538
rect 53228 43484 53284 43486
rect 53116 42924 53172 42980
rect 54348 44098 54404 44100
rect 54348 44046 54350 44098
rect 54350 44046 54402 44098
rect 54402 44046 54404 44098
rect 54348 44044 54404 44046
rect 55804 46508 55860 46564
rect 55020 45052 55076 45108
rect 55132 45218 55188 45220
rect 55132 45166 55134 45218
rect 55134 45166 55186 45218
rect 55186 45166 55188 45218
rect 55132 45164 55188 45166
rect 55132 44828 55188 44884
rect 54908 43708 54964 43764
rect 53900 42978 53956 42980
rect 53900 42926 53902 42978
rect 53902 42926 53954 42978
rect 53954 42926 53956 42978
rect 53900 42924 53956 42926
rect 52444 41970 52500 41972
rect 52444 41918 52446 41970
rect 52446 41918 52498 41970
rect 52498 41918 52500 41970
rect 52444 41916 52500 41918
rect 53116 41970 53172 41972
rect 53116 41918 53118 41970
rect 53118 41918 53170 41970
rect 53170 41918 53172 41970
rect 53116 41916 53172 41918
rect 53676 41916 53732 41972
rect 52892 41410 52948 41412
rect 52892 41358 52894 41410
rect 52894 41358 52946 41410
rect 52946 41358 52948 41410
rect 52892 41356 52948 41358
rect 52668 41298 52724 41300
rect 52668 41246 52670 41298
rect 52670 41246 52722 41298
rect 52722 41246 52724 41298
rect 52668 41244 52724 41246
rect 53564 40962 53620 40964
rect 53564 40910 53566 40962
rect 53566 40910 53618 40962
rect 53618 40910 53620 40962
rect 53564 40908 53620 40910
rect 53116 40348 53172 40404
rect 55244 44546 55300 44548
rect 55244 44494 55246 44546
rect 55246 44494 55298 44546
rect 55298 44494 55300 44546
rect 55244 44492 55300 44494
rect 55132 42924 55188 42980
rect 55692 45106 55748 45108
rect 55692 45054 55694 45106
rect 55694 45054 55746 45106
rect 55746 45054 55748 45106
rect 55692 45052 55748 45054
rect 55356 44268 55412 44324
rect 55468 44044 55524 44100
rect 57036 45164 57092 45220
rect 56140 44546 56196 44548
rect 56140 44494 56142 44546
rect 56142 44494 56194 44546
rect 56194 44494 56196 44546
rect 56140 44492 56196 44494
rect 57820 60674 57876 60676
rect 57820 60622 57822 60674
rect 57822 60622 57874 60674
rect 57874 60622 57876 60674
rect 57820 60620 57876 60622
rect 57708 60562 57764 60564
rect 57708 60510 57710 60562
rect 57710 60510 57762 60562
rect 57762 60510 57764 60562
rect 57708 60508 57764 60510
rect 58044 60002 58100 60004
rect 58044 59950 58046 60002
rect 58046 59950 58098 60002
rect 58098 59950 58100 60002
rect 58044 59948 58100 59950
rect 58156 59218 58212 59220
rect 58156 59166 58158 59218
rect 58158 59166 58210 59218
rect 58210 59166 58212 59218
rect 58156 59164 58212 59166
rect 57708 54572 57764 54628
rect 57596 52220 57652 52276
rect 56588 44322 56644 44324
rect 56588 44270 56590 44322
rect 56590 44270 56642 44322
rect 56642 44270 56644 44322
rect 56588 44268 56644 44270
rect 55692 43932 55748 43988
rect 54796 41916 54852 41972
rect 55356 41804 55412 41860
rect 56364 43708 56420 43764
rect 56252 41916 56308 41972
rect 54124 39058 54180 39060
rect 54124 39006 54126 39058
rect 54126 39006 54178 39058
rect 54178 39006 54180 39058
rect 54124 39004 54180 39006
rect 53676 38668 53732 38724
rect 55916 40908 55972 40964
rect 56028 40236 56084 40292
rect 56812 43708 56868 43764
rect 56700 41970 56756 41972
rect 56700 41918 56702 41970
rect 56702 41918 56754 41970
rect 56754 41918 56756 41970
rect 56700 41916 56756 41918
rect 57036 41804 57092 41860
rect 57260 41692 57316 41748
rect 57484 41858 57540 41860
rect 57484 41806 57486 41858
rect 57486 41806 57538 41858
rect 57538 41806 57540 41858
rect 57484 41804 57540 41806
rect 57596 41692 57652 41748
rect 57372 41468 57428 41524
rect 57596 41244 57652 41300
rect 56924 40908 56980 40964
rect 57484 40402 57540 40404
rect 57484 40350 57486 40402
rect 57486 40350 57538 40402
rect 57538 40350 57540 40402
rect 57484 40348 57540 40350
rect 57036 40236 57092 40292
rect 57484 40012 57540 40068
rect 56364 39004 56420 39060
rect 56812 39004 56868 39060
rect 57596 38834 57652 38836
rect 57596 38782 57598 38834
rect 57598 38782 57650 38834
rect 57650 38782 57652 38834
rect 57596 38780 57652 38782
rect 54908 38050 54964 38052
rect 54908 37998 54910 38050
rect 54910 37998 54962 38050
rect 54962 37998 54964 38050
rect 54908 37996 54964 37998
rect 55356 38050 55412 38052
rect 55356 37998 55358 38050
rect 55358 37998 55410 38050
rect 55410 37998 55412 38050
rect 55356 37996 55412 37998
rect 52892 35698 52948 35700
rect 52892 35646 52894 35698
rect 52894 35646 52946 35698
rect 52946 35646 52948 35698
rect 52892 35644 52948 35646
rect 53116 35474 53172 35476
rect 53116 35422 53118 35474
rect 53118 35422 53170 35474
rect 53170 35422 53172 35474
rect 53116 35420 53172 35422
rect 52332 31164 52388 31220
rect 52668 32620 52724 32676
rect 51772 30268 51828 30324
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 51100 29650 51156 29652
rect 51100 29598 51102 29650
rect 51102 29598 51154 29650
rect 51154 29598 51156 29650
rect 51100 29596 51156 29598
rect 50988 29426 51044 29428
rect 50988 29374 50990 29426
rect 50990 29374 51042 29426
rect 51042 29374 51044 29426
rect 50988 29372 51044 29374
rect 50652 28812 50708 28868
rect 51548 29538 51604 29540
rect 51548 29486 51550 29538
rect 51550 29486 51602 29538
rect 51602 29486 51604 29538
rect 51548 29484 51604 29486
rect 51436 28700 51492 28756
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50092 28028 50148 28084
rect 49980 25788 50036 25844
rect 50316 27804 50372 27860
rect 52780 32060 52836 32116
rect 53452 34690 53508 34692
rect 53452 34638 53454 34690
rect 53454 34638 53506 34690
rect 53506 34638 53508 34690
rect 53452 34636 53508 34638
rect 53452 33234 53508 33236
rect 53452 33182 53454 33234
rect 53454 33182 53506 33234
rect 53506 33182 53508 33234
rect 53452 33180 53508 33182
rect 53116 31500 53172 31556
rect 52668 30268 52724 30324
rect 53228 29932 53284 29988
rect 53004 29484 53060 29540
rect 53228 29372 53284 29428
rect 51660 28028 51716 28084
rect 52668 27916 52724 27972
rect 52780 28476 52836 28532
rect 51436 27858 51492 27860
rect 51436 27806 51438 27858
rect 51438 27806 51490 27858
rect 51490 27806 51492 27858
rect 51436 27804 51492 27806
rect 53004 28530 53060 28532
rect 53004 28478 53006 28530
rect 53006 28478 53058 28530
rect 53058 28478 53060 28530
rect 53004 28476 53060 28478
rect 53564 28530 53620 28532
rect 53564 28478 53566 28530
rect 53566 28478 53618 28530
rect 53618 28478 53620 28530
rect 53564 28476 53620 28478
rect 53340 27804 53396 27860
rect 55580 36316 55636 36372
rect 54012 35308 54068 35364
rect 54012 34636 54068 34692
rect 53788 33292 53844 33348
rect 55356 35698 55412 35700
rect 55356 35646 55358 35698
rect 55358 35646 55410 35698
rect 55410 35646 55412 35698
rect 55356 35644 55412 35646
rect 54012 33180 54068 33236
rect 53900 32786 53956 32788
rect 53900 32734 53902 32786
rect 53902 32734 53954 32786
rect 53954 32734 53956 32786
rect 53900 32732 53956 32734
rect 54908 32732 54964 32788
rect 55580 34076 55636 34132
rect 55020 33292 55076 33348
rect 55580 32732 55636 32788
rect 54796 32674 54852 32676
rect 54796 32622 54798 32674
rect 54798 32622 54850 32674
rect 54850 32622 54852 32674
rect 54796 32620 54852 32622
rect 55244 32060 55300 32116
rect 55132 30380 55188 30436
rect 54572 29986 54628 29988
rect 54572 29934 54574 29986
rect 54574 29934 54626 29986
rect 54626 29934 54628 29986
rect 54572 29932 54628 29934
rect 54908 29986 54964 29988
rect 54908 29934 54910 29986
rect 54910 29934 54962 29986
rect 54962 29934 54964 29986
rect 54908 29932 54964 29934
rect 53452 27692 53508 27748
rect 53004 26962 53060 26964
rect 53004 26910 53006 26962
rect 53006 26910 53058 26962
rect 53058 26910 53060 26962
rect 53004 26908 53060 26910
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 46956 25452 47012 25508
rect 45836 25340 45892 25396
rect 50204 25228 50260 25284
rect 45724 24556 45780 24612
rect 45164 23884 45220 23940
rect 45500 23996 45556 24052
rect 46060 23938 46116 23940
rect 46060 23886 46062 23938
rect 46062 23886 46114 23938
rect 46114 23886 46116 23938
rect 46060 23884 46116 23886
rect 45052 23324 45108 23380
rect 44940 23266 44996 23268
rect 44940 23214 44942 23266
rect 44942 23214 44994 23266
rect 44994 23214 44996 23266
rect 44940 23212 44996 23214
rect 45836 23324 45892 23380
rect 45612 23212 45668 23268
rect 46508 22988 46564 23044
rect 46172 22652 46228 22708
rect 45612 22370 45668 22372
rect 45612 22318 45614 22370
rect 45614 22318 45666 22370
rect 45666 22318 45668 22370
rect 45612 22316 45668 22318
rect 45388 22204 45444 22260
rect 45164 19852 45220 19908
rect 45948 22204 46004 22260
rect 52332 25564 52388 25620
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51436 23660 51492 23716
rect 46844 23324 46900 23380
rect 46732 22370 46788 22372
rect 46732 22318 46734 22370
rect 46734 22318 46786 22370
rect 46786 22318 46788 22370
rect 46732 22316 46788 22318
rect 46284 19964 46340 20020
rect 46172 19404 46228 19460
rect 44716 18956 44772 19012
rect 45276 18620 45332 18676
rect 44716 18508 44772 18564
rect 45948 18620 46004 18676
rect 44492 18450 44548 18452
rect 44492 18398 44494 18450
rect 44494 18398 44546 18450
rect 44546 18398 44548 18450
rect 44492 18396 44548 18398
rect 44940 17666 44996 17668
rect 44940 17614 44942 17666
rect 44942 17614 44994 17666
rect 44994 17614 44996 17666
rect 44940 17612 44996 17614
rect 45276 17836 45332 17892
rect 44492 17388 44548 17444
rect 43708 13634 43764 13636
rect 43708 13582 43710 13634
rect 43710 13582 43762 13634
rect 43762 13582 43764 13634
rect 43708 13580 43764 13582
rect 42924 13020 42980 13076
rect 42588 12796 42644 12852
rect 42364 12236 42420 12292
rect 41692 11900 41748 11956
rect 41020 11452 41076 11508
rect 42028 11340 42084 11396
rect 42140 12066 42196 12068
rect 42140 12014 42142 12066
rect 42142 12014 42194 12066
rect 42194 12014 42196 12066
rect 42140 12012 42196 12014
rect 41692 10834 41748 10836
rect 41692 10782 41694 10834
rect 41694 10782 41746 10834
rect 41746 10782 41748 10834
rect 41692 10780 41748 10782
rect 42140 10780 42196 10836
rect 42252 11116 42308 11172
rect 42252 10610 42308 10612
rect 42252 10558 42254 10610
rect 42254 10558 42306 10610
rect 42306 10558 42308 10610
rect 42252 10556 42308 10558
rect 40572 9212 40628 9268
rect 42588 9772 42644 9828
rect 40460 8204 40516 8260
rect 40012 8092 40068 8148
rect 41916 7980 41972 8036
rect 39900 7868 39956 7924
rect 40796 7868 40852 7924
rect 40012 7698 40068 7700
rect 40012 7646 40014 7698
rect 40014 7646 40066 7698
rect 40066 7646 40068 7698
rect 40012 7644 40068 7646
rect 40124 7586 40180 7588
rect 40124 7534 40126 7586
rect 40126 7534 40178 7586
rect 40178 7534 40180 7586
rect 40124 7532 40180 7534
rect 40684 7420 40740 7476
rect 41468 7698 41524 7700
rect 41468 7646 41470 7698
rect 41470 7646 41522 7698
rect 41522 7646 41524 7698
rect 41468 7644 41524 7646
rect 40460 6636 40516 6692
rect 41580 7532 41636 7588
rect 40236 6578 40292 6580
rect 40236 6526 40238 6578
rect 40238 6526 40290 6578
rect 40290 6526 40292 6578
rect 40236 6524 40292 6526
rect 40012 6076 40068 6132
rect 39564 5292 39620 5348
rect 40348 5234 40404 5236
rect 40348 5182 40350 5234
rect 40350 5182 40402 5234
rect 40402 5182 40404 5234
rect 40348 5180 40404 5182
rect 38220 5068 38276 5124
rect 39116 5122 39172 5124
rect 39116 5070 39118 5122
rect 39118 5070 39170 5122
rect 39170 5070 39172 5122
rect 39116 5068 39172 5070
rect 40908 5180 40964 5236
rect 40796 4396 40852 4452
rect 42140 7756 42196 7812
rect 43036 11506 43092 11508
rect 43036 11454 43038 11506
rect 43038 11454 43090 11506
rect 43090 11454 43092 11506
rect 43036 11452 43092 11454
rect 42924 10668 42980 10724
rect 43148 10610 43204 10612
rect 43148 10558 43150 10610
rect 43150 10558 43202 10610
rect 43202 10558 43204 10610
rect 43148 10556 43204 10558
rect 44044 14364 44100 14420
rect 44156 13692 44212 13748
rect 44044 12850 44100 12852
rect 44044 12798 44046 12850
rect 44046 12798 44098 12850
rect 44098 12798 44100 12850
rect 44044 12796 44100 12798
rect 43932 10722 43988 10724
rect 43932 10670 43934 10722
rect 43934 10670 43986 10722
rect 43986 10670 43988 10722
rect 43932 10668 43988 10670
rect 42924 10108 42980 10164
rect 43484 9938 43540 9940
rect 43484 9886 43486 9938
rect 43486 9886 43538 9938
rect 43538 9886 43540 9938
rect 43484 9884 43540 9886
rect 43820 9826 43876 9828
rect 43820 9774 43822 9826
rect 43822 9774 43874 9826
rect 43874 9774 43876 9826
rect 43820 9772 43876 9774
rect 42812 9266 42868 9268
rect 42812 9214 42814 9266
rect 42814 9214 42866 9266
rect 42866 9214 42868 9266
rect 42812 9212 42868 9214
rect 43484 9266 43540 9268
rect 43484 9214 43486 9266
rect 43486 9214 43538 9266
rect 43538 9214 43540 9266
rect 43484 9212 43540 9214
rect 42588 7196 42644 7252
rect 41804 6690 41860 6692
rect 41804 6638 41806 6690
rect 41806 6638 41858 6690
rect 41858 6638 41860 6690
rect 41804 6636 41860 6638
rect 43708 7644 43764 7700
rect 43260 7586 43316 7588
rect 43260 7534 43262 7586
rect 43262 7534 43314 7586
rect 43314 7534 43316 7586
rect 43260 7532 43316 7534
rect 43820 7474 43876 7476
rect 43820 7422 43822 7474
rect 43822 7422 43874 7474
rect 43874 7422 43876 7474
rect 43820 7420 43876 7422
rect 43260 6748 43316 6804
rect 45052 15820 45108 15876
rect 45388 15874 45444 15876
rect 45388 15822 45390 15874
rect 45390 15822 45442 15874
rect 45442 15822 45444 15874
rect 45388 15820 45444 15822
rect 45724 15874 45780 15876
rect 45724 15822 45726 15874
rect 45726 15822 45778 15874
rect 45778 15822 45780 15874
rect 45724 15820 45780 15822
rect 45724 15260 45780 15316
rect 44716 15202 44772 15204
rect 44716 15150 44718 15202
rect 44718 15150 44770 15202
rect 44770 15150 44772 15202
rect 44716 15148 44772 15150
rect 44716 14418 44772 14420
rect 44716 14366 44718 14418
rect 44718 14366 44770 14418
rect 44770 14366 44772 14418
rect 44716 14364 44772 14366
rect 44492 13916 44548 13972
rect 44940 13858 44996 13860
rect 44940 13806 44942 13858
rect 44942 13806 44994 13858
rect 44994 13806 44996 13858
rect 44940 13804 44996 13806
rect 45276 12850 45332 12852
rect 45276 12798 45278 12850
rect 45278 12798 45330 12850
rect 45330 12798 45332 12850
rect 45276 12796 45332 12798
rect 44716 12684 44772 12740
rect 45612 12738 45668 12740
rect 45612 12686 45614 12738
rect 45614 12686 45666 12738
rect 45666 12686 45668 12738
rect 45612 12684 45668 12686
rect 45500 12572 45556 12628
rect 44604 10668 44660 10724
rect 44380 10556 44436 10612
rect 42924 6578 42980 6580
rect 42924 6526 42926 6578
rect 42926 6526 42978 6578
rect 42978 6526 42980 6578
rect 42924 6524 42980 6526
rect 43260 6412 43316 6468
rect 43932 6412 43988 6468
rect 43820 6076 43876 6132
rect 41244 5180 41300 5236
rect 41692 4450 41748 4452
rect 41692 4398 41694 4450
rect 41694 4398 41746 4450
rect 41746 4398 41748 4450
rect 41692 4396 41748 4398
rect 44940 8258 44996 8260
rect 44940 8206 44942 8258
rect 44942 8206 44994 8258
rect 44994 8206 44996 8258
rect 44940 8204 44996 8206
rect 47964 23100 48020 23156
rect 47180 22652 47236 22708
rect 46956 21756 47012 21812
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 52444 25340 52500 25396
rect 52780 25282 52836 25284
rect 52780 25230 52782 25282
rect 52782 25230 52834 25282
rect 52834 25230 52836 25282
rect 52780 25228 52836 25230
rect 53452 26962 53508 26964
rect 53452 26910 53454 26962
rect 53454 26910 53506 26962
rect 53506 26910 53508 26962
rect 53452 26908 53508 26910
rect 53004 25506 53060 25508
rect 53004 25454 53006 25506
rect 53006 25454 53058 25506
rect 53058 25454 53060 25506
rect 53004 25452 53060 25454
rect 53676 27804 53732 27860
rect 54236 27746 54292 27748
rect 54236 27694 54238 27746
rect 54238 27694 54290 27746
rect 54290 27694 54292 27746
rect 54236 27692 54292 27694
rect 53676 26850 53732 26852
rect 53676 26798 53678 26850
rect 53678 26798 53730 26850
rect 53730 26798 53732 26850
rect 53676 26796 53732 26798
rect 53564 25564 53620 25620
rect 53452 25506 53508 25508
rect 53452 25454 53454 25506
rect 53454 25454 53506 25506
rect 53506 25454 53508 25506
rect 53452 25452 53508 25454
rect 52892 24834 52948 24836
rect 52892 24782 52894 24834
rect 52894 24782 52946 24834
rect 52946 24782 52948 24834
rect 52892 24780 52948 24782
rect 55356 30940 55412 30996
rect 55132 28476 55188 28532
rect 55356 28700 55412 28756
rect 55132 27858 55188 27860
rect 55132 27806 55134 27858
rect 55134 27806 55186 27858
rect 55186 27806 55188 27858
rect 55132 27804 55188 27806
rect 54460 27020 54516 27076
rect 55468 27970 55524 27972
rect 55468 27918 55470 27970
rect 55470 27918 55522 27970
rect 55522 27918 55524 27970
rect 55468 27916 55524 27918
rect 54236 26908 54292 26964
rect 53564 25340 53620 25396
rect 53340 24668 53396 24724
rect 52668 23772 52724 23828
rect 53004 23714 53060 23716
rect 53004 23662 53006 23714
rect 53006 23662 53058 23714
rect 53058 23662 53060 23714
rect 53004 23660 53060 23662
rect 52220 23212 52276 23268
rect 50428 23100 50484 23156
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 50764 22988 50820 23044
rect 51212 22988 51268 23044
rect 48188 22428 48244 22484
rect 50204 22428 50260 22484
rect 46844 20018 46900 20020
rect 46844 19966 46846 20018
rect 46846 19966 46898 20018
rect 46898 19966 46900 20018
rect 46844 19964 46900 19966
rect 46732 19906 46788 19908
rect 46732 19854 46734 19906
rect 46734 19854 46786 19906
rect 46786 19854 46788 19906
rect 46732 19852 46788 19854
rect 46956 19740 47012 19796
rect 46732 18508 46788 18564
rect 46620 17442 46676 17444
rect 46620 17390 46622 17442
rect 46622 17390 46674 17442
rect 46674 17390 46676 17442
rect 46620 17388 46676 17390
rect 45612 8258 45668 8260
rect 45612 8206 45614 8258
rect 45614 8206 45666 8258
rect 45666 8206 45668 8258
rect 45612 8204 45668 8206
rect 46396 8258 46452 8260
rect 46396 8206 46398 8258
rect 46398 8206 46450 8258
rect 46450 8206 46452 8258
rect 46396 8204 46452 8206
rect 45836 7756 45892 7812
rect 46172 7644 46228 7700
rect 45052 6524 45108 6580
rect 46620 15202 46676 15204
rect 46620 15150 46622 15202
rect 46622 15150 46674 15202
rect 46674 15150 46676 15202
rect 46620 15148 46676 15150
rect 47292 19964 47348 20020
rect 47180 19234 47236 19236
rect 47180 19182 47182 19234
rect 47182 19182 47234 19234
rect 47234 19182 47236 19234
rect 47180 19180 47236 19182
rect 47180 17666 47236 17668
rect 47180 17614 47182 17666
rect 47182 17614 47234 17666
rect 47234 17614 47236 17666
rect 47180 17612 47236 17614
rect 49644 21810 49700 21812
rect 49644 21758 49646 21810
rect 49646 21758 49698 21810
rect 49698 21758 49700 21810
rect 49644 21756 49700 21758
rect 49756 21698 49812 21700
rect 49756 21646 49758 21698
rect 49758 21646 49810 21698
rect 49810 21646 49812 21698
rect 49756 21644 49812 21646
rect 47516 19740 47572 19796
rect 47628 19404 47684 19460
rect 47964 19964 48020 20020
rect 47740 19292 47796 19348
rect 47852 19852 47908 19908
rect 47404 17442 47460 17444
rect 47404 17390 47406 17442
rect 47406 17390 47458 17442
rect 47458 17390 47460 17442
rect 47404 17388 47460 17390
rect 47852 15986 47908 15988
rect 47852 15934 47854 15986
rect 47854 15934 47906 15986
rect 47906 15934 47908 15986
rect 47852 15932 47908 15934
rect 47180 15820 47236 15876
rect 47740 15820 47796 15876
rect 47180 15372 47236 15428
rect 46844 15314 46900 15316
rect 46844 15262 46846 15314
rect 46846 15262 46898 15314
rect 46898 15262 46900 15314
rect 46844 15260 46900 15262
rect 47292 15484 47348 15540
rect 49980 17612 50036 17668
rect 49308 16882 49364 16884
rect 49308 16830 49310 16882
rect 49310 16830 49362 16882
rect 49362 16830 49364 16882
rect 49308 16828 49364 16830
rect 49084 16716 49140 16772
rect 48860 15372 48916 15428
rect 48972 15484 49028 15540
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50876 21644 50932 21700
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50316 19180 50372 19236
rect 50764 19292 50820 19348
rect 50316 18732 50372 18788
rect 50764 19010 50820 19012
rect 50764 18958 50766 19010
rect 50766 18958 50818 19010
rect 50818 18958 50820 19010
rect 50764 18956 50820 18958
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50428 18620 50484 18676
rect 51324 18060 51380 18116
rect 50652 17666 50708 17668
rect 50652 17614 50654 17666
rect 50654 17614 50706 17666
rect 50706 17614 50708 17666
rect 50652 17612 50708 17614
rect 51548 18396 51604 18452
rect 50876 17612 50932 17668
rect 50988 17724 51044 17780
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50316 16828 50372 16884
rect 51212 17106 51268 17108
rect 51212 17054 51214 17106
rect 51214 17054 51266 17106
rect 51266 17054 51268 17106
rect 51212 17052 51268 17054
rect 49420 15426 49476 15428
rect 49420 15374 49422 15426
rect 49422 15374 49474 15426
rect 49474 15374 49476 15426
rect 49420 15372 49476 15374
rect 47628 14364 47684 14420
rect 47404 13692 47460 13748
rect 46956 11564 47012 11620
rect 46956 10892 47012 10948
rect 46844 10108 46900 10164
rect 48076 14530 48132 14532
rect 48076 14478 48078 14530
rect 48078 14478 48130 14530
rect 48130 14478 48132 14530
rect 48076 14476 48132 14478
rect 48300 14364 48356 14420
rect 47516 13804 47572 13860
rect 47852 12850 47908 12852
rect 47852 12798 47854 12850
rect 47854 12798 47906 12850
rect 47906 12798 47908 12850
rect 47852 12796 47908 12798
rect 47516 12572 47572 12628
rect 49308 14700 49364 14756
rect 49980 15372 50036 15428
rect 50540 15986 50596 15988
rect 50540 15934 50542 15986
rect 50542 15934 50594 15986
rect 50594 15934 50596 15986
rect 50540 15932 50596 15934
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50204 15202 50260 15204
rect 50204 15150 50206 15202
rect 50206 15150 50258 15202
rect 50258 15150 50260 15202
rect 50204 15148 50260 15150
rect 50652 15036 50708 15092
rect 50540 14754 50596 14756
rect 50540 14702 50542 14754
rect 50542 14702 50594 14754
rect 50594 14702 50596 14754
rect 50540 14700 50596 14702
rect 50428 14588 50484 14644
rect 50204 14530 50260 14532
rect 50204 14478 50206 14530
rect 50206 14478 50258 14530
rect 50258 14478 50260 14530
rect 50204 14476 50260 14478
rect 51212 14812 51268 14868
rect 50764 14642 50820 14644
rect 50764 14590 50766 14642
rect 50766 14590 50818 14642
rect 50818 14590 50820 14642
rect 50764 14588 50820 14590
rect 50540 14252 50596 14308
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 51212 14530 51268 14532
rect 51212 14478 51214 14530
rect 51214 14478 51266 14530
rect 51266 14478 51268 14530
rect 51212 14476 51268 14478
rect 52220 18450 52276 18452
rect 52220 18398 52222 18450
rect 52222 18398 52274 18450
rect 52274 18398 52276 18450
rect 52220 18396 52276 18398
rect 52444 18284 52500 18340
rect 51660 17106 51716 17108
rect 51660 17054 51662 17106
rect 51662 17054 51714 17106
rect 51714 17054 51716 17106
rect 51660 17052 51716 17054
rect 52332 18226 52388 18228
rect 52332 18174 52334 18226
rect 52334 18174 52386 18226
rect 52386 18174 52388 18226
rect 52332 18172 52388 18174
rect 52108 17836 52164 17892
rect 51996 17052 52052 17108
rect 51660 16828 51716 16884
rect 52332 17836 52388 17892
rect 52220 16716 52276 16772
rect 51660 15484 51716 15540
rect 51436 15202 51492 15204
rect 51436 15150 51438 15202
rect 51438 15150 51490 15202
rect 51490 15150 51492 15202
rect 51436 15148 51492 15150
rect 51884 14812 51940 14868
rect 52108 15260 52164 15316
rect 52108 14530 52164 14532
rect 52108 14478 52110 14530
rect 52110 14478 52162 14530
rect 52162 14478 52164 14530
rect 52108 14476 52164 14478
rect 51772 14418 51828 14420
rect 51772 14366 51774 14418
rect 51774 14366 51826 14418
rect 51826 14366 51828 14418
rect 51772 14364 51828 14366
rect 50988 14252 51044 14308
rect 50204 13746 50260 13748
rect 50204 13694 50206 13746
rect 50206 13694 50258 13746
rect 50258 13694 50260 13746
rect 50204 13692 50260 13694
rect 51548 14306 51604 14308
rect 51548 14254 51550 14306
rect 51550 14254 51602 14306
rect 51602 14254 51604 14306
rect 51548 14252 51604 14254
rect 50316 13580 50372 13636
rect 49532 12460 49588 12516
rect 49756 13020 49812 13076
rect 49756 12402 49812 12404
rect 49756 12350 49758 12402
rect 49758 12350 49810 12402
rect 49810 12350 49812 12402
rect 49756 12348 49812 12350
rect 50204 12572 50260 12628
rect 48412 11564 48468 11620
rect 49868 11564 49924 11620
rect 47852 11452 47908 11508
rect 48860 11506 48916 11508
rect 48860 11454 48862 11506
rect 48862 11454 48914 11506
rect 48914 11454 48916 11506
rect 48860 11452 48916 11454
rect 49644 11452 49700 11508
rect 50092 11506 50148 11508
rect 50092 11454 50094 11506
rect 50094 11454 50146 11506
rect 50146 11454 50148 11506
rect 50092 11452 50148 11454
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50316 12236 50372 12292
rect 50652 12402 50708 12404
rect 50652 12350 50654 12402
rect 50654 12350 50706 12402
rect 50706 12350 50708 12402
rect 50652 12348 50708 12350
rect 50988 11900 51044 11956
rect 51100 11564 51156 11620
rect 51436 12348 51492 12404
rect 52444 17388 52500 17444
rect 53564 23212 53620 23268
rect 53676 23714 53732 23716
rect 53676 23662 53678 23714
rect 53678 23662 53730 23714
rect 53730 23662 53732 23714
rect 53676 23660 53732 23662
rect 58156 55298 58212 55300
rect 58156 55246 58158 55298
rect 58158 55246 58210 55298
rect 58210 55246 58212 55298
rect 58156 55244 58212 55246
rect 58156 54236 58212 54292
rect 58156 52780 58212 52836
rect 58156 52220 58212 52276
rect 58156 51548 58212 51604
rect 58156 49196 58212 49252
rect 58044 45890 58100 45892
rect 58044 45838 58046 45890
rect 58046 45838 58098 45890
rect 58098 45838 58100 45890
rect 58044 45836 58100 45838
rect 58156 45330 58212 45332
rect 58156 45278 58158 45330
rect 58158 45278 58210 45330
rect 58210 45278 58212 45330
rect 58156 45276 58212 45278
rect 58380 40012 58436 40068
rect 57708 38444 57764 38500
rect 58044 38834 58100 38836
rect 58044 38782 58046 38834
rect 58046 38782 58098 38834
rect 58098 38782 58100 38834
rect 58044 38780 58100 38782
rect 58044 38332 58100 38388
rect 58268 38444 58324 38500
rect 56700 37996 56756 38052
rect 56028 36204 56084 36260
rect 57036 36482 57092 36484
rect 57036 36430 57038 36482
rect 57038 36430 57090 36482
rect 57090 36430 57092 36482
rect 57036 36428 57092 36430
rect 56700 36370 56756 36372
rect 56700 36318 56702 36370
rect 56702 36318 56754 36370
rect 56754 36318 56756 36370
rect 56700 36316 56756 36318
rect 57148 36258 57204 36260
rect 57148 36206 57150 36258
rect 57150 36206 57202 36258
rect 57202 36206 57204 36258
rect 57148 36204 57204 36206
rect 56476 35698 56532 35700
rect 56476 35646 56478 35698
rect 56478 35646 56530 35698
rect 56530 35646 56532 35698
rect 56476 35644 56532 35646
rect 56812 35308 56868 35364
rect 56924 35644 56980 35700
rect 56924 34076 56980 34132
rect 56028 32060 56084 32116
rect 57260 34130 57316 34132
rect 57260 34078 57262 34130
rect 57262 34078 57314 34130
rect 57314 34078 57316 34130
rect 57260 34076 57316 34078
rect 57932 36428 57988 36484
rect 57820 35644 57876 35700
rect 57708 35308 57764 35364
rect 57148 33404 57204 33460
rect 57148 33234 57204 33236
rect 57148 33182 57150 33234
rect 57150 33182 57202 33234
rect 57202 33182 57204 33234
rect 57148 33180 57204 33182
rect 57036 33122 57092 33124
rect 57036 33070 57038 33122
rect 57038 33070 57090 33122
rect 57090 33070 57092 33122
rect 57036 33068 57092 33070
rect 56588 30994 56644 30996
rect 56588 30942 56590 30994
rect 56590 30942 56642 30994
rect 56642 30942 56644 30994
rect 56588 30940 56644 30942
rect 56924 30940 56980 30996
rect 57484 33346 57540 33348
rect 57484 33294 57486 33346
rect 57486 33294 57538 33346
rect 57538 33294 57540 33346
rect 57484 33292 57540 33294
rect 57596 33122 57652 33124
rect 57596 33070 57598 33122
rect 57598 33070 57650 33122
rect 57650 33070 57652 33122
rect 57596 33068 57652 33070
rect 58044 33068 58100 33124
rect 57036 29932 57092 29988
rect 56924 29650 56980 29652
rect 56924 29598 56926 29650
rect 56926 29598 56978 29650
rect 56978 29598 56980 29650
rect 56924 29596 56980 29598
rect 57372 29596 57428 29652
rect 56588 28754 56644 28756
rect 56588 28702 56590 28754
rect 56590 28702 56642 28754
rect 56642 28702 56644 28754
rect 56588 28700 56644 28702
rect 56588 28476 56644 28532
rect 57260 27970 57316 27972
rect 57260 27918 57262 27970
rect 57262 27918 57314 27970
rect 57314 27918 57316 27970
rect 57260 27916 57316 27918
rect 56924 27580 56980 27636
rect 56028 26460 56084 26516
rect 56812 27132 56868 27188
rect 57036 26514 57092 26516
rect 57036 26462 57038 26514
rect 57038 26462 57090 26514
rect 57090 26462 57092 26514
rect 57036 26460 57092 26462
rect 58156 32060 58212 32116
rect 58156 31388 58212 31444
rect 57708 29932 57764 29988
rect 58156 29596 58212 29652
rect 58044 28700 58100 28756
rect 57932 27970 57988 27972
rect 57932 27918 57934 27970
rect 57934 27918 57986 27970
rect 57986 27918 57988 27970
rect 57932 27916 57988 27918
rect 57932 27634 57988 27636
rect 57932 27582 57934 27634
rect 57934 27582 57986 27634
rect 57986 27582 57988 27634
rect 57932 27580 57988 27582
rect 57596 26124 57652 26180
rect 57484 25676 57540 25732
rect 56588 24668 56644 24724
rect 55916 24444 55972 24500
rect 57596 25282 57652 25284
rect 57596 25230 57598 25282
rect 57598 25230 57650 25282
rect 57650 25230 57652 25282
rect 57596 25228 57652 25230
rect 55132 23324 55188 23380
rect 56700 23378 56756 23380
rect 56700 23326 56702 23378
rect 56702 23326 56754 23378
rect 56754 23326 56756 23378
rect 56700 23324 56756 23326
rect 54124 23266 54180 23268
rect 54124 23214 54126 23266
rect 54126 23214 54178 23266
rect 54178 23214 54180 23266
rect 54124 23212 54180 23214
rect 53900 22988 53956 23044
rect 54684 23042 54740 23044
rect 54684 22990 54686 23042
rect 54686 22990 54738 23042
rect 54738 22990 54740 23042
rect 54684 22988 54740 22990
rect 54572 22258 54628 22260
rect 54572 22206 54574 22258
rect 54574 22206 54626 22258
rect 54626 22206 54628 22258
rect 54572 22204 54628 22206
rect 56588 23266 56644 23268
rect 56588 23214 56590 23266
rect 56590 23214 56642 23266
rect 56642 23214 56644 23266
rect 56588 23212 56644 23214
rect 57148 24722 57204 24724
rect 57148 24670 57150 24722
rect 57150 24670 57202 24722
rect 57202 24670 57204 24722
rect 57148 24668 57204 24670
rect 56812 22370 56868 22372
rect 56812 22318 56814 22370
rect 56814 22318 56866 22370
rect 56866 22318 56868 22370
rect 56812 22316 56868 22318
rect 57036 22258 57092 22260
rect 57036 22206 57038 22258
rect 57038 22206 57090 22258
rect 57090 22206 57092 22258
rect 57036 22204 57092 22206
rect 55132 21980 55188 22036
rect 56924 22092 56980 22148
rect 57484 23436 57540 23492
rect 57932 23212 57988 23268
rect 57372 22370 57428 22372
rect 57372 22318 57374 22370
rect 57374 22318 57426 22370
rect 57426 22318 57428 22370
rect 57372 22316 57428 22318
rect 58268 28476 58324 28532
rect 58156 27916 58212 27972
rect 58156 27186 58212 27188
rect 58156 27134 58158 27186
rect 58158 27134 58210 27186
rect 58210 27134 58212 27186
rect 58156 27132 58212 27134
rect 58380 26236 58436 26292
rect 58156 25228 58212 25284
rect 58156 24444 58212 24500
rect 57148 21980 57204 22036
rect 57596 22146 57652 22148
rect 57596 22094 57598 22146
rect 57598 22094 57650 22146
rect 57650 22094 57652 22146
rect 57596 22092 57652 22094
rect 54908 19180 54964 19236
rect 53788 18956 53844 19012
rect 52668 18284 52724 18340
rect 52780 17890 52836 17892
rect 52780 17838 52782 17890
rect 52782 17838 52834 17890
rect 52834 17838 52836 17890
rect 52780 17836 52836 17838
rect 52668 17052 52724 17108
rect 52780 17388 52836 17444
rect 53228 18338 53284 18340
rect 53228 18286 53230 18338
rect 53230 18286 53282 18338
rect 53282 18286 53284 18338
rect 53228 18284 53284 18286
rect 54460 18338 54516 18340
rect 54460 18286 54462 18338
rect 54462 18286 54514 18338
rect 54514 18286 54516 18338
rect 54460 18284 54516 18286
rect 53564 18172 53620 18228
rect 54572 18226 54628 18228
rect 54572 18174 54574 18226
rect 54574 18174 54626 18226
rect 54626 18174 54628 18226
rect 54572 18172 54628 18174
rect 53340 17724 53396 17780
rect 53564 17554 53620 17556
rect 53564 17502 53566 17554
rect 53566 17502 53618 17554
rect 53618 17502 53620 17554
rect 53564 17500 53620 17502
rect 53116 17442 53172 17444
rect 53116 17390 53118 17442
rect 53118 17390 53170 17442
rect 53170 17390 53172 17442
rect 53116 17388 53172 17390
rect 53340 17276 53396 17332
rect 52892 16882 52948 16884
rect 52892 16830 52894 16882
rect 52894 16830 52946 16882
rect 52946 16830 52948 16882
rect 52892 16828 52948 16830
rect 52332 15538 52388 15540
rect 52332 15486 52334 15538
rect 52334 15486 52386 15538
rect 52386 15486 52388 15538
rect 52332 15484 52388 15486
rect 52556 15148 52612 15204
rect 54124 17836 54180 17892
rect 54348 17778 54404 17780
rect 54348 17726 54350 17778
rect 54350 17726 54402 17778
rect 54402 17726 54404 17778
rect 54348 17724 54404 17726
rect 54908 17612 54964 17668
rect 53788 17388 53844 17444
rect 53788 16828 53844 16884
rect 53340 16770 53396 16772
rect 53340 16718 53342 16770
rect 53342 16718 53394 16770
rect 53394 16718 53396 16770
rect 53340 16716 53396 16718
rect 52780 14642 52836 14644
rect 52780 14590 52782 14642
rect 52782 14590 52834 14642
rect 52834 14590 52836 14642
rect 52780 14588 52836 14590
rect 51884 13692 51940 13748
rect 52668 13746 52724 13748
rect 52668 13694 52670 13746
rect 52670 13694 52722 13746
rect 52722 13694 52724 13746
rect 52668 13692 52724 13694
rect 52780 13634 52836 13636
rect 52780 13582 52782 13634
rect 52782 13582 52834 13634
rect 52834 13582 52836 13634
rect 52780 13580 52836 13582
rect 53004 14476 53060 14532
rect 53564 15036 53620 15092
rect 53564 14588 53620 14644
rect 54236 15090 54292 15092
rect 54236 15038 54238 15090
rect 54238 15038 54290 15090
rect 54290 15038 54292 15090
rect 54236 15036 54292 15038
rect 55132 17276 55188 17332
rect 55020 16828 55076 16884
rect 56476 18172 56532 18228
rect 57820 17948 57876 18004
rect 57148 17666 57204 17668
rect 57148 17614 57150 17666
rect 57150 17614 57202 17666
rect 57202 17614 57204 17666
rect 57148 17612 57204 17614
rect 58156 17554 58212 17556
rect 58156 17502 58158 17554
rect 58158 17502 58210 17554
rect 58210 17502 58212 17554
rect 58156 17500 58212 17502
rect 55244 16716 55300 16772
rect 57372 16716 57428 16772
rect 54348 14642 54404 14644
rect 54348 14590 54350 14642
rect 54350 14590 54402 14642
rect 54402 14590 54404 14642
rect 54348 14588 54404 14590
rect 56476 15036 56532 15092
rect 53340 14418 53396 14420
rect 53340 14366 53342 14418
rect 53342 14366 53394 14418
rect 53394 14366 53396 14418
rect 53340 14364 53396 14366
rect 53116 14306 53172 14308
rect 53116 14254 53118 14306
rect 53118 14254 53170 14306
rect 53170 14254 53172 14306
rect 53116 14252 53172 14254
rect 55356 13692 55412 13748
rect 55244 13634 55300 13636
rect 55244 13582 55246 13634
rect 55246 13582 55298 13634
rect 55298 13582 55300 13634
rect 55244 13580 55300 13582
rect 51324 11564 51380 11620
rect 51660 11900 51716 11956
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 49532 10332 49588 10388
rect 52220 12290 52276 12292
rect 52220 12238 52222 12290
rect 52222 12238 52274 12290
rect 52274 12238 52276 12290
rect 52220 12236 52276 12238
rect 52668 12290 52724 12292
rect 52668 12238 52670 12290
rect 52670 12238 52722 12290
rect 52722 12238 52724 12290
rect 52668 12236 52724 12238
rect 52108 11394 52164 11396
rect 52108 11342 52110 11394
rect 52110 11342 52162 11394
rect 52162 11342 52164 11394
rect 52108 11340 52164 11342
rect 51772 11228 51828 11284
rect 50652 10498 50708 10500
rect 50652 10446 50654 10498
rect 50654 10446 50706 10498
rect 50706 10446 50708 10498
rect 50652 10444 50708 10446
rect 52892 12962 52948 12964
rect 52892 12910 52894 12962
rect 52894 12910 52946 12962
rect 52946 12910 52948 12962
rect 52892 12908 52948 12910
rect 56028 13746 56084 13748
rect 56028 13694 56030 13746
rect 56030 13694 56082 13746
rect 56082 13694 56084 13746
rect 56028 13692 56084 13694
rect 56700 13692 56756 13748
rect 55356 11564 55412 11620
rect 57260 11676 57316 11732
rect 52780 11340 52836 11396
rect 55580 11452 55636 11508
rect 56028 11506 56084 11508
rect 56028 11454 56030 11506
rect 56030 11454 56082 11506
rect 56082 11454 56084 11506
rect 56028 11452 56084 11454
rect 54796 11282 54852 11284
rect 54796 11230 54798 11282
rect 54798 11230 54850 11282
rect 54850 11230 54852 11282
rect 54796 11228 54852 11230
rect 51996 10834 52052 10836
rect 51996 10782 51998 10834
rect 51998 10782 52050 10834
rect 52050 10782 52052 10834
rect 51996 10780 52052 10782
rect 50204 9996 50260 10052
rect 47292 9212 47348 9268
rect 49756 9212 49812 9268
rect 46620 7756 46676 7812
rect 47404 8316 47460 8372
rect 46396 6524 46452 6580
rect 47292 8092 47348 8148
rect 51212 9996 51268 10052
rect 51100 9714 51156 9716
rect 51100 9662 51102 9714
rect 51102 9662 51154 9714
rect 51154 9662 51156 9714
rect 51100 9660 51156 9662
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 48636 8316 48692 8372
rect 47628 8258 47684 8260
rect 47628 8206 47630 8258
rect 47630 8206 47682 8258
rect 47682 8206 47684 8258
rect 47628 8204 47684 8206
rect 47516 8092 47572 8148
rect 47964 7644 48020 7700
rect 47180 6524 47236 6580
rect 45052 5906 45108 5908
rect 45052 5854 45054 5906
rect 45054 5854 45106 5906
rect 45106 5854 45108 5906
rect 45052 5852 45108 5854
rect 44940 5628 44996 5684
rect 44604 5068 44660 5124
rect 45276 5628 45332 5684
rect 45500 5122 45556 5124
rect 45500 5070 45502 5122
rect 45502 5070 45554 5122
rect 45554 5070 45556 5122
rect 45500 5068 45556 5070
rect 46508 6018 46564 6020
rect 46508 5966 46510 6018
rect 46510 5966 46562 6018
rect 46562 5966 46564 6018
rect 46508 5964 46564 5966
rect 46732 5906 46788 5908
rect 46732 5854 46734 5906
rect 46734 5854 46786 5906
rect 46786 5854 46788 5906
rect 46732 5852 46788 5854
rect 46396 5122 46452 5124
rect 46396 5070 46398 5122
rect 46398 5070 46450 5122
rect 46450 5070 46452 5122
rect 46396 5068 46452 5070
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 47068 6018 47124 6020
rect 47068 5966 47070 6018
rect 47070 5966 47122 6018
rect 47122 5966 47124 6018
rect 47068 5964 47124 5966
rect 48412 6412 48468 6468
rect 48300 6076 48356 6132
rect 47068 5122 47124 5124
rect 47068 5070 47070 5122
rect 47070 5070 47122 5122
rect 47122 5070 47124 5122
rect 47068 5068 47124 5070
rect 46956 4508 47012 4564
rect 46956 4284 47012 4340
rect 46060 4172 46116 4228
rect 47068 4226 47124 4228
rect 47068 4174 47070 4226
rect 47070 4174 47122 4226
rect 47122 4174 47124 4226
rect 47068 4172 47124 4174
rect 49644 8316 49700 8372
rect 48972 8258 49028 8260
rect 48972 8206 48974 8258
rect 48974 8206 49026 8258
rect 49026 8206 49028 8258
rect 48972 8204 49028 8206
rect 49420 8034 49476 8036
rect 49420 7982 49422 8034
rect 49422 7982 49474 8034
rect 49474 7982 49476 8034
rect 49420 7980 49476 7982
rect 48748 7644 48804 7700
rect 49868 7474 49924 7476
rect 49868 7422 49870 7474
rect 49870 7422 49922 7474
rect 49922 7422 49924 7474
rect 49868 7420 49924 7422
rect 49756 7362 49812 7364
rect 49756 7310 49758 7362
rect 49758 7310 49810 7362
rect 49810 7310 49812 7362
rect 49756 7308 49812 7310
rect 50204 8370 50260 8372
rect 50204 8318 50206 8370
rect 50206 8318 50258 8370
rect 50258 8318 50260 8370
rect 50204 8316 50260 8318
rect 51100 8370 51156 8372
rect 51100 8318 51102 8370
rect 51102 8318 51154 8370
rect 51154 8318 51156 8370
rect 51100 8316 51156 8318
rect 50764 8258 50820 8260
rect 50764 8206 50766 8258
rect 50766 8206 50818 8258
rect 50818 8206 50820 8258
rect 50764 8204 50820 8206
rect 50428 8092 50484 8148
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 51436 9884 51492 9940
rect 52108 10108 52164 10164
rect 53228 10108 53284 10164
rect 52332 9884 52388 9940
rect 51660 9772 51716 9828
rect 52892 9826 52948 9828
rect 52892 9774 52894 9826
rect 52894 9774 52946 9826
rect 52946 9774 52948 9826
rect 52892 9772 52948 9774
rect 52556 9660 52612 9716
rect 52892 9602 52948 9604
rect 52892 9550 52894 9602
rect 52894 9550 52946 9602
rect 52946 9550 52948 9602
rect 52892 9548 52948 9550
rect 54460 9548 54516 9604
rect 58156 10610 58212 10612
rect 58156 10558 58158 10610
rect 58158 10558 58210 10610
rect 58210 10558 58212 10610
rect 58156 10556 58212 10558
rect 51996 8204 52052 8260
rect 51324 8092 51380 8148
rect 50876 7586 50932 7588
rect 50876 7534 50878 7586
rect 50878 7534 50930 7586
rect 50930 7534 50932 7586
rect 50876 7532 50932 7534
rect 50652 7474 50708 7476
rect 50652 7422 50654 7474
rect 50654 7422 50706 7474
rect 50706 7422 50708 7474
rect 50652 7420 50708 7422
rect 50092 7308 50148 7364
rect 49420 6578 49476 6580
rect 49420 6526 49422 6578
rect 49422 6526 49474 6578
rect 49474 6526 49476 6578
rect 49420 6524 49476 6526
rect 50204 6748 50260 6804
rect 50652 6748 50708 6804
rect 50428 6636 50484 6692
rect 51436 7644 51492 7700
rect 51660 7420 51716 7476
rect 51548 7362 51604 7364
rect 51548 7310 51550 7362
rect 51550 7310 51602 7362
rect 51602 7310 51604 7362
rect 51548 7308 51604 7310
rect 52444 7362 52500 7364
rect 52444 7310 52446 7362
rect 52446 7310 52498 7362
rect 52498 7310 52500 7362
rect 52444 7308 52500 7310
rect 51548 6748 51604 6804
rect 52668 6802 52724 6804
rect 52668 6750 52670 6802
rect 52670 6750 52722 6802
rect 52722 6750 52724 6802
rect 52668 6748 52724 6750
rect 52556 6636 52612 6692
rect 54796 6690 54852 6692
rect 54796 6638 54798 6690
rect 54798 6638 54850 6690
rect 54850 6638 54852 6690
rect 54796 6636 54852 6638
rect 48748 4562 48804 4564
rect 48748 4510 48750 4562
rect 48750 4510 48802 4562
rect 48802 4510 48804 4562
rect 48748 4508 48804 4510
rect 50428 6412 50484 6468
rect 50316 5122 50372 5124
rect 50316 5070 50318 5122
rect 50318 5070 50370 5122
rect 50370 5070 50372 5122
rect 50316 5068 50372 5070
rect 48524 4172 48580 4228
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51212 6412 51268 6468
rect 53340 4956 53396 5012
rect 51324 4898 51380 4900
rect 51324 4846 51326 4898
rect 51326 4846 51378 4898
rect 51378 4846 51380 4898
rect 51324 4844 51380 4846
rect 52668 4844 52724 4900
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 55468 4956 55524 5012
rect 57596 4338 57652 4340
rect 57596 4286 57598 4338
rect 57598 4286 57650 4338
rect 57650 4286 57652 4338
rect 57596 4284 57652 4286
rect 57372 4226 57428 4228
rect 57372 4174 57374 4226
rect 57374 4174 57426 4226
rect 57426 4174 57428 4226
rect 57372 4172 57428 4174
rect 58156 4172 58212 4228
rect 58156 3612 58212 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 4722 66780 4732 66836
rect 4788 66780 5516 66836
rect 5572 66780 5582 66836
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 24882 66444 24892 66500
rect 24948 66444 26124 66500
rect 26180 66444 26190 66500
rect 38994 66444 39004 66500
rect 39060 66444 40796 66500
rect 40852 66444 40862 66500
rect 45042 66444 45052 66500
rect 45108 66444 48412 66500
rect 48468 66444 48478 66500
rect 49074 66444 49084 66500
rect 49140 66444 52220 66500
rect 52276 66444 52286 66500
rect 53106 66444 53116 66500
rect 53172 66444 56028 66500
rect 56084 66444 56094 66500
rect 59200 66164 60000 66192
rect 43026 66108 43036 66164
rect 43092 66108 46172 66164
rect 46228 66108 46238 66164
rect 58146 66108 58156 66164
rect 58212 66108 60000 66164
rect 59200 66080 60000 66108
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 51090 65548 51100 65604
rect 51156 65548 51166 65604
rect 51100 65492 51156 65548
rect 20178 65436 20188 65492
rect 20244 65436 20860 65492
rect 20916 65436 20926 65492
rect 33730 65436 33740 65492
rect 33796 65436 34860 65492
rect 34916 65436 35532 65492
rect 35588 65436 35598 65492
rect 41010 65436 41020 65492
rect 41076 65436 42700 65492
rect 42756 65436 42766 65492
rect 51100 65436 52332 65492
rect 52388 65436 52398 65492
rect 57586 65436 57596 65492
rect 57652 65436 58156 65492
rect 58212 65436 58222 65492
rect 17602 65324 17612 65380
rect 17668 65324 19516 65380
rect 19572 65324 19582 65380
rect 34962 65324 34972 65380
rect 35028 65324 35644 65380
rect 35700 65324 35710 65380
rect 38546 65324 38556 65380
rect 38612 65324 41132 65380
rect 41188 65324 42028 65380
rect 42084 65324 44380 65380
rect 44436 65324 44446 65380
rect 46498 65324 46508 65380
rect 46564 65324 47740 65380
rect 47796 65324 47806 65380
rect 51762 65324 51772 65380
rect 51828 65324 54124 65380
rect 54180 65324 54190 65380
rect 54898 65324 54908 65380
rect 54964 65324 55468 65380
rect 55524 65324 55534 65380
rect 37426 65212 37436 65268
rect 37492 65212 40124 65268
rect 40180 65212 40190 65268
rect 55346 65100 55356 65156
rect 55412 65100 57148 65156
rect 57204 65100 57214 65156
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 22530 64876 22540 64932
rect 22596 64876 23548 64932
rect 23604 64876 23614 64932
rect 30258 64876 30268 64932
rect 30324 64876 55244 64932
rect 55300 64876 55310 64932
rect 10098 64764 10108 64820
rect 10164 64764 12796 64820
rect 12852 64764 12862 64820
rect 8754 64652 8764 64708
rect 8820 64652 9436 64708
rect 9492 64652 12684 64708
rect 12740 64652 13580 64708
rect 13636 64652 16828 64708
rect 16884 64652 16894 64708
rect 17938 64652 17948 64708
rect 18004 64652 20188 64708
rect 20244 64652 20254 64708
rect 27794 64652 27804 64708
rect 27860 64652 29148 64708
rect 29204 64652 29484 64708
rect 29540 64652 30380 64708
rect 30436 64652 30446 64708
rect 36642 64652 36652 64708
rect 36708 64652 37100 64708
rect 37156 64652 38556 64708
rect 38612 64652 38622 64708
rect 11330 64540 11340 64596
rect 11396 64540 12572 64596
rect 12628 64540 12638 64596
rect 30930 64540 30940 64596
rect 30996 64540 32956 64596
rect 33012 64540 33022 64596
rect 20850 64428 20860 64484
rect 20916 64428 21420 64484
rect 21476 64428 21868 64484
rect 21924 64428 23212 64484
rect 23268 64428 23996 64484
rect 24052 64428 25452 64484
rect 25508 64428 25518 64484
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 26674 64204 26684 64260
rect 26740 64204 27468 64260
rect 27524 64204 28140 64260
rect 28196 64204 28206 64260
rect 12562 64092 12572 64148
rect 12628 64092 13804 64148
rect 13860 64092 13870 64148
rect 32620 64036 32676 64540
rect 33282 64428 33292 64484
rect 33348 64428 34636 64484
rect 34692 64428 34702 64484
rect 52098 64428 52108 64484
rect 52164 64428 52780 64484
rect 52836 64428 54908 64484
rect 54964 64428 54974 64484
rect 43652 64316 47516 64372
rect 47572 64316 47582 64372
rect 43652 64148 43708 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 45602 64204 45612 64260
rect 45668 64204 46508 64260
rect 46564 64204 46574 64260
rect 46946 64204 46956 64260
rect 47012 64204 50484 64260
rect 50428 64148 50484 64204
rect 39218 64092 39228 64148
rect 39284 64092 41580 64148
rect 41636 64092 43708 64148
rect 44930 64092 44940 64148
rect 44996 64092 49588 64148
rect 50428 64092 54236 64148
rect 54292 64092 54572 64148
rect 54628 64092 54638 64148
rect 12786 63980 12796 64036
rect 12852 63980 13692 64036
rect 13748 63980 14140 64036
rect 14196 63980 14206 64036
rect 32610 63980 32620 64036
rect 32676 63980 32686 64036
rect 44818 63980 44828 64036
rect 44884 63980 46060 64036
rect 46116 63980 46126 64036
rect 49532 63924 49588 64092
rect 55234 63980 55244 64036
rect 55300 63980 55804 64036
rect 55860 63980 55870 64036
rect 5730 63868 5740 63924
rect 5796 63868 8764 63924
rect 8820 63868 8830 63924
rect 12226 63868 12236 63924
rect 12292 63868 12908 63924
rect 12964 63868 14252 63924
rect 14308 63868 14318 63924
rect 16706 63868 16716 63924
rect 16772 63868 17612 63924
rect 17668 63868 17678 63924
rect 32498 63868 32508 63924
rect 32564 63868 33180 63924
rect 33236 63868 33246 63924
rect 43362 63868 43372 63924
rect 43428 63868 43820 63924
rect 43876 63868 43886 63924
rect 45154 63868 45164 63924
rect 45220 63868 45948 63924
rect 46004 63868 46014 63924
rect 49522 63868 49532 63924
rect 49588 63868 51324 63924
rect 51380 63868 51390 63924
rect 23650 63756 23660 63812
rect 23716 63756 32396 63812
rect 32452 63756 32462 63812
rect 55122 63756 55132 63812
rect 55188 63756 56364 63812
rect 56420 63756 56430 63812
rect 26338 63644 26348 63700
rect 26404 63644 27244 63700
rect 27300 63644 28252 63700
rect 28308 63644 28318 63700
rect 55906 63644 55916 63700
rect 55972 63644 57372 63700
rect 57428 63644 57438 63700
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 47730 63420 47740 63476
rect 47796 63420 50652 63476
rect 50708 63420 55020 63476
rect 55076 63420 55086 63476
rect 21074 63308 21084 63364
rect 21140 63308 22316 63364
rect 22372 63308 22382 63364
rect 24770 63196 24780 63252
rect 24836 63196 26236 63252
rect 26292 63196 26302 63252
rect 49970 63196 49980 63252
rect 50036 63196 51100 63252
rect 51156 63196 51166 63252
rect 52994 63196 53004 63252
rect 53060 63196 53900 63252
rect 53956 63196 55244 63252
rect 55300 63196 55310 63252
rect 13122 63084 13132 63140
rect 13188 63084 15484 63140
rect 15540 63084 17276 63140
rect 17332 63084 17342 63140
rect 26674 63084 26684 63140
rect 26740 63084 27132 63140
rect 27188 63084 27198 63140
rect 30146 63084 30156 63140
rect 30212 63084 30940 63140
rect 30996 63084 31276 63140
rect 31332 63084 31342 63140
rect 43474 63084 43484 63140
rect 43540 63084 44044 63140
rect 44100 63084 44940 63140
rect 44996 63084 45006 63140
rect 46050 63084 46060 63140
rect 46116 63084 47292 63140
rect 47348 63084 47740 63140
rect 47796 63084 47806 63140
rect 49074 63084 49084 63140
rect 49140 63084 49644 63140
rect 49700 63084 50764 63140
rect 50820 63084 50830 63140
rect 6514 62972 6524 63028
rect 6580 62972 7308 63028
rect 7364 62972 7644 63028
rect 7700 62972 7710 63028
rect 16482 62972 16492 63028
rect 16548 62972 17612 63028
rect 17668 62972 17678 63028
rect 26450 62972 26460 63028
rect 26516 62972 27244 63028
rect 27300 62972 27310 63028
rect 41010 62972 41020 63028
rect 41076 62972 41804 63028
rect 41860 62972 44156 63028
rect 44212 62972 45052 63028
rect 45108 62972 45118 63028
rect 16258 62860 16268 62916
rect 16324 62860 17388 62916
rect 17444 62860 17948 62916
rect 18004 62860 18014 62916
rect 26114 62860 26124 62916
rect 26180 62860 27020 62916
rect 27076 62860 27086 62916
rect 27570 62860 27580 62916
rect 27636 62860 28476 62916
rect 28532 62860 28542 62916
rect 28914 62860 28924 62916
rect 28980 62860 29484 62916
rect 29540 62860 29550 62916
rect 31490 62860 31500 62916
rect 31556 62860 32060 62916
rect 32116 62860 32844 62916
rect 32900 62860 32910 62916
rect 41906 62860 41916 62916
rect 41972 62860 42924 62916
rect 42980 62860 42990 62916
rect 45266 62860 45276 62916
rect 45332 62860 47180 62916
rect 47236 62860 47246 62916
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 7084 62524 8540 62580
rect 8596 62524 8606 62580
rect 39442 62524 39452 62580
rect 39508 62524 48692 62580
rect 48850 62524 48860 62580
rect 48916 62524 52108 62580
rect 52164 62524 52174 62580
rect 55010 62524 55020 62580
rect 55076 62524 55580 62580
rect 55636 62524 55646 62580
rect 7084 62356 7140 62524
rect 48636 62468 48692 62524
rect 7858 62412 7868 62468
rect 7924 62412 10556 62468
rect 10612 62412 10622 62468
rect 10882 62412 10892 62468
rect 10948 62412 18956 62468
rect 19012 62412 19022 62468
rect 20402 62412 20412 62468
rect 20468 62412 20860 62468
rect 20916 62412 32060 62468
rect 32116 62412 32956 62468
rect 33012 62412 33022 62468
rect 37874 62412 37884 62468
rect 37940 62412 45276 62468
rect 45332 62412 45342 62468
rect 46050 62412 46060 62468
rect 46116 62412 46508 62468
rect 46564 62412 46574 62468
rect 48636 62412 52444 62468
rect 52500 62412 53228 62468
rect 53284 62412 53294 62468
rect 6738 62300 6748 62356
rect 6804 62300 7084 62356
rect 7140 62300 7150 62356
rect 7970 62300 7980 62356
rect 8036 62300 9548 62356
rect 9604 62300 10220 62356
rect 10276 62300 10286 62356
rect 11890 62300 11900 62356
rect 11956 62300 13580 62356
rect 13636 62300 13646 62356
rect 18162 62300 18172 62356
rect 18228 62300 19516 62356
rect 19572 62300 19582 62356
rect 36306 62300 36316 62356
rect 36372 62300 41244 62356
rect 41300 62300 41310 62356
rect 42690 62300 42700 62356
rect 42756 62300 43484 62356
rect 43540 62300 43550 62356
rect 43652 62300 43932 62356
rect 43988 62300 43998 62356
rect 44930 62300 44940 62356
rect 44996 62300 45724 62356
rect 45780 62300 45790 62356
rect 27234 62188 27244 62244
rect 27300 62188 28364 62244
rect 28420 62188 29484 62244
rect 29540 62188 29550 62244
rect 36754 62188 36764 62244
rect 36820 62188 41020 62244
rect 41076 62188 42252 62244
rect 42308 62188 42318 62244
rect 43586 62188 43596 62244
rect 43652 62188 43708 62300
rect 50082 62188 50092 62244
rect 50148 62188 51660 62244
rect 51716 62188 51726 62244
rect 52882 62188 52892 62244
rect 52948 62188 54124 62244
rect 54180 62188 54190 62244
rect 25890 62076 25900 62132
rect 25956 62076 27692 62132
rect 27748 62076 27758 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 48850 61852 48860 61908
rect 48916 61852 50988 61908
rect 51044 61852 51054 61908
rect 11778 61628 11788 61684
rect 11844 61628 12236 61684
rect 12292 61628 12684 61684
rect 12740 61628 15596 61684
rect 15652 61628 15662 61684
rect 54124 61572 54180 62188
rect 54124 61516 55468 61572
rect 55524 61516 55534 61572
rect 35634 61404 35644 61460
rect 35700 61404 37212 61460
rect 37268 61404 37278 61460
rect 42018 61404 42028 61460
rect 42084 61404 43708 61460
rect 43764 61404 44156 61460
rect 44212 61404 44222 61460
rect 6178 61292 6188 61348
rect 6244 61292 6860 61348
rect 6916 61292 6926 61348
rect 22642 61292 22652 61348
rect 22708 61292 25564 61348
rect 25620 61292 41020 61348
rect 41076 61292 41086 61348
rect 28130 61180 28140 61236
rect 28196 61180 34748 61236
rect 34804 61180 35420 61236
rect 35476 61180 36092 61236
rect 36148 61180 36158 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 29586 61068 29596 61124
rect 29652 61068 34636 61124
rect 34692 61068 35196 61124
rect 35252 61068 35868 61124
rect 35924 61068 35934 61124
rect 25442 60956 25452 61012
rect 25508 60956 26012 61012
rect 26068 60956 26078 61012
rect 38322 60956 38332 61012
rect 38388 60956 39956 61012
rect 49046 60956 49084 61012
rect 49140 60956 49150 61012
rect 49746 60956 49756 61012
rect 49812 60956 50428 61012
rect 50484 60956 50988 61012
rect 51044 60956 51436 61012
rect 51492 60956 51502 61012
rect 54450 60956 54460 61012
rect 54516 60956 55244 61012
rect 55300 60956 56700 61012
rect 56756 60956 57932 61012
rect 57988 60956 57998 61012
rect 10994 60844 11004 60900
rect 11060 60844 13244 60900
rect 13300 60844 13310 60900
rect 16258 60844 16268 60900
rect 16324 60844 17500 60900
rect 17556 60844 17566 60900
rect 27794 60844 27804 60900
rect 27860 60844 33852 60900
rect 33908 60844 34748 60900
rect 34804 60844 34814 60900
rect 35410 60844 35420 60900
rect 35476 60844 37548 60900
rect 37604 60844 37614 60900
rect 38612 60844 39116 60900
rect 39172 60844 39182 60900
rect 38612 60788 38668 60844
rect 39900 60788 39956 60956
rect 49084 60900 49140 60956
rect 49084 60844 50204 60900
rect 50260 60844 50270 60900
rect 54338 60844 54348 60900
rect 54404 60844 55804 60900
rect 55860 60844 56588 60900
rect 56644 60844 56654 60900
rect 10210 60732 10220 60788
rect 10276 60732 10780 60788
rect 10836 60732 13356 60788
rect 13412 60732 13422 60788
rect 15698 60732 15708 60788
rect 15764 60732 27748 60788
rect 27906 60732 27916 60788
rect 27972 60732 28924 60788
rect 28980 60732 28990 60788
rect 32386 60732 32396 60788
rect 32452 60732 37772 60788
rect 37828 60732 38668 60788
rect 39890 60732 39900 60788
rect 39956 60732 39966 60788
rect 40226 60732 40236 60788
rect 40292 60732 51660 60788
rect 51716 60732 53004 60788
rect 53060 60732 53070 60788
rect 27692 60676 27748 60732
rect 5618 60620 5628 60676
rect 5684 60620 6300 60676
rect 6356 60620 6366 60676
rect 21746 60620 21756 60676
rect 21812 60620 23212 60676
rect 23268 60620 23548 60676
rect 23604 60620 25676 60676
rect 25732 60620 25742 60676
rect 25890 60620 25900 60676
rect 25956 60620 27132 60676
rect 27188 60620 27198 60676
rect 27682 60620 27692 60676
rect 27748 60620 28700 60676
rect 28756 60620 28766 60676
rect 37314 60620 37324 60676
rect 37380 60620 37996 60676
rect 38052 60620 38668 60676
rect 38724 60620 39004 60676
rect 39060 60620 39070 60676
rect 49522 60620 49532 60676
rect 49588 60620 49756 60676
rect 49812 60620 49822 60676
rect 50978 60620 50988 60676
rect 51044 60620 52780 60676
rect 52836 60620 52846 60676
rect 57138 60620 57148 60676
rect 57204 60620 57820 60676
rect 57876 60620 57886 60676
rect 25900 60564 25956 60620
rect 12562 60508 12572 60564
rect 12628 60508 13804 60564
rect 13860 60508 13870 60564
rect 25442 60508 25452 60564
rect 25508 60508 25956 60564
rect 27234 60508 27244 60564
rect 27300 60508 28028 60564
rect 28084 60508 29932 60564
rect 29988 60508 29998 60564
rect 32050 60508 32060 60564
rect 32116 60508 33068 60564
rect 33124 60508 33134 60564
rect 34738 60508 34748 60564
rect 34804 60508 36988 60564
rect 37044 60508 37054 60564
rect 39890 60508 39900 60564
rect 39956 60508 41468 60564
rect 41524 60508 41916 60564
rect 41972 60508 42476 60564
rect 42532 60508 42542 60564
rect 53330 60508 53340 60564
rect 53396 60508 54684 60564
rect 54740 60508 56700 60564
rect 56756 60508 57708 60564
rect 57764 60508 57774 60564
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 18834 60284 18844 60340
rect 18900 60284 20188 60340
rect 20244 60284 20254 60340
rect 26852 60284 33180 60340
rect 33236 60284 33246 60340
rect 26852 60228 26908 60284
rect 17602 60172 17612 60228
rect 17668 60172 26908 60228
rect 28354 60172 28364 60228
rect 28420 60172 29260 60228
rect 29316 60172 29326 60228
rect 44258 60172 44268 60228
rect 44324 60172 48860 60228
rect 48916 60172 48926 60228
rect 51202 60172 51212 60228
rect 51268 60172 51884 60228
rect 51940 60172 51950 60228
rect 2818 60060 2828 60116
rect 2884 60060 5124 60116
rect 10546 60060 10556 60116
rect 10612 60060 12796 60116
rect 12852 60060 15148 60116
rect 18162 60060 18172 60116
rect 18228 60060 19852 60116
rect 19908 60060 19918 60116
rect 20132 60060 26908 60116
rect 5068 60004 5124 60060
rect 5068 59948 5908 60004
rect 9090 59948 9100 60004
rect 9156 59948 11788 60004
rect 11844 59948 11854 60004
rect 12450 59948 12460 60004
rect 12516 59948 14140 60004
rect 14196 59948 14206 60004
rect 15092 59948 15148 60060
rect 20132 60004 20188 60060
rect 15204 59948 15214 60004
rect 15586 59948 15596 60004
rect 15652 59948 20188 60004
rect 5852 59780 5908 59948
rect 26852 59892 26908 60060
rect 27458 59948 27468 60004
rect 27524 59948 29372 60004
rect 29428 59948 29438 60004
rect 30370 59948 30380 60004
rect 30436 59948 32396 60004
rect 32452 59948 32462 60004
rect 40226 59948 40236 60004
rect 40292 59948 44940 60004
rect 44996 59948 45006 60004
rect 52098 59948 52108 60004
rect 52164 59948 53340 60004
rect 53396 59948 54236 60004
rect 54292 59948 54302 60004
rect 54898 59948 54908 60004
rect 54964 59948 58044 60004
rect 58100 59948 58110 60004
rect 16146 59836 16156 59892
rect 16212 59836 18060 59892
rect 18116 59836 18126 59892
rect 23986 59836 23996 59892
rect 24052 59836 26572 59892
rect 26628 59836 26638 59892
rect 26852 59836 38164 59892
rect 38108 59780 38164 59836
rect 5842 59724 5852 59780
rect 5908 59724 8428 59780
rect 8484 59724 11340 59780
rect 11396 59724 12796 59780
rect 12852 59724 12862 59780
rect 15026 59724 15036 59780
rect 15092 59724 16940 59780
rect 16996 59724 17006 59780
rect 31154 59724 31164 59780
rect 31220 59724 33628 59780
rect 33684 59724 33694 59780
rect 38098 59724 38108 59780
rect 38164 59724 38174 59780
rect 40786 59724 40796 59780
rect 40852 59724 41468 59780
rect 41524 59724 41534 59780
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 40674 59500 40684 59556
rect 40740 59500 41244 59556
rect 41300 59500 41310 59556
rect 3490 59388 3500 59444
rect 3556 59388 7644 59444
rect 7700 59388 7710 59444
rect 16706 59388 16716 59444
rect 16772 59388 18172 59444
rect 18228 59388 18238 59444
rect 41794 59388 41804 59444
rect 41860 59388 42812 59444
rect 42868 59388 44156 59444
rect 44212 59388 44222 59444
rect 47058 59388 47068 59444
rect 47124 59388 48300 59444
rect 48356 59388 50428 59444
rect 50484 59388 51436 59444
rect 51492 59388 54684 59444
rect 54740 59388 54750 59444
rect 56690 59388 56700 59444
rect 56756 59388 57372 59444
rect 57428 59388 57438 59444
rect 7522 59276 7532 59332
rect 7588 59276 8204 59332
rect 8260 59276 16660 59332
rect 17602 59276 17612 59332
rect 17668 59276 18060 59332
rect 18116 59276 18126 59332
rect 36194 59276 36204 59332
rect 36260 59276 37212 59332
rect 37268 59276 37278 59332
rect 42354 59276 42364 59332
rect 42420 59276 43036 59332
rect 43092 59276 43102 59332
rect 48178 59276 48188 59332
rect 48244 59276 49532 59332
rect 49588 59276 49598 59332
rect 16604 59220 16660 59276
rect 59200 59220 60000 59248
rect 15922 59164 15932 59220
rect 15988 59164 16380 59220
rect 16436 59164 16446 59220
rect 16604 59164 20300 59220
rect 20356 59164 21084 59220
rect 21140 59164 21150 59220
rect 41234 59164 41244 59220
rect 41300 59164 43260 59220
rect 43316 59164 43326 59220
rect 43810 59164 43820 59220
rect 43876 59164 45276 59220
rect 45332 59164 45724 59220
rect 45780 59164 48636 59220
rect 48692 59164 55692 59220
rect 55748 59164 56812 59220
rect 56868 59164 56878 59220
rect 58146 59164 58156 59220
rect 58212 59164 60000 59220
rect 59200 59136 60000 59164
rect 12786 59052 12796 59108
rect 12852 59052 16492 59108
rect 16548 59052 16558 59108
rect 18050 59052 18060 59108
rect 18116 59052 20188 59108
rect 31602 59052 31612 59108
rect 31668 59052 32284 59108
rect 32340 59052 33404 59108
rect 33460 59052 33470 59108
rect 39218 59052 39228 59108
rect 39284 59052 41020 59108
rect 41076 59052 41086 59108
rect 20132 58996 20188 59052
rect 20132 58940 37324 58996
rect 37380 58940 37390 58996
rect 38994 58940 39004 58996
rect 39060 58940 39452 58996
rect 39508 58940 41916 58996
rect 41972 58940 41982 58996
rect 12226 58828 12236 58884
rect 12292 58828 14364 58884
rect 14420 58828 14430 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 43250 58716 43260 58772
rect 43316 58716 48860 58772
rect 48916 58716 48926 58772
rect 37762 58492 37772 58548
rect 37828 58492 38556 58548
rect 38612 58492 41020 58548
rect 41076 58492 41804 58548
rect 41860 58492 42364 58548
rect 42420 58492 42430 58548
rect 45266 58492 45276 58548
rect 45332 58492 46956 58548
rect 47012 58492 47022 58548
rect 13794 58380 13804 58436
rect 13860 58380 14924 58436
rect 14980 58380 14990 58436
rect 16370 58380 16380 58436
rect 16436 58380 16446 58436
rect 25218 58380 25228 58436
rect 25284 58380 26684 58436
rect 26740 58380 26750 58436
rect 43138 58380 43148 58436
rect 43204 58380 44828 58436
rect 44884 58380 44894 58436
rect 0 58324 800 58352
rect 16380 58324 16436 58380
rect 0 58268 1708 58324
rect 1764 58268 1774 58324
rect 10994 58268 11004 58324
rect 11060 58268 11788 58324
rect 11844 58268 11854 58324
rect 16380 58268 16604 58324
rect 16660 58268 16670 58324
rect 29810 58268 29820 58324
rect 29876 58268 30492 58324
rect 30548 58268 30558 58324
rect 41122 58268 41132 58324
rect 41188 58268 52556 58324
rect 52612 58268 53004 58324
rect 53060 58268 53070 58324
rect 0 58240 800 58268
rect 2482 58156 2492 58212
rect 2548 58156 3948 58212
rect 4004 58156 4014 58212
rect 5506 58156 5516 58212
rect 5572 58156 5740 58212
rect 5796 58156 5806 58212
rect 5058 58044 5068 58100
rect 5124 58044 5852 58100
rect 5908 58044 5918 58100
rect 30370 58044 30380 58100
rect 30436 58044 30446 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 30380 57876 30436 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 19730 57820 19740 57876
rect 19796 57820 20300 57876
rect 20356 57820 30436 57876
rect 1810 57708 1820 57764
rect 1876 57708 2828 57764
rect 2884 57708 2894 57764
rect 3826 57708 3836 57764
rect 3892 57708 4172 57764
rect 4228 57708 4956 57764
rect 5012 57708 5022 57764
rect 14914 57708 14924 57764
rect 14980 57708 15484 57764
rect 15540 57708 15550 57764
rect 20738 57708 20748 57764
rect 20804 57708 26012 57764
rect 26068 57708 26078 57764
rect 28242 57708 28252 57764
rect 28308 57708 35980 57764
rect 36036 57708 37660 57764
rect 37716 57708 37726 57764
rect 8418 57596 8428 57652
rect 8484 57596 9436 57652
rect 9492 57596 9502 57652
rect 10098 57596 10108 57652
rect 10164 57596 10668 57652
rect 10724 57596 10734 57652
rect 19394 57596 19404 57652
rect 19460 57596 20300 57652
rect 20356 57596 20366 57652
rect 20748 57540 20804 57708
rect 30146 57596 30156 57652
rect 30212 57596 30940 57652
rect 30996 57596 31006 57652
rect 43586 57596 43596 57652
rect 43652 57596 44492 57652
rect 44548 57596 44558 57652
rect 51426 57596 51436 57652
rect 51492 57596 51502 57652
rect 51436 57540 51492 57596
rect 4610 57484 4620 57540
rect 4676 57484 5628 57540
rect 5684 57484 5694 57540
rect 11890 57484 11900 57540
rect 11956 57484 12460 57540
rect 12516 57484 13356 57540
rect 13412 57484 13916 57540
rect 13972 57484 13982 57540
rect 19058 57484 19068 57540
rect 19124 57484 20804 57540
rect 32274 57484 32284 57540
rect 32340 57484 32844 57540
rect 32900 57484 33180 57540
rect 33236 57484 33740 57540
rect 33796 57484 33806 57540
rect 42578 57484 42588 57540
rect 42644 57484 43148 57540
rect 43204 57484 43214 57540
rect 51090 57484 51100 57540
rect 51156 57484 51492 57540
rect 34962 57372 34972 57428
rect 35028 57372 37772 57428
rect 37828 57372 37838 57428
rect 47058 57372 47068 57428
rect 47124 57372 48188 57428
rect 48244 57372 49420 57428
rect 49476 57372 49486 57428
rect 30034 57260 30044 57316
rect 30100 57260 30604 57316
rect 30660 57260 31612 57316
rect 31668 57260 31678 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 5842 57036 5852 57092
rect 5908 57036 6188 57092
rect 6244 57036 6254 57092
rect 9986 57036 9996 57092
rect 10052 57036 10444 57092
rect 10500 57036 10510 57092
rect 10770 57036 10780 57092
rect 10836 57036 12236 57092
rect 12292 57036 12302 57092
rect 32386 56924 32396 56980
rect 32452 56924 33740 56980
rect 33796 56924 33806 56980
rect 4050 56812 4060 56868
rect 4116 56812 4508 56868
rect 4564 56812 4844 56868
rect 4900 56812 5516 56868
rect 5572 56812 5582 56868
rect 6850 56812 6860 56868
rect 6916 56812 11284 56868
rect 19842 56812 19852 56868
rect 19908 56812 20748 56868
rect 20804 56812 20814 56868
rect 26674 56812 26684 56868
rect 26740 56812 27748 56868
rect 36418 56812 36428 56868
rect 36484 56812 37100 56868
rect 37156 56812 37166 56868
rect 37986 56812 37996 56868
rect 38052 56812 42252 56868
rect 42308 56812 42318 56868
rect 11228 56756 11284 56812
rect 5282 56700 5292 56756
rect 5348 56700 6636 56756
rect 6692 56700 9772 56756
rect 9828 56700 9838 56756
rect 11218 56700 11228 56756
rect 11284 56700 12012 56756
rect 12068 56700 12078 56756
rect 13682 56700 13692 56756
rect 13748 56700 14252 56756
rect 14308 56700 15148 56756
rect 15204 56700 15214 56756
rect 26786 56700 26796 56756
rect 26852 56700 27132 56756
rect 27188 56700 27198 56756
rect 27692 56644 27748 56812
rect 35186 56700 35196 56756
rect 35252 56700 36092 56756
rect 36148 56700 37324 56756
rect 37380 56700 38220 56756
rect 38276 56700 38286 56756
rect 42914 56700 42924 56756
rect 42980 56700 43260 56756
rect 43316 56700 43326 56756
rect 12562 56588 12572 56644
rect 12628 56588 13916 56644
rect 13972 56588 14588 56644
rect 14644 56588 14654 56644
rect 27682 56588 27692 56644
rect 27748 56588 27758 56644
rect 51986 56476 51996 56532
rect 52052 56476 52780 56532
rect 52836 56476 52846 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 8194 56252 8204 56308
rect 8260 56252 8764 56308
rect 8820 56252 9884 56308
rect 9940 56252 9950 56308
rect 12898 56252 12908 56308
rect 12964 56252 14588 56308
rect 14644 56252 14654 56308
rect 47618 56252 47628 56308
rect 47684 56252 47964 56308
rect 48020 56252 49980 56308
rect 50036 56252 50046 56308
rect 50306 56252 50316 56308
rect 50372 56252 50876 56308
rect 50932 56252 50942 56308
rect 8306 56140 8316 56196
rect 8372 56140 8988 56196
rect 9044 56140 9054 56196
rect 13346 56140 13356 56196
rect 13412 56140 14028 56196
rect 14084 56140 14094 56196
rect 22978 56140 22988 56196
rect 23044 56140 23660 56196
rect 23716 56140 24164 56196
rect 32498 56140 32508 56196
rect 32564 56140 35644 56196
rect 35700 56140 36204 56196
rect 36260 56140 36270 56196
rect 48178 56140 48188 56196
rect 48244 56140 48748 56196
rect 48804 56140 48814 56196
rect 14242 56028 14252 56084
rect 14308 56028 15148 56084
rect 15204 56028 15214 56084
rect 24108 55972 24164 56140
rect 35970 56028 35980 56084
rect 36036 56028 37212 56084
rect 37268 56028 37278 56084
rect 38612 56028 39004 56084
rect 39060 56028 39070 56084
rect 50306 56028 50316 56084
rect 50372 56028 51436 56084
rect 51492 56028 51884 56084
rect 51940 56028 51950 56084
rect 38612 55972 38668 56028
rect 24098 55916 24108 55972
rect 24164 55916 24174 55972
rect 36306 55916 36316 55972
rect 36372 55916 38668 55972
rect 41682 55916 41692 55972
rect 41748 55916 42924 55972
rect 42980 55916 42990 55972
rect 45490 55916 45500 55972
rect 45556 55916 46396 55972
rect 46452 55916 46462 55972
rect 15922 55804 15932 55860
rect 15988 55804 27020 55860
rect 27076 55804 27086 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 4844 55580 5068 55636
rect 5124 55580 6636 55636
rect 6692 55580 7196 55636
rect 7252 55580 7262 55636
rect 21298 55580 21308 55636
rect 21364 55580 25340 55636
rect 25396 55580 25406 55636
rect 4844 55524 4900 55580
rect 4386 55468 4396 55524
rect 4452 55468 4900 55524
rect 6178 55468 6188 55524
rect 6244 55468 10332 55524
rect 10388 55468 11004 55524
rect 11060 55468 11070 55524
rect 11778 55468 11788 55524
rect 11844 55468 13020 55524
rect 13076 55468 13086 55524
rect 23650 55468 23660 55524
rect 23716 55468 24444 55524
rect 24500 55468 24510 55524
rect 35186 55468 35196 55524
rect 35252 55468 35980 55524
rect 36036 55468 36046 55524
rect 53890 55468 53900 55524
rect 53956 55468 54908 55524
rect 54964 55468 54974 55524
rect 55122 55468 55132 55524
rect 55188 55468 55198 55524
rect 55132 55412 55188 55468
rect 13122 55356 13132 55412
rect 13188 55356 14028 55412
rect 14084 55356 14924 55412
rect 14980 55356 14990 55412
rect 33730 55356 33740 55412
rect 33796 55356 34860 55412
rect 34916 55356 34926 55412
rect 41570 55356 41580 55412
rect 41636 55356 42140 55412
rect 42196 55356 46732 55412
rect 46788 55356 46798 55412
rect 55132 55356 56476 55412
rect 56532 55356 56542 55412
rect 11330 55244 11340 55300
rect 11396 55244 13468 55300
rect 13524 55244 14476 55300
rect 14532 55244 14542 55300
rect 31602 55244 31612 55300
rect 31668 55244 32284 55300
rect 32340 55244 32956 55300
rect 33012 55244 33022 55300
rect 44258 55244 44268 55300
rect 44324 55244 44940 55300
rect 44996 55244 45006 55300
rect 55010 55244 55020 55300
rect 55076 55244 58156 55300
rect 58212 55244 58222 55300
rect 30706 55132 30716 55188
rect 30772 55132 31500 55188
rect 31556 55132 31566 55188
rect 38322 55132 38332 55188
rect 38388 55132 39564 55188
rect 39620 55132 39630 55188
rect 46946 55132 46956 55188
rect 47012 55132 49308 55188
rect 49364 55132 49980 55188
rect 50036 55132 50046 55188
rect 2818 55020 2828 55076
rect 2884 55020 3052 55076
rect 3108 55020 3724 55076
rect 3780 55020 3790 55076
rect 12674 55020 12684 55076
rect 12740 55020 13580 55076
rect 13636 55020 13646 55076
rect 27010 55020 27020 55076
rect 27076 55020 27916 55076
rect 27972 55020 29372 55076
rect 29428 55020 29438 55076
rect 40450 55020 40460 55076
rect 40516 55020 41468 55076
rect 41524 55020 42364 55076
rect 42420 55020 42430 55076
rect 49522 55020 49532 55076
rect 49588 55020 50428 55076
rect 50484 55020 50494 55076
rect 52882 55020 52892 55076
rect 52948 55020 53788 55076
rect 53844 55020 53854 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 41794 54684 41804 54740
rect 41860 54684 42476 54740
rect 42532 54684 42542 54740
rect 51314 54684 51324 54740
rect 51380 54684 51884 54740
rect 51940 54684 53116 54740
rect 53172 54684 53182 54740
rect 3154 54572 3164 54628
rect 3220 54572 3948 54628
rect 4004 54572 5404 54628
rect 5460 54572 5470 54628
rect 26674 54572 26684 54628
rect 26740 54572 26908 54628
rect 39442 54572 39452 54628
rect 39508 54572 40796 54628
rect 40852 54572 40862 54628
rect 46050 54572 46060 54628
rect 46116 54572 46844 54628
rect 46900 54572 49196 54628
rect 49252 54572 49262 54628
rect 55122 54572 55132 54628
rect 55188 54572 56812 54628
rect 56868 54572 57708 54628
rect 57764 54572 57774 54628
rect 26852 54516 26908 54572
rect 4610 54460 4620 54516
rect 4676 54460 5180 54516
rect 5236 54460 5246 54516
rect 12562 54460 12572 54516
rect 12628 54460 14476 54516
rect 14532 54460 15372 54516
rect 15428 54460 15438 54516
rect 15820 54460 18284 54516
rect 18340 54460 19068 54516
rect 19124 54460 19628 54516
rect 19684 54460 19694 54516
rect 26852 54460 27580 54516
rect 27636 54460 27646 54516
rect 46386 54460 46396 54516
rect 46452 54460 46956 54516
rect 47012 54460 47022 54516
rect 50306 54460 50316 54516
rect 50372 54460 50876 54516
rect 50932 54460 51660 54516
rect 51716 54460 51726 54516
rect 15820 54404 15876 54460
rect 6850 54348 6860 54404
rect 6916 54348 15876 54404
rect 16034 54348 16044 54404
rect 16100 54348 20188 54404
rect 28466 54348 28476 54404
rect 28532 54348 29148 54404
rect 29204 54348 29214 54404
rect 31042 54348 31052 54404
rect 31108 54348 31948 54404
rect 32004 54348 32014 54404
rect 46834 54348 46844 54404
rect 46900 54348 47852 54404
rect 47908 54348 47918 54404
rect 56130 54348 56140 54404
rect 56196 54348 56700 54404
rect 56756 54348 56766 54404
rect 20132 54292 20188 54348
rect 20132 54236 32508 54292
rect 32564 54236 33180 54292
rect 33236 54236 33246 54292
rect 54898 54236 54908 54292
rect 54964 54236 57148 54292
rect 57204 54236 58156 54292
rect 58212 54236 58222 54292
rect 54786 54124 54796 54180
rect 54852 54124 55132 54180
rect 55188 54124 55198 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 41010 54012 41020 54068
rect 41076 54012 42476 54068
rect 42532 54012 44268 54068
rect 44324 54012 44334 54068
rect 3378 53900 3388 53956
rect 3444 53900 4284 53956
rect 4340 53900 4350 53956
rect 23314 53900 23324 53956
rect 23380 53900 24780 53956
rect 24836 53900 29204 53956
rect 29362 53900 29372 53956
rect 29428 53900 31276 53956
rect 31332 53900 31342 53956
rect 51650 53900 51660 53956
rect 51716 53900 52668 53956
rect 52724 53900 52734 53956
rect 29148 53844 29204 53900
rect 17826 53788 17836 53844
rect 17892 53788 18732 53844
rect 18788 53788 18798 53844
rect 20514 53788 20524 53844
rect 20580 53788 20590 53844
rect 21186 53788 21196 53844
rect 21252 53788 22316 53844
rect 22372 53788 22382 53844
rect 28130 53788 28140 53844
rect 28196 53788 28924 53844
rect 28980 53788 28990 53844
rect 29148 53788 30380 53844
rect 30436 53788 31388 53844
rect 31444 53788 31454 53844
rect 36194 53788 36204 53844
rect 36260 53788 37100 53844
rect 37156 53788 37166 53844
rect 37986 53788 37996 53844
rect 38052 53788 42028 53844
rect 42084 53788 42094 53844
rect 47842 53788 47852 53844
rect 47908 53788 52780 53844
rect 52836 53788 52846 53844
rect 52994 53788 53004 53844
rect 53060 53788 55804 53844
rect 55860 53788 55870 53844
rect 20524 53732 20580 53788
rect 19842 53676 19852 53732
rect 19908 53676 20580 53732
rect 20636 53676 30716 53732
rect 30772 53676 30782 53732
rect 34514 53676 34524 53732
rect 34580 53676 36428 53732
rect 36484 53676 36494 53732
rect 39554 53676 39564 53732
rect 39620 53676 40236 53732
rect 40292 53676 40302 53732
rect 44258 53676 44268 53732
rect 44324 53676 45836 53732
rect 45892 53676 45902 53732
rect 20636 53620 20692 53676
rect 17938 53564 17948 53620
rect 18004 53564 18014 53620
rect 19394 53564 19404 53620
rect 19460 53564 20636 53620
rect 20692 53564 20702 53620
rect 23090 53564 23100 53620
rect 23156 53564 23548 53620
rect 23604 53564 24332 53620
rect 24388 53564 24398 53620
rect 39442 53564 39452 53620
rect 39508 53564 40908 53620
rect 40964 53564 45500 53620
rect 45556 53564 45566 53620
rect 17948 53508 18004 53564
rect 20076 53508 20132 53564
rect 51660 53508 51716 53788
rect 5954 53452 5964 53508
rect 6020 53452 7196 53508
rect 7252 53452 7262 53508
rect 7410 53452 7420 53508
rect 7476 53452 8092 53508
rect 8148 53452 8652 53508
rect 8708 53452 8718 53508
rect 17948 53452 18844 53508
rect 18900 53452 19628 53508
rect 19684 53452 19694 53508
rect 20066 53452 20076 53508
rect 20132 53452 20142 53508
rect 23202 53452 23212 53508
rect 23268 53452 23884 53508
rect 23940 53452 23950 53508
rect 28914 53452 28924 53508
rect 28980 53452 30044 53508
rect 30100 53452 30604 53508
rect 30660 53452 30670 53508
rect 38546 53452 38556 53508
rect 38612 53452 41020 53508
rect 41076 53452 41086 53508
rect 51650 53452 51660 53508
rect 51716 53452 51726 53508
rect 52770 53452 52780 53508
rect 52836 53452 53676 53508
rect 53732 53452 53742 53508
rect 40002 53340 40012 53396
rect 40068 53340 41356 53396
rect 41412 53340 41422 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 20626 53228 20636 53284
rect 20692 53228 21308 53284
rect 21364 53228 21374 53284
rect 47506 53228 47516 53284
rect 47572 53228 47964 53284
rect 48020 53228 48030 53284
rect 7634 53116 7644 53172
rect 7700 53116 8540 53172
rect 8596 53116 8606 53172
rect 24658 53116 24668 53172
rect 24724 53116 25340 53172
rect 25396 53116 25406 53172
rect 31266 53116 31276 53172
rect 31332 53116 32172 53172
rect 32228 53116 32238 53172
rect 35970 53116 35980 53172
rect 36036 53116 36316 53172
rect 36372 53116 37324 53172
rect 37380 53116 37390 53172
rect 46834 53116 46844 53172
rect 46900 53116 51548 53172
rect 51604 53116 51614 53172
rect 12898 53004 12908 53060
rect 12964 53004 14812 53060
rect 14868 53004 14878 53060
rect 35634 53004 35644 53060
rect 35700 53004 36652 53060
rect 36708 53004 36718 53060
rect 50978 53004 50988 53060
rect 51044 53004 51660 53060
rect 51716 53004 51726 53060
rect 17490 52892 17500 52948
rect 17556 52892 20636 52948
rect 20692 52892 20702 52948
rect 23090 52892 23100 52948
rect 23156 52892 24220 52948
rect 24276 52892 24286 52948
rect 30818 52892 30828 52948
rect 30884 52892 31276 52948
rect 31332 52892 31342 52948
rect 34402 52892 34412 52948
rect 34468 52892 35980 52948
rect 36036 52892 36764 52948
rect 36820 52892 36830 52948
rect 46386 52892 46396 52948
rect 46452 52892 46732 52948
rect 46788 52892 47516 52948
rect 47572 52892 47582 52948
rect 7298 52780 7308 52836
rect 7364 52780 8428 52836
rect 8484 52780 8494 52836
rect 10658 52780 10668 52836
rect 10724 52780 12348 52836
rect 12404 52780 12414 52836
rect 20290 52780 20300 52836
rect 20356 52780 20524 52836
rect 20580 52780 20590 52836
rect 30706 52780 30716 52836
rect 30772 52780 31948 52836
rect 32004 52780 32014 52836
rect 33282 52780 33292 52836
rect 33348 52780 33516 52836
rect 33572 52780 33582 52836
rect 43810 52780 43820 52836
rect 43876 52780 46508 52836
rect 46564 52780 46574 52836
rect 57362 52780 57372 52836
rect 57428 52780 58156 52836
rect 58212 52780 58222 52836
rect 4274 52668 4284 52724
rect 4340 52668 4956 52724
rect 5012 52668 10220 52724
rect 10276 52668 10286 52724
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 8194 52444 8204 52500
rect 8260 52444 8652 52500
rect 8708 52444 10108 52500
rect 10164 52444 11452 52500
rect 11508 52444 11518 52500
rect 47170 52444 47180 52500
rect 47236 52444 51324 52500
rect 51380 52444 51390 52500
rect 16482 52332 16492 52388
rect 16548 52332 32508 52388
rect 32564 52332 33292 52388
rect 33348 52332 33358 52388
rect 56130 52332 56140 52388
rect 56196 52332 56588 52388
rect 56644 52332 56654 52388
rect 59200 52276 60000 52304
rect 3938 52220 3948 52276
rect 4004 52220 4620 52276
rect 4676 52220 6860 52276
rect 6916 52220 6926 52276
rect 14914 52220 14924 52276
rect 14980 52220 15988 52276
rect 19170 52220 19180 52276
rect 19236 52220 20300 52276
rect 20356 52220 20366 52276
rect 20738 52220 20748 52276
rect 20804 52220 23100 52276
rect 23156 52220 23166 52276
rect 32386 52220 32396 52276
rect 32452 52220 33740 52276
rect 33796 52220 33806 52276
rect 45490 52220 45500 52276
rect 45556 52220 46732 52276
rect 46788 52220 46798 52276
rect 53330 52220 53340 52276
rect 53396 52220 57596 52276
rect 57652 52220 57662 52276
rect 58146 52220 58156 52276
rect 58212 52220 60000 52276
rect 15932 52164 15988 52220
rect 59200 52192 60000 52220
rect 10770 52108 10780 52164
rect 10836 52108 12796 52164
rect 12852 52108 13356 52164
rect 13412 52108 13692 52164
rect 13748 52108 13758 52164
rect 14466 52108 14476 52164
rect 14532 52108 15260 52164
rect 15316 52108 15326 52164
rect 15922 52108 15932 52164
rect 15988 52108 15998 52164
rect 30930 52108 30940 52164
rect 30996 52108 31836 52164
rect 31892 52108 31902 52164
rect 33394 52108 33404 52164
rect 33460 52108 35644 52164
rect 35700 52108 35710 52164
rect 53218 52108 53228 52164
rect 53284 52108 53676 52164
rect 53732 52108 54124 52164
rect 54180 52108 55132 52164
rect 55188 52108 55198 52164
rect 7970 51996 7980 52052
rect 8036 51996 8764 52052
rect 8820 51996 8830 52052
rect 40114 51996 40124 52052
rect 40180 51996 43148 52052
rect 43204 51996 44156 52052
rect 44212 51996 44222 52052
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 11778 51548 11788 51604
rect 11844 51548 13244 51604
rect 13300 51548 13468 51604
rect 13524 51548 13804 51604
rect 13860 51548 13870 51604
rect 42466 51548 42476 51604
rect 42532 51548 43260 51604
rect 43316 51548 43708 51604
rect 43764 51548 43774 51604
rect 48290 51548 48300 51604
rect 48356 51548 48748 51604
rect 48804 51548 48814 51604
rect 55458 51548 55468 51604
rect 55524 51548 57036 51604
rect 57092 51548 58156 51604
rect 58212 51548 58222 51604
rect 3378 51436 3388 51492
rect 3444 51436 5068 51492
rect 5124 51436 5134 51492
rect 22418 51436 22428 51492
rect 22484 51436 23772 51492
rect 23828 51436 23838 51492
rect 54674 51436 54684 51492
rect 54740 51436 56812 51492
rect 56868 51436 56878 51492
rect 4274 51324 4284 51380
rect 4340 51324 4396 51380
rect 4452 51324 4462 51380
rect 28466 51324 28476 51380
rect 28532 51324 29148 51380
rect 29204 51324 29214 51380
rect 43250 51324 43260 51380
rect 43316 51324 47292 51380
rect 47348 51324 47358 51380
rect 52434 51324 52444 51380
rect 52500 51324 52510 51380
rect 56466 51324 56476 51380
rect 56532 51324 56542 51380
rect 3266 51212 3276 51268
rect 3332 51212 3948 51268
rect 4004 51212 4014 51268
rect 36754 51212 36764 51268
rect 36820 51212 37772 51268
rect 37828 51212 38556 51268
rect 38612 51212 38622 51268
rect 41794 51212 41804 51268
rect 41860 51212 42252 51268
rect 42308 51212 43596 51268
rect 43652 51212 43662 51268
rect 52444 51156 52500 51324
rect 56476 51268 56532 51324
rect 55346 51212 55356 51268
rect 55412 51212 56532 51268
rect 41234 51100 41244 51156
rect 41300 51100 41692 51156
rect 41748 51100 41758 51156
rect 51090 51100 51100 51156
rect 51156 51100 51772 51156
rect 51828 51100 52500 51156
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 29026 50764 29036 50820
rect 29092 50764 32284 50820
rect 32340 50764 32350 50820
rect 41010 50764 41020 50820
rect 41076 50764 41804 50820
rect 41860 50764 41870 50820
rect 53218 50764 53228 50820
rect 53284 50764 54012 50820
rect 54068 50764 54078 50820
rect 3938 50652 3948 50708
rect 4004 50652 5516 50708
rect 5572 50652 11676 50708
rect 11732 50652 12236 50708
rect 12292 50652 12302 50708
rect 29362 50652 29372 50708
rect 29428 50652 30940 50708
rect 30996 50652 31006 50708
rect 45836 50652 51212 50708
rect 51268 50652 51278 50708
rect 45836 50596 45892 50652
rect 3602 50540 3612 50596
rect 3668 50540 5628 50596
rect 5684 50540 5694 50596
rect 28354 50540 28364 50596
rect 28420 50540 29260 50596
rect 29316 50540 29326 50596
rect 29586 50540 29596 50596
rect 29652 50540 30156 50596
rect 30212 50540 30222 50596
rect 41458 50540 41468 50596
rect 41524 50540 42812 50596
rect 42868 50540 42878 50596
rect 44146 50540 44156 50596
rect 44212 50540 44828 50596
rect 44884 50540 45836 50596
rect 45892 50540 45902 50596
rect 46050 50540 46060 50596
rect 46116 50540 46732 50596
rect 46788 50540 47628 50596
rect 47684 50540 47694 50596
rect 4162 50428 4172 50484
rect 4228 50428 5740 50484
rect 5796 50428 5806 50484
rect 26226 50428 26236 50484
rect 26292 50428 30604 50484
rect 30660 50428 30670 50484
rect 30818 50428 30828 50484
rect 30884 50428 30894 50484
rect 4246 50316 4284 50372
rect 4340 50316 4350 50372
rect 4620 50260 4676 50428
rect 30828 50372 30884 50428
rect 29922 50316 29932 50372
rect 29988 50316 30884 50372
rect 4620 50204 4732 50260
rect 4788 50204 4798 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 2482 49980 2492 50036
rect 2548 49980 4508 50036
rect 4564 49980 4574 50036
rect 10770 49980 10780 50036
rect 10836 49980 11116 50036
rect 11172 49980 12348 50036
rect 12404 49980 14028 50036
rect 14084 49980 14094 50036
rect 19506 49980 19516 50036
rect 19572 49980 26908 50036
rect 28690 49980 28700 50036
rect 28756 49980 29820 50036
rect 29876 49980 29886 50036
rect 39330 49980 39340 50036
rect 39396 49980 41020 50036
rect 41076 49980 42140 50036
rect 42196 49980 42206 50036
rect 8978 49868 8988 49924
rect 9044 49868 10220 49924
rect 10276 49868 10286 49924
rect 19282 49868 19292 49924
rect 19348 49868 20188 49924
rect 20244 49868 20254 49924
rect 26852 49812 26908 49980
rect 37650 49868 37660 49924
rect 37716 49868 38556 49924
rect 38612 49868 38622 49924
rect 39218 49868 39228 49924
rect 39284 49868 51212 49924
rect 51268 49868 51660 49924
rect 51716 49868 51726 49924
rect 8866 49756 8876 49812
rect 8932 49756 9324 49812
rect 9380 49756 10332 49812
rect 10388 49756 12684 49812
rect 12740 49756 12750 49812
rect 13234 49756 13244 49812
rect 13300 49756 14252 49812
rect 14308 49756 14318 49812
rect 19506 49756 19516 49812
rect 19572 49756 21420 49812
rect 21476 49756 21486 49812
rect 26852 49756 29036 49812
rect 29092 49756 30492 49812
rect 30548 49756 30558 49812
rect 32722 49756 32732 49812
rect 32788 49756 33404 49812
rect 33460 49756 33470 49812
rect 34178 49756 34188 49812
rect 34244 49756 35084 49812
rect 35140 49756 35150 49812
rect 41458 49756 41468 49812
rect 41524 49756 42252 49812
rect 42308 49756 42318 49812
rect 50754 49756 50764 49812
rect 50820 49756 51100 49812
rect 51156 49756 52668 49812
rect 52724 49756 54460 49812
rect 54516 49756 54526 49812
rect 19170 49644 19180 49700
rect 19236 49644 20524 49700
rect 20580 49644 31052 49700
rect 31108 49644 32508 49700
rect 32564 49644 32574 49700
rect 42130 49644 42140 49700
rect 42196 49644 43372 49700
rect 43428 49644 43438 49700
rect 14690 49532 14700 49588
rect 14756 49532 15596 49588
rect 15652 49532 15662 49588
rect 47394 49532 47404 49588
rect 47460 49532 48860 49588
rect 48916 49532 48926 49588
rect 27346 49420 27356 49476
rect 27412 49420 34860 49476
rect 34916 49420 34926 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 16258 49196 16268 49252
rect 16324 49196 32284 49252
rect 32340 49196 32956 49252
rect 33012 49196 33180 49252
rect 33236 49196 33740 49252
rect 33796 49196 33806 49252
rect 54898 49196 54908 49252
rect 54964 49196 55468 49252
rect 55524 49196 56028 49252
rect 56084 49196 58156 49252
rect 58212 49196 58222 49252
rect 8530 49084 8540 49140
rect 8596 49084 9100 49140
rect 9156 49084 9166 49140
rect 17378 49084 17388 49140
rect 17444 49084 20076 49140
rect 20132 49084 20142 49140
rect 23538 49084 23548 49140
rect 23604 49084 24444 49140
rect 24500 49084 25788 49140
rect 25844 49084 25854 49140
rect 5394 48972 5404 49028
rect 5460 48972 6076 49028
rect 6132 48972 10108 49028
rect 10164 48972 10174 49028
rect 16706 48972 16716 49028
rect 16772 48972 19068 49028
rect 19124 48972 22540 49028
rect 22596 48972 22988 49028
rect 23044 48972 25116 49028
rect 25172 48972 25182 49028
rect 30930 48972 30940 49028
rect 30996 48972 31724 49028
rect 31780 48972 31790 49028
rect 50866 48972 50876 49028
rect 50932 48972 51548 49028
rect 51604 48972 51614 49028
rect 6738 48860 6748 48916
rect 6804 48860 9324 48916
rect 9380 48860 9390 48916
rect 19954 48860 19964 48916
rect 20020 48860 20188 48916
rect 20514 48860 20524 48916
rect 20580 48860 21420 48916
rect 21476 48860 21486 48916
rect 20132 48804 20188 48860
rect 8418 48748 8428 48804
rect 8484 48748 9660 48804
rect 9716 48748 9726 48804
rect 20132 48748 20412 48804
rect 20468 48748 21308 48804
rect 21364 48748 21374 48804
rect 30482 48748 30492 48804
rect 30548 48748 35084 48804
rect 35140 48748 35150 48804
rect 20290 48636 20300 48692
rect 20356 48636 21532 48692
rect 21588 48636 21598 48692
rect 54674 48636 54684 48692
rect 54740 48636 55692 48692
rect 55748 48636 55758 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 8306 48412 8316 48468
rect 8372 48412 9548 48468
rect 9604 48412 9614 48468
rect 20962 48412 20972 48468
rect 21028 48412 21980 48468
rect 22036 48412 23324 48468
rect 23380 48412 23390 48468
rect 53890 48412 53900 48468
rect 53956 48412 53966 48468
rect 53900 48356 53956 48412
rect 8082 48300 8092 48356
rect 8148 48300 9212 48356
rect 9268 48300 9278 48356
rect 10546 48300 10556 48356
rect 10612 48300 11340 48356
rect 11396 48300 11406 48356
rect 42354 48300 42364 48356
rect 42420 48300 43372 48356
rect 43428 48300 43438 48356
rect 49186 48300 49196 48356
rect 49252 48300 53956 48356
rect 54786 48300 54796 48356
rect 54852 48300 55468 48356
rect 55524 48300 55534 48356
rect 14018 48188 14028 48244
rect 14084 48188 15484 48244
rect 15540 48188 15932 48244
rect 15988 48188 15998 48244
rect 26114 48188 26124 48244
rect 26180 48188 27468 48244
rect 27524 48188 27534 48244
rect 43026 48188 43036 48244
rect 43092 48188 43484 48244
rect 43540 48188 43550 48244
rect 54226 48188 54236 48244
rect 54292 48188 54908 48244
rect 54964 48188 56252 48244
rect 56308 48188 56318 48244
rect 4946 48076 4956 48132
rect 5012 48076 5628 48132
rect 5684 48076 5694 48132
rect 11106 48076 11116 48132
rect 11172 48076 12908 48132
rect 12964 48076 13804 48132
rect 13860 48076 14140 48132
rect 14196 48076 14206 48132
rect 23874 48076 23884 48132
rect 23940 48076 24668 48132
rect 24724 48076 24892 48132
rect 24948 48076 24958 48132
rect 41570 48076 41580 48132
rect 41636 48076 42588 48132
rect 42644 48076 42654 48132
rect 43586 47964 43596 48020
rect 43652 47964 49644 48020
rect 49700 47964 49710 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 26898 47740 26908 47796
rect 26964 47740 27244 47796
rect 27300 47740 27310 47796
rect 9538 47628 9548 47684
rect 9604 47628 11116 47684
rect 11172 47628 11182 47684
rect 21522 47628 21532 47684
rect 21588 47628 22652 47684
rect 22708 47628 22718 47684
rect 35410 47628 35420 47684
rect 35476 47628 36652 47684
rect 36708 47628 37436 47684
rect 37492 47628 37502 47684
rect 1810 47516 1820 47572
rect 1876 47516 5068 47572
rect 5124 47516 5134 47572
rect 23090 47516 23100 47572
rect 23156 47516 24332 47572
rect 24388 47516 24398 47572
rect 37986 47516 37996 47572
rect 38052 47516 41692 47572
rect 41748 47516 41758 47572
rect 42130 47516 42140 47572
rect 42196 47516 42924 47572
rect 42980 47516 43596 47572
rect 43652 47516 44268 47572
rect 44324 47516 44828 47572
rect 44884 47516 44894 47572
rect 9650 47404 9660 47460
rect 9716 47404 11116 47460
rect 11172 47404 11788 47460
rect 11844 47404 11854 47460
rect 14914 47404 14924 47460
rect 14980 47404 15372 47460
rect 15428 47404 15438 47460
rect 23650 47404 23660 47460
rect 23716 47404 24556 47460
rect 24612 47404 24622 47460
rect 27906 47404 27916 47460
rect 27972 47404 34636 47460
rect 34692 47404 34972 47460
rect 35028 47404 35038 47460
rect 36418 47404 36428 47460
rect 36484 47404 38444 47460
rect 38500 47404 38510 47460
rect 49858 47404 49868 47460
rect 49924 47404 52668 47460
rect 52724 47404 53676 47460
rect 53732 47404 53742 47460
rect 4610 47292 4620 47348
rect 4676 47292 5292 47348
rect 5348 47292 5740 47348
rect 5796 47292 5806 47348
rect 15026 47292 15036 47348
rect 15092 47292 15708 47348
rect 15764 47292 17836 47348
rect 17892 47292 17902 47348
rect 18274 47292 18284 47348
rect 18340 47292 23716 47348
rect 11778 47180 11788 47236
rect 11844 47180 12684 47236
rect 12740 47180 13020 47236
rect 13076 47180 15148 47236
rect 15092 47124 15148 47180
rect 20188 47180 21084 47236
rect 21140 47180 21150 47236
rect 15092 47068 19684 47124
rect 5394 46956 5404 47012
rect 5460 46956 6188 47012
rect 6244 46956 13692 47012
rect 13748 46956 13758 47012
rect 19628 46900 19684 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 20188 46900 20244 47180
rect 23660 47124 23716 47292
rect 26852 47292 27244 47348
rect 27300 47292 28252 47348
rect 28308 47292 28318 47348
rect 24322 47180 24332 47236
rect 24388 47180 24668 47236
rect 24724 47180 25452 47236
rect 25508 47180 25518 47236
rect 26852 47124 26908 47292
rect 37090 47180 37100 47236
rect 37156 47180 37660 47236
rect 37716 47180 38556 47236
rect 38612 47180 38622 47236
rect 43474 47180 43484 47236
rect 43540 47180 44828 47236
rect 44884 47180 47740 47236
rect 47796 47180 47806 47236
rect 48850 47180 48860 47236
rect 48916 47180 49756 47236
rect 49812 47180 49980 47236
rect 50036 47180 50046 47236
rect 23650 47068 23660 47124
rect 23716 47068 23726 47124
rect 24882 47068 24892 47124
rect 24948 47068 26908 47124
rect 28354 47068 28364 47124
rect 28420 47068 28588 47124
rect 28644 47068 29372 47124
rect 29428 47068 29438 47124
rect 36082 47068 36092 47124
rect 36148 47068 39004 47124
rect 39060 47068 39070 47124
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 25442 46956 25452 47012
rect 25508 46956 43708 47012
rect 43922 46956 43932 47012
rect 43988 46956 45276 47012
rect 45332 46956 45948 47012
rect 46004 46956 46014 47012
rect 43652 46900 43708 46956
rect 12338 46844 12348 46900
rect 12404 46844 13356 46900
rect 13412 46844 14812 46900
rect 14868 46844 18508 46900
rect 18564 46844 18574 46900
rect 19628 46844 20188 46900
rect 20244 46844 20282 46900
rect 24546 46844 24556 46900
rect 24612 46844 34748 46900
rect 34804 46844 34814 46900
rect 43652 46844 48804 46900
rect 48748 46788 48804 46844
rect 10546 46732 10556 46788
rect 10612 46732 12796 46788
rect 12852 46732 12862 46788
rect 28690 46732 28700 46788
rect 28756 46732 29820 46788
rect 29876 46732 29886 46788
rect 31462 46732 31500 46788
rect 31556 46732 31566 46788
rect 39890 46732 39900 46788
rect 39956 46732 43260 46788
rect 43316 46732 43708 46788
rect 48738 46732 48748 46788
rect 48804 46732 48814 46788
rect 43652 46676 43708 46732
rect 14242 46620 14252 46676
rect 14308 46620 14700 46676
rect 14756 46620 14766 46676
rect 19394 46620 19404 46676
rect 19460 46620 23548 46676
rect 23604 46620 25228 46676
rect 25284 46620 25294 46676
rect 35858 46620 35868 46676
rect 35924 46620 36652 46676
rect 36708 46620 37436 46676
rect 37492 46620 37502 46676
rect 37650 46620 37660 46676
rect 37716 46620 38892 46676
rect 38948 46620 38958 46676
rect 43652 46620 44492 46676
rect 44548 46620 44558 46676
rect 45378 46620 45388 46676
rect 45444 46620 45724 46676
rect 45780 46620 45790 46676
rect 49298 46620 49308 46676
rect 49364 46620 49756 46676
rect 49812 46620 50540 46676
rect 50596 46620 50606 46676
rect 2706 46508 2716 46564
rect 2772 46508 3388 46564
rect 3444 46508 3454 46564
rect 14466 46508 14476 46564
rect 14532 46508 14924 46564
rect 14980 46508 14990 46564
rect 15362 46508 15372 46564
rect 15428 46508 26012 46564
rect 26068 46508 26078 46564
rect 26226 46508 26236 46564
rect 26292 46508 27356 46564
rect 27412 46508 27422 46564
rect 31378 46508 31388 46564
rect 31444 46508 31724 46564
rect 31780 46508 31790 46564
rect 31938 46508 31948 46564
rect 32004 46508 32508 46564
rect 32564 46508 32844 46564
rect 32900 46508 37548 46564
rect 37604 46508 37614 46564
rect 41010 46508 41020 46564
rect 41076 46508 41692 46564
rect 41748 46508 41758 46564
rect 45042 46508 45052 46564
rect 45108 46508 45836 46564
rect 45892 46508 45902 46564
rect 50306 46508 50316 46564
rect 50372 46508 52108 46564
rect 52164 46508 52174 46564
rect 54786 46508 54796 46564
rect 54852 46508 55804 46564
rect 55860 46508 55870 46564
rect 19730 46396 19740 46452
rect 19796 46396 20188 46452
rect 20132 46340 20188 46396
rect 26852 46396 35756 46452
rect 35812 46396 36316 46452
rect 36372 46396 37100 46452
rect 37156 46396 37166 46452
rect 39554 46396 39564 46452
rect 39620 46396 40908 46452
rect 40964 46396 40974 46452
rect 43652 46396 47628 46452
rect 47684 46396 53004 46452
rect 53060 46396 53070 46452
rect 26852 46340 26908 46396
rect 43652 46340 43708 46396
rect 20132 46284 26908 46340
rect 38210 46284 38220 46340
rect 38276 46284 43708 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 30146 46172 30156 46228
rect 30212 46172 31052 46228
rect 31108 46172 31948 46228
rect 32004 46172 32014 46228
rect 22978 46060 22988 46116
rect 23044 46060 23660 46116
rect 23716 46060 23726 46116
rect 9986 45948 9996 46004
rect 10052 45948 10556 46004
rect 10612 45948 10622 46004
rect 13570 45948 13580 46004
rect 13636 45948 19068 46004
rect 19124 45948 19134 46004
rect 27458 45948 27468 46004
rect 27524 45948 27534 46004
rect 29810 45948 29820 46004
rect 29876 45948 31052 46004
rect 31108 45948 31118 46004
rect 27468 45892 27524 45948
rect 15810 45836 15820 45892
rect 15876 45836 17052 45892
rect 17108 45836 17118 45892
rect 27010 45836 27020 45892
rect 27076 45836 27244 45892
rect 27300 45836 27524 45892
rect 37202 45836 37212 45892
rect 37268 45836 37548 45892
rect 37604 45836 37614 45892
rect 48402 45836 48412 45892
rect 48468 45836 49532 45892
rect 49588 45836 49598 45892
rect 54898 45836 54908 45892
rect 54964 45836 58044 45892
rect 58100 45836 58110 45892
rect 8754 45724 8764 45780
rect 8820 45724 9996 45780
rect 10052 45724 14812 45780
rect 14868 45724 15484 45780
rect 15540 45724 15550 45780
rect 16258 45724 16268 45780
rect 16324 45724 17724 45780
rect 17780 45724 17790 45780
rect 18386 45724 18396 45780
rect 18452 45724 26236 45780
rect 26292 45724 26302 45780
rect 32050 45724 32060 45780
rect 32116 45724 33180 45780
rect 33236 45724 33246 45780
rect 49298 45724 49308 45780
rect 49364 45724 49980 45780
rect 50036 45724 50046 45780
rect 20738 45612 20748 45668
rect 20804 45612 21420 45668
rect 21476 45612 37996 45668
rect 38052 45612 38444 45668
rect 38500 45612 48076 45668
rect 48132 45612 48142 45668
rect 14018 45500 14028 45556
rect 14084 45500 14812 45556
rect 14868 45500 14878 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 9426 45388 9436 45444
rect 9492 45388 12796 45444
rect 12852 45388 13580 45444
rect 13636 45388 13646 45444
rect 59200 45332 60000 45360
rect 8866 45276 8876 45332
rect 8932 45276 9772 45332
rect 9828 45276 9838 45332
rect 11666 45276 11676 45332
rect 11732 45276 16828 45332
rect 16884 45276 16894 45332
rect 22306 45276 22316 45332
rect 22372 45276 23212 45332
rect 23268 45276 23278 45332
rect 34402 45276 34412 45332
rect 34468 45276 36204 45332
rect 36260 45276 36652 45332
rect 36708 45276 38892 45332
rect 38948 45276 38958 45332
rect 48290 45276 48300 45332
rect 48356 45276 48748 45332
rect 48804 45276 48814 45332
rect 53330 45276 53340 45332
rect 53396 45276 54908 45332
rect 54964 45276 54974 45332
rect 58146 45276 58156 45332
rect 58212 45276 60000 45332
rect 7522 45164 7532 45220
rect 7588 45164 8204 45220
rect 8260 45164 10108 45220
rect 10164 45164 10174 45220
rect 21634 45164 21644 45220
rect 21700 45164 22204 45220
rect 22260 45164 22270 45220
rect 31490 45164 31500 45220
rect 31556 45164 34076 45220
rect 34132 45164 34142 45220
rect 49074 45164 49084 45220
rect 49140 45164 50428 45220
rect 50484 45164 50988 45220
rect 51044 45164 51054 45220
rect 53340 45108 53396 45276
rect 59200 45248 60000 45276
rect 55122 45164 55132 45220
rect 55188 45164 57036 45220
rect 57092 45164 57102 45220
rect 6066 45052 6076 45108
rect 6132 45052 9436 45108
rect 9492 45052 9502 45108
rect 15138 45052 15148 45108
rect 15204 45052 15820 45108
rect 15876 45052 15886 45108
rect 21746 45052 21756 45108
rect 21812 45052 22428 45108
rect 22484 45052 22494 45108
rect 27906 45052 27916 45108
rect 27972 45052 28476 45108
rect 28532 45052 29148 45108
rect 29204 45052 29214 45108
rect 49970 45052 49980 45108
rect 50036 45052 53396 45108
rect 55010 45052 55020 45108
rect 55076 45052 55692 45108
rect 55748 45052 55758 45108
rect 22306 44940 22316 44996
rect 22372 44940 23100 44996
rect 23156 44940 23166 44996
rect 24658 44940 24668 44996
rect 24724 44940 25564 44996
rect 25620 44940 25630 44996
rect 32386 44940 32396 44996
rect 32452 44940 33292 44996
rect 33348 44940 33358 44996
rect 33954 44940 33964 44996
rect 34020 44940 35420 44996
rect 35476 44940 35486 44996
rect 51874 44940 51884 44996
rect 51940 44940 52892 44996
rect 52948 44940 52958 44996
rect 51090 44828 51100 44884
rect 51156 44828 51436 44884
rect 51492 44828 55132 44884
rect 55188 44828 55198 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 5170 44492 5180 44548
rect 5236 44492 6020 44548
rect 54562 44492 54572 44548
rect 54628 44492 55244 44548
rect 55300 44492 56140 44548
rect 56196 44492 56206 44548
rect 5964 44436 6020 44492
rect 3378 44380 3388 44436
rect 3444 44380 4508 44436
rect 4564 44380 5628 44436
rect 5684 44380 5694 44436
rect 5954 44380 5964 44436
rect 6020 44380 15596 44436
rect 15652 44380 15662 44436
rect 23426 44380 23436 44436
rect 23492 44380 24108 44436
rect 24164 44380 24174 44436
rect 25554 44380 25564 44436
rect 25620 44380 31388 44436
rect 31444 44380 32060 44436
rect 32116 44380 32284 44436
rect 32340 44380 32350 44436
rect 13468 44324 13524 44380
rect 4834 44268 4844 44324
rect 4900 44268 6188 44324
rect 6244 44268 6254 44324
rect 13458 44268 13468 44324
rect 13524 44268 13534 44324
rect 15092 44268 15484 44324
rect 15540 44268 15550 44324
rect 15810 44268 15820 44324
rect 15876 44268 16156 44324
rect 16212 44268 17500 44324
rect 17556 44268 17566 44324
rect 18498 44268 18508 44324
rect 18564 44268 20972 44324
rect 21028 44268 21038 44324
rect 21634 44268 21644 44324
rect 21700 44268 22092 44324
rect 22148 44268 24444 44324
rect 24500 44268 24510 44324
rect 24770 44268 24780 44324
rect 24836 44268 25340 44324
rect 25396 44268 25406 44324
rect 31154 44268 31164 44324
rect 31220 44268 31948 44324
rect 32004 44268 32396 44324
rect 32452 44268 32462 44324
rect 33058 44268 33068 44324
rect 33124 44268 33740 44324
rect 33796 44268 33806 44324
rect 38882 44268 38892 44324
rect 38948 44268 40796 44324
rect 40852 44268 42140 44324
rect 42196 44268 42206 44324
rect 55346 44268 55356 44324
rect 55412 44268 56588 44324
rect 56644 44268 56654 44324
rect 15092 44100 15148 44268
rect 12562 44044 12572 44100
rect 12628 44044 13804 44100
rect 13860 44044 15148 44100
rect 33740 44100 33796 44268
rect 34066 44156 34076 44212
rect 34132 44156 34916 44212
rect 34860 44100 34916 44156
rect 33740 44044 34636 44100
rect 34692 44044 34702 44100
rect 34850 44044 34860 44100
rect 34916 44044 43708 44100
rect 54338 44044 54348 44100
rect 54404 44044 55468 44100
rect 55524 44044 55534 44100
rect 43652 43988 43708 44044
rect 12114 43932 12124 43988
rect 12180 43932 12684 43988
rect 12740 43932 12750 43988
rect 22530 43932 22540 43988
rect 22596 43932 22876 43988
rect 22932 43932 23212 43988
rect 23268 43932 23660 43988
rect 23716 43932 36764 43988
rect 36820 43932 36830 43988
rect 43652 43932 44268 43988
rect 44324 43932 44334 43988
rect 55682 43932 55692 43988
rect 55748 43932 55758 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 35634 43820 35644 43876
rect 35700 43820 38220 43876
rect 38276 43820 38286 43876
rect 55692 43764 55748 43932
rect 2370 43708 2380 43764
rect 2436 43708 2604 43764
rect 2660 43708 2670 43764
rect 51762 43708 51772 43764
rect 51828 43708 54908 43764
rect 54964 43708 54974 43764
rect 55692 43708 56364 43764
rect 56420 43708 56812 43764
rect 56868 43708 56878 43764
rect 53564 43652 53620 43708
rect 3332 43596 5516 43652
rect 5572 43596 5582 43652
rect 16370 43596 16380 43652
rect 16436 43596 20524 43652
rect 20580 43596 20590 43652
rect 29810 43596 29820 43652
rect 29876 43596 30940 43652
rect 30996 43596 31006 43652
rect 40114 43596 40124 43652
rect 40180 43596 44156 43652
rect 44212 43596 44222 43652
rect 53554 43596 53564 43652
rect 53620 43596 53630 43652
rect 3332 43540 3388 43596
rect 1810 43484 1820 43540
rect 1876 43484 3388 43540
rect 3602 43484 3612 43540
rect 3668 43484 5068 43540
rect 5124 43484 5134 43540
rect 16930 43484 16940 43540
rect 16996 43484 17612 43540
rect 17668 43484 17678 43540
rect 20962 43484 20972 43540
rect 21028 43484 33740 43540
rect 33796 43484 41020 43540
rect 41076 43484 41468 43540
rect 41524 43484 52780 43540
rect 52836 43484 53228 43540
rect 53284 43484 53294 43540
rect 19730 43372 19740 43428
rect 19796 43372 22316 43428
rect 22372 43372 22382 43428
rect 40338 43372 40348 43428
rect 40404 43372 42252 43428
rect 42308 43372 42318 43428
rect 42466 43372 42476 43428
rect 42532 43372 43036 43428
rect 43092 43372 44940 43428
rect 44996 43372 45388 43428
rect 45444 43372 45454 43428
rect 46610 43372 46620 43428
rect 46676 43372 46844 43428
rect 46900 43372 48188 43428
rect 48244 43372 48254 43428
rect 19618 43148 19628 43204
rect 19684 43148 20860 43204
rect 20916 43148 22092 43204
rect 22148 43148 22158 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 13010 43036 13020 43092
rect 13076 43036 13916 43092
rect 13972 43036 33180 43092
rect 33236 43036 33246 43092
rect 3602 42924 3612 42980
rect 3668 42924 3948 42980
rect 4004 42924 4014 42980
rect 17266 42924 17276 42980
rect 17332 42924 20188 42980
rect 20244 42924 20254 42980
rect 42242 42924 42252 42980
rect 42308 42924 43596 42980
rect 43652 42924 43662 42980
rect 44146 42924 44156 42980
rect 44212 42924 45612 42980
rect 45668 42924 45678 42980
rect 53106 42924 53116 42980
rect 53172 42924 53900 42980
rect 53956 42924 55132 42980
rect 55188 42924 55198 42980
rect 14914 42812 14924 42868
rect 14980 42812 16828 42868
rect 16884 42812 16894 42868
rect 28354 42812 28364 42868
rect 28420 42812 29932 42868
rect 29988 42812 29998 42868
rect 8754 42700 8764 42756
rect 8820 42700 11788 42756
rect 11844 42700 11854 42756
rect 15922 42700 15932 42756
rect 15988 42700 16492 42756
rect 16548 42700 16558 42756
rect 26002 42700 26012 42756
rect 26068 42700 27132 42756
rect 27188 42700 29148 42756
rect 29204 42700 29214 42756
rect 37762 42700 37772 42756
rect 37828 42700 39452 42756
rect 39508 42700 39518 42756
rect 45602 42700 45612 42756
rect 45668 42700 46620 42756
rect 46676 42700 46686 42756
rect 8306 42588 8316 42644
rect 8372 42588 9100 42644
rect 9156 42588 9166 42644
rect 15932 42588 18060 42644
rect 18116 42588 20300 42644
rect 20356 42588 20366 42644
rect 27682 42588 27692 42644
rect 27748 42588 29708 42644
rect 29764 42588 31276 42644
rect 31332 42588 31342 42644
rect 50194 42588 50204 42644
rect 50260 42588 51660 42644
rect 51716 42588 51726 42644
rect 15932 42532 15988 42588
rect 6066 42476 6076 42532
rect 6132 42476 8988 42532
rect 9044 42476 9054 42532
rect 15922 42476 15932 42532
rect 15988 42476 15998 42532
rect 16818 42476 16828 42532
rect 16884 42476 21420 42532
rect 21476 42476 21486 42532
rect 28466 42476 28476 42532
rect 28532 42476 30940 42532
rect 30996 42476 31006 42532
rect 43698 42476 43708 42532
rect 43764 42476 45164 42532
rect 45220 42476 45948 42532
rect 46004 42476 46396 42532
rect 46452 42476 46462 42532
rect 15810 42364 15820 42420
rect 15876 42364 16268 42420
rect 16324 42364 16334 42420
rect 28018 42364 28028 42420
rect 28084 42364 28364 42420
rect 28420 42364 28430 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 28924 42308 28980 42476
rect 43922 42364 43932 42420
rect 43988 42364 45500 42420
rect 45556 42364 45566 42420
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 8866 42252 8876 42308
rect 8932 42252 9660 42308
rect 9716 42252 9726 42308
rect 28914 42252 28924 42308
rect 28980 42252 28990 42308
rect 9874 42140 9884 42196
rect 9940 42140 10556 42196
rect 10612 42140 10622 42196
rect 17826 42140 17836 42196
rect 17892 42140 20972 42196
rect 21028 42140 21038 42196
rect 28802 42140 28812 42196
rect 28868 42140 30044 42196
rect 30100 42140 30110 42196
rect 35308 42140 36428 42196
rect 36484 42140 38108 42196
rect 38164 42140 38174 42196
rect 22642 42028 22652 42084
rect 22708 42028 24556 42084
rect 24612 42028 24622 42084
rect 27234 42028 27244 42084
rect 27300 42028 27916 42084
rect 27972 42028 28476 42084
rect 28532 42028 28542 42084
rect 33730 42028 33740 42084
rect 33796 42028 34076 42084
rect 34132 42028 34142 42084
rect 35308 41972 35364 42140
rect 35522 42028 35532 42084
rect 35588 42028 39228 42084
rect 39284 42028 39294 42084
rect 8194 41916 8204 41972
rect 8260 41916 8764 41972
rect 8820 41916 9660 41972
rect 9716 41916 9726 41972
rect 13458 41916 13468 41972
rect 13524 41916 14140 41972
rect 14196 41916 14206 41972
rect 14466 41916 14476 41972
rect 14532 41916 15260 41972
rect 15316 41916 15326 41972
rect 15474 41916 15484 41972
rect 15540 41916 20300 41972
rect 20356 41916 21084 41972
rect 21140 41916 21150 41972
rect 28018 41916 28028 41972
rect 28084 41916 29484 41972
rect 29540 41916 29550 41972
rect 33516 41916 35364 41972
rect 38210 41916 38220 41972
rect 38276 41916 38892 41972
rect 38948 41916 38958 41972
rect 40338 41916 40348 41972
rect 40404 41916 41804 41972
rect 41860 41916 41870 41972
rect 43652 41916 45724 41972
rect 45780 41916 46844 41972
rect 46900 41916 46910 41972
rect 49186 41916 49196 41972
rect 49252 41916 50204 41972
rect 50260 41916 52444 41972
rect 52500 41916 53116 41972
rect 53172 41916 53676 41972
rect 53732 41916 54796 41972
rect 54852 41916 56252 41972
rect 56308 41916 56700 41972
rect 56756 41916 56766 41972
rect 14802 41804 14812 41860
rect 14868 41804 17388 41860
rect 17444 41804 17454 41860
rect 19394 41804 19404 41860
rect 19460 41804 21196 41860
rect 21252 41804 21262 41860
rect 28130 41804 28140 41860
rect 28196 41804 30492 41860
rect 30548 41804 30558 41860
rect 33516 41748 33572 41916
rect 43652 41860 43708 41916
rect 38098 41804 38108 41860
rect 38164 41804 43708 41860
rect 55346 41804 55356 41860
rect 55412 41804 57036 41860
rect 57092 41804 57102 41860
rect 57446 41804 57484 41860
rect 57540 41804 57550 41860
rect 2818 41692 2828 41748
rect 2884 41692 3276 41748
rect 3332 41692 15148 41748
rect 15698 41692 15708 41748
rect 15764 41692 16380 41748
rect 16436 41692 19964 41748
rect 20020 41692 20748 41748
rect 20804 41692 20814 41748
rect 24210 41692 24220 41748
rect 24276 41692 26572 41748
rect 26628 41692 26638 41748
rect 26852 41692 33572 41748
rect 33730 41692 33740 41748
rect 33796 41692 36876 41748
rect 36932 41692 36942 41748
rect 57250 41692 57260 41748
rect 57316 41692 57596 41748
rect 57652 41692 57662 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 15092 41524 15148 41692
rect 16930 41580 16940 41636
rect 16996 41580 21420 41636
rect 21476 41580 21486 41636
rect 13794 41468 13804 41524
rect 13860 41468 13870 41524
rect 15092 41468 18060 41524
rect 18116 41468 21308 41524
rect 21364 41468 21374 41524
rect 13804 41412 13860 41468
rect 26852 41412 26908 41692
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 30146 41468 30156 41524
rect 30212 41468 32508 41524
rect 32564 41468 33404 41524
rect 33460 41468 33628 41524
rect 33684 41468 34412 41524
rect 34468 41468 34478 41524
rect 57362 41468 57372 41524
rect 57428 41468 57652 41524
rect 13804 41356 26908 41412
rect 49858 41356 49868 41412
rect 49924 41356 50428 41412
rect 51874 41356 51884 41412
rect 51940 41356 52892 41412
rect 52948 41356 52958 41412
rect 50372 41300 50428 41356
rect 57596 41300 57652 41468
rect 9538 41244 9548 41300
rect 9604 41244 9996 41300
rect 10052 41244 11788 41300
rect 11844 41244 11854 41300
rect 16706 41244 16716 41300
rect 16772 41244 20076 41300
rect 20132 41244 20142 41300
rect 23762 41244 23772 41300
rect 23828 41244 25228 41300
rect 25284 41244 25294 41300
rect 27132 41244 27468 41300
rect 27524 41244 27972 41300
rect 44258 41244 44268 41300
rect 44324 41244 45164 41300
rect 45220 41244 45230 41300
rect 50372 41244 50540 41300
rect 50596 41244 50606 41300
rect 51986 41244 51996 41300
rect 52052 41244 52668 41300
rect 52724 41244 52734 41300
rect 57586 41244 57596 41300
rect 57652 41244 57662 41300
rect 5170 41132 5180 41188
rect 5236 41132 5516 41188
rect 5572 41132 5582 41188
rect 8194 41132 8204 41188
rect 8260 41132 8652 41188
rect 8708 41132 10108 41188
rect 10164 41132 10174 41188
rect 14690 41132 14700 41188
rect 14756 41132 15820 41188
rect 15876 41132 16156 41188
rect 16212 41132 16222 41188
rect 18274 41132 18284 41188
rect 18340 41132 19852 41188
rect 19908 41132 19918 41188
rect 25554 41132 25564 41188
rect 25620 41132 26012 41188
rect 26068 41132 26908 41188
rect 26964 41132 26974 41188
rect 27132 41076 27188 41244
rect 27682 41132 27692 41188
rect 27748 41132 27758 41188
rect 27692 41076 27748 41132
rect 27916 41076 27972 41244
rect 32498 41132 32508 41188
rect 32564 41132 33516 41188
rect 33572 41132 33582 41188
rect 36082 41132 36092 41188
rect 36148 41132 37660 41188
rect 37716 41132 40348 41188
rect 40404 41132 40414 41188
rect 50642 41132 50652 41188
rect 50708 41132 51660 41188
rect 51716 41132 51726 41188
rect 5282 41020 5292 41076
rect 5348 41020 5852 41076
rect 5908 41020 11004 41076
rect 11060 41020 11070 41076
rect 12338 41020 12348 41076
rect 12404 41020 13916 41076
rect 13972 41020 13982 41076
rect 18946 41020 18956 41076
rect 19012 41020 20524 41076
rect 20580 41020 20590 41076
rect 26450 41020 26460 41076
rect 26516 41020 27188 41076
rect 27244 41020 27356 41076
rect 27412 41020 27748 41076
rect 27906 41020 27916 41076
rect 27972 41020 27982 41076
rect 33170 41020 33180 41076
rect 33236 41020 34188 41076
rect 34244 41020 34748 41076
rect 34804 41020 34814 41076
rect 41122 41020 41132 41076
rect 41188 41020 42252 41076
rect 42308 41020 42318 41076
rect 27244 40964 27300 41020
rect 4274 40908 4284 40964
rect 4340 40908 5068 40964
rect 5124 40908 5740 40964
rect 5796 40908 5806 40964
rect 12450 40908 12460 40964
rect 12516 40908 13692 40964
rect 13748 40908 14812 40964
rect 14868 40908 14878 40964
rect 22306 40908 22316 40964
rect 22372 40908 24332 40964
rect 24388 40908 24398 40964
rect 25554 40908 25564 40964
rect 25620 40908 27300 40964
rect 27458 40908 27468 40964
rect 27524 40908 27534 40964
rect 28018 40908 28028 40964
rect 28084 40908 35084 40964
rect 35140 40908 35644 40964
rect 35700 40908 35710 40964
rect 44146 40908 44156 40964
rect 44212 40908 44492 40964
rect 44548 40908 45164 40964
rect 45220 40908 49644 40964
rect 49700 40908 49710 40964
rect 53554 40908 53564 40964
rect 53620 40908 55916 40964
rect 55972 40908 56924 40964
rect 56980 40908 56990 40964
rect 27468 40852 27524 40908
rect 20290 40796 20300 40852
rect 20356 40796 20366 40852
rect 22978 40796 22988 40852
rect 23044 40796 23436 40852
rect 23492 40796 23502 40852
rect 23874 40796 23884 40852
rect 23940 40796 27524 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 12786 40572 12796 40628
rect 12852 40572 14028 40628
rect 14084 40572 14094 40628
rect 20300 40516 20356 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 23090 40684 23100 40740
rect 23156 40684 41804 40740
rect 41860 40684 41870 40740
rect 20962 40572 20972 40628
rect 21028 40572 21420 40628
rect 21476 40572 21486 40628
rect 20972 40516 21028 40572
rect 3042 40460 3052 40516
rect 3108 40460 4060 40516
rect 4116 40460 4126 40516
rect 19170 40460 19180 40516
rect 19236 40460 21028 40516
rect 3938 40348 3948 40404
rect 4004 40348 5292 40404
rect 5348 40348 5358 40404
rect 10994 40348 11004 40404
rect 11060 40348 14476 40404
rect 14532 40348 14542 40404
rect 18386 40348 18396 40404
rect 18452 40348 20300 40404
rect 20356 40348 20366 40404
rect 23100 40292 23156 40684
rect 23314 40572 23324 40628
rect 23380 40572 23772 40628
rect 23828 40572 23838 40628
rect 24434 40572 24444 40628
rect 24500 40572 28924 40628
rect 28980 40572 29708 40628
rect 29764 40572 29774 40628
rect 23884 40460 27804 40516
rect 27860 40460 27870 40516
rect 30258 40460 30268 40516
rect 30324 40460 31164 40516
rect 31220 40460 34972 40516
rect 35028 40460 35038 40516
rect 38098 40460 38108 40516
rect 38164 40460 43372 40516
rect 43428 40460 43438 40516
rect 23884 40404 23940 40460
rect 23874 40348 23884 40404
rect 23940 40348 23950 40404
rect 27234 40348 27244 40404
rect 27300 40348 27580 40404
rect 27636 40348 29484 40404
rect 29540 40348 29550 40404
rect 40226 40348 40236 40404
rect 40292 40348 41244 40404
rect 41300 40348 41468 40404
rect 41524 40348 41534 40404
rect 51650 40348 51660 40404
rect 51716 40348 53116 40404
rect 53172 40348 53182 40404
rect 57446 40348 57484 40404
rect 57540 40348 57550 40404
rect 20738 40236 20748 40292
rect 20804 40236 23156 40292
rect 56018 40236 56028 40292
rect 56084 40236 57036 40292
rect 57092 40236 57102 40292
rect 13794 40124 13804 40180
rect 13860 40124 15148 40180
rect 15204 40124 15214 40180
rect 16482 40124 16492 40180
rect 16548 40124 17388 40180
rect 17444 40124 17454 40180
rect 26338 40124 26348 40180
rect 26404 40124 28588 40180
rect 28644 40124 28654 40180
rect 57474 40012 57484 40068
rect 57540 40012 58380 40068
rect 58436 40012 58446 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 44594 39788 44604 39844
rect 44660 39788 45836 39844
rect 45892 39788 45902 39844
rect 48738 39788 48748 39844
rect 48804 39788 49084 39844
rect 49140 39788 49150 39844
rect 1810 39676 1820 39732
rect 1876 39676 5068 39732
rect 5124 39676 5404 39732
rect 5460 39676 5470 39732
rect 17714 39676 17724 39732
rect 17780 39676 18844 39732
rect 18900 39676 18910 39732
rect 22194 39676 22204 39732
rect 22260 39676 23436 39732
rect 23492 39676 25004 39732
rect 25060 39676 26124 39732
rect 26180 39676 26190 39732
rect 31490 39676 31500 39732
rect 31556 39676 32172 39732
rect 32228 39676 32238 39732
rect 35186 39676 35196 39732
rect 35252 39676 37100 39732
rect 37156 39676 37166 39732
rect 12898 39564 12908 39620
rect 12964 39564 14140 39620
rect 14196 39564 14588 39620
rect 14644 39564 14654 39620
rect 16370 39564 16380 39620
rect 16436 39564 17500 39620
rect 17556 39564 19068 39620
rect 19124 39564 19134 39620
rect 20150 39564 20188 39620
rect 20244 39564 20254 39620
rect 23650 39564 23660 39620
rect 23716 39564 24668 39620
rect 24724 39564 26236 39620
rect 26292 39564 26302 39620
rect 43810 39564 43820 39620
rect 43876 39564 47404 39620
rect 47460 39564 47470 39620
rect 15474 39452 15484 39508
rect 15540 39452 16492 39508
rect 16548 39452 16558 39508
rect 25554 39452 25564 39508
rect 25620 39452 26572 39508
rect 26628 39452 26638 39508
rect 44258 39452 44268 39508
rect 44324 39452 45052 39508
rect 45108 39452 45724 39508
rect 45780 39452 45790 39508
rect 12562 39340 12572 39396
rect 12628 39340 24052 39396
rect 24210 39340 24220 39396
rect 24276 39340 27468 39396
rect 27524 39340 27534 39396
rect 30930 39340 30940 39396
rect 30996 39340 32060 39396
rect 32116 39340 32126 39396
rect 23996 39284 24052 39340
rect 23996 39228 30156 39284
rect 30212 39228 30222 39284
rect 42242 39228 42252 39284
rect 42308 39228 48748 39284
rect 48804 39228 48972 39284
rect 49028 39228 49038 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 22418 39116 22428 39172
rect 22484 39116 23212 39172
rect 23268 39116 23278 39172
rect 7858 39004 7868 39060
rect 7924 39004 12348 39060
rect 12404 39004 12414 39060
rect 26674 39004 26684 39060
rect 26740 39004 27692 39060
rect 27748 39004 27758 39060
rect 30370 39004 30380 39060
rect 30436 39004 31276 39060
rect 31332 39004 31342 39060
rect 54114 39004 54124 39060
rect 54180 39004 56364 39060
rect 56420 39004 56812 39060
rect 56868 39004 56878 39060
rect 12002 38892 12012 38948
rect 12068 38892 12908 38948
rect 12964 38892 12974 38948
rect 18834 38892 18844 38948
rect 18900 38892 19292 38948
rect 19348 38892 20412 38948
rect 20468 38892 20478 38948
rect 24322 38892 24332 38948
rect 24388 38892 27132 38948
rect 27188 38892 27198 38948
rect 36754 38892 36764 38948
rect 36820 38892 39004 38948
rect 39060 38892 39070 38948
rect 5842 38780 5852 38836
rect 5908 38780 6636 38836
rect 6692 38780 7868 38836
rect 7924 38780 7934 38836
rect 11442 38780 11452 38836
rect 11508 38780 12572 38836
rect 12628 38780 13132 38836
rect 13188 38780 13198 38836
rect 15810 38780 15820 38836
rect 15876 38780 16828 38836
rect 16884 38780 18060 38836
rect 18116 38780 18126 38836
rect 23874 38780 23884 38836
rect 23940 38780 26348 38836
rect 26404 38780 26414 38836
rect 26852 38780 28028 38836
rect 28084 38780 28094 38836
rect 30034 38780 30044 38836
rect 30100 38780 30940 38836
rect 30996 38780 31006 38836
rect 37090 38780 37100 38836
rect 37156 38780 46060 38836
rect 46116 38780 46228 38836
rect 57586 38780 57596 38836
rect 57652 38780 58044 38836
rect 58100 38780 58110 38836
rect 26852 38724 26908 38780
rect 46172 38724 46228 38780
rect 4162 38668 4172 38724
rect 4228 38668 7532 38724
rect 7588 38668 7598 38724
rect 10770 38668 10780 38724
rect 10836 38668 11676 38724
rect 11732 38668 12460 38724
rect 12516 38668 12526 38724
rect 17714 38668 17724 38724
rect 17780 38668 17948 38724
rect 18004 38668 18620 38724
rect 18676 38668 18686 38724
rect 24546 38668 24556 38724
rect 24612 38668 25676 38724
rect 25732 38668 25742 38724
rect 26002 38668 26012 38724
rect 26068 38668 26908 38724
rect 29922 38668 29932 38724
rect 29988 38668 34748 38724
rect 34804 38668 34814 38724
rect 35196 38668 37548 38724
rect 37604 38668 37614 38724
rect 46162 38668 46172 38724
rect 46228 38668 46238 38724
rect 49410 38668 49420 38724
rect 49476 38668 53676 38724
rect 53732 38668 53742 38724
rect 35196 38612 35252 38668
rect 6402 38556 6412 38612
rect 6468 38556 7420 38612
rect 7476 38556 7980 38612
rect 8036 38556 8046 38612
rect 12226 38556 12236 38612
rect 12292 38556 12572 38612
rect 12628 38556 15372 38612
rect 15428 38556 15438 38612
rect 18498 38556 18508 38612
rect 18564 38556 19852 38612
rect 19908 38556 19918 38612
rect 28354 38556 28364 38612
rect 28420 38556 30828 38612
rect 30884 38556 30894 38612
rect 31052 38556 35252 38612
rect 39666 38556 39676 38612
rect 39732 38556 40236 38612
rect 40292 38556 40302 38612
rect 7074 38444 7084 38500
rect 7140 38444 13524 38500
rect 15138 38444 15148 38500
rect 15204 38444 15484 38500
rect 15540 38444 15550 38500
rect 26114 38444 26124 38500
rect 26180 38444 26908 38500
rect 26964 38444 29260 38500
rect 29316 38444 29326 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 13468 38388 13524 38444
rect 31052 38388 31108 38556
rect 31938 38444 31948 38500
rect 32004 38444 34076 38500
rect 34132 38444 34142 38500
rect 57698 38444 57708 38500
rect 57764 38444 58268 38500
rect 58324 38444 58334 38500
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 59200 38388 60000 38416
rect 11778 38332 11788 38388
rect 11844 38332 13244 38388
rect 13300 38332 13310 38388
rect 13468 38332 20188 38388
rect 20244 38332 21308 38388
rect 21364 38332 21374 38388
rect 26786 38332 26796 38388
rect 26852 38332 31108 38388
rect 58034 38332 58044 38388
rect 58100 38332 60000 38388
rect 59200 38304 60000 38332
rect 9874 38220 9884 38276
rect 9940 38220 11900 38276
rect 11956 38220 11966 38276
rect 14578 38220 14588 38276
rect 14644 38220 15372 38276
rect 15428 38220 15438 38276
rect 16034 38220 16044 38276
rect 16100 38220 18956 38276
rect 19012 38220 20636 38276
rect 20692 38220 20702 38276
rect 15586 38108 15596 38164
rect 15652 38108 15764 38164
rect 16146 38108 16156 38164
rect 16212 38108 16604 38164
rect 16660 38108 17948 38164
rect 18004 38108 18014 38164
rect 24658 38108 24668 38164
rect 24724 38108 27020 38164
rect 27076 38108 27086 38164
rect 37874 38108 37884 38164
rect 37940 38108 38780 38164
rect 38836 38108 38846 38164
rect 45714 38108 45724 38164
rect 45780 38108 46396 38164
rect 46452 38108 46462 38164
rect 4050 37996 4060 38052
rect 4116 37996 11116 38052
rect 11172 37996 11182 38052
rect 14018 37996 14028 38052
rect 14084 37996 14094 38052
rect 14802 37996 14812 38052
rect 14868 37996 15484 38052
rect 15540 37996 15550 38052
rect 14028 37828 14084 37996
rect 15708 37940 15764 38108
rect 17602 37996 17612 38052
rect 17668 37996 18508 38052
rect 18564 37996 18574 38052
rect 26562 37996 26572 38052
rect 26628 37996 27468 38052
rect 27524 37996 28252 38052
rect 28308 37996 28588 38052
rect 28644 37996 29148 38052
rect 29204 37996 29214 38052
rect 46022 37996 46060 38052
rect 46116 37996 46126 38052
rect 54898 37996 54908 38052
rect 54964 37996 55356 38052
rect 55412 37996 56700 38052
rect 56756 37996 56766 38052
rect 15708 37884 17052 37940
rect 17108 37884 18956 37940
rect 19012 37884 19022 37940
rect 22978 37884 22988 37940
rect 23044 37884 23996 37940
rect 24052 37884 24062 37940
rect 27570 37884 27580 37940
rect 27636 37884 28140 37940
rect 28196 37884 29260 37940
rect 29316 37884 29326 37940
rect 30594 37884 30604 37940
rect 30660 37884 31500 37940
rect 31556 37884 31566 37940
rect 33954 37884 33964 37940
rect 34020 37884 37212 37940
rect 37268 37884 38668 37940
rect 38724 37884 38734 37940
rect 46610 37884 46620 37940
rect 46676 37884 48524 37940
rect 48580 37884 48590 37940
rect 14028 37772 15260 37828
rect 15316 37772 18620 37828
rect 18676 37772 18686 37828
rect 26002 37772 26012 37828
rect 26068 37772 28364 37828
rect 28420 37772 28430 37828
rect 28690 37772 28700 37828
rect 28756 37772 30828 37828
rect 30884 37772 30894 37828
rect 34514 37772 34524 37828
rect 34580 37772 35308 37828
rect 36866 37772 36876 37828
rect 36932 37772 37436 37828
rect 37492 37772 37502 37828
rect 15586 37660 15596 37716
rect 15652 37660 15932 37716
rect 15988 37660 15998 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 35252 37604 35308 37772
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 23538 37548 23548 37604
rect 23604 37548 23996 37604
rect 24052 37548 24062 37604
rect 35252 37548 35532 37604
rect 35588 37548 37828 37604
rect 2706 37436 2716 37492
rect 2772 37436 3612 37492
rect 3668 37436 3678 37492
rect 19618 37436 19628 37492
rect 19684 37436 20188 37492
rect 20244 37436 20254 37492
rect 23874 37436 23884 37492
rect 23940 37436 25340 37492
rect 25396 37436 27580 37492
rect 27636 37436 27646 37492
rect 31266 37436 31276 37492
rect 31332 37436 37100 37492
rect 37156 37436 37166 37492
rect 37772 37380 37828 37548
rect 37986 37436 37996 37492
rect 38052 37436 38062 37492
rect 3042 37324 3052 37380
rect 3108 37324 3948 37380
rect 4004 37324 4014 37380
rect 8418 37324 8428 37380
rect 8484 37324 8764 37380
rect 8820 37324 8830 37380
rect 9874 37324 9884 37380
rect 9940 37324 10892 37380
rect 10948 37324 10958 37380
rect 11330 37324 11340 37380
rect 11396 37324 12460 37380
rect 12516 37324 12526 37380
rect 14802 37324 14812 37380
rect 14868 37324 16828 37380
rect 16884 37324 16894 37380
rect 19394 37324 19404 37380
rect 19460 37324 20300 37380
rect 20356 37324 20366 37380
rect 26114 37324 26124 37380
rect 26180 37324 27132 37380
rect 27188 37324 27198 37380
rect 30258 37324 30268 37380
rect 30324 37324 31388 37380
rect 31444 37324 34412 37380
rect 34468 37324 34478 37380
rect 34626 37324 34636 37380
rect 34692 37324 35756 37380
rect 35812 37324 35822 37380
rect 37762 37324 37772 37380
rect 37828 37324 37838 37380
rect 11340 37268 11396 37324
rect 3154 37212 3164 37268
rect 3220 37212 3724 37268
rect 3780 37212 3790 37268
rect 4610 37212 4620 37268
rect 4676 37212 5180 37268
rect 5236 37212 7868 37268
rect 7924 37212 7934 37268
rect 8530 37212 8540 37268
rect 8596 37212 9324 37268
rect 9380 37212 11396 37268
rect 15474 37212 15484 37268
rect 15540 37212 16044 37268
rect 16100 37212 16110 37268
rect 16370 37212 16380 37268
rect 16436 37212 17276 37268
rect 17332 37212 17342 37268
rect 19058 37212 19068 37268
rect 19124 37212 20412 37268
rect 20468 37212 20478 37268
rect 26786 37212 26796 37268
rect 26852 37212 29372 37268
rect 29428 37212 29438 37268
rect 33506 37212 33516 37268
rect 33572 37212 34300 37268
rect 34356 37212 35644 37268
rect 35700 37212 35710 37268
rect 8754 37100 8764 37156
rect 8820 37100 9436 37156
rect 9492 37100 9502 37156
rect 15810 37100 15820 37156
rect 15876 37100 16268 37156
rect 16324 37100 16334 37156
rect 18498 37100 18508 37156
rect 18564 37100 19740 37156
rect 19796 37100 20748 37156
rect 20804 37100 20814 37156
rect 22866 37100 22876 37156
rect 22932 37100 25228 37156
rect 25284 37100 25294 37156
rect 31490 37100 31500 37156
rect 31556 37100 34076 37156
rect 34132 37100 34142 37156
rect 9090 36988 9100 37044
rect 9156 36988 9548 37044
rect 9604 36988 10220 37044
rect 10276 36988 10556 37044
rect 10612 36988 10622 37044
rect 10994 36988 11004 37044
rect 11060 36988 11900 37044
rect 11956 36988 11966 37044
rect 23996 36932 24052 37100
rect 37996 37044 38052 37436
rect 38770 37324 38780 37380
rect 38836 37324 39564 37380
rect 39620 37324 39630 37380
rect 39218 37100 39228 37156
rect 39284 37100 39676 37156
rect 39732 37100 40908 37156
rect 40964 37100 40974 37156
rect 41234 37100 41244 37156
rect 41300 37100 43036 37156
rect 43092 37100 43102 37156
rect 33058 36988 33068 37044
rect 33124 36988 35980 37044
rect 36036 36988 37772 37044
rect 37828 36988 38052 37044
rect 17154 36876 17164 36932
rect 17220 36876 20300 36932
rect 20356 36876 20366 36932
rect 23986 36876 23996 36932
rect 24052 36876 24062 36932
rect 25218 36876 25228 36932
rect 25284 36876 26012 36932
rect 26068 36876 26078 36932
rect 37314 36876 37324 36932
rect 37380 36876 37660 36932
rect 37716 36876 37726 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 8754 36540 8764 36596
rect 8820 36540 9772 36596
rect 9828 36540 9838 36596
rect 15922 36428 15932 36484
rect 15988 36428 16828 36484
rect 16884 36428 17948 36484
rect 18004 36428 18014 36484
rect 24322 36428 24332 36484
rect 24388 36428 26908 36484
rect 26964 36428 26974 36484
rect 35410 36428 35420 36484
rect 35476 36428 37212 36484
rect 37268 36428 38556 36484
rect 38612 36428 39228 36484
rect 39284 36428 39294 36484
rect 57026 36428 57036 36484
rect 57092 36428 57932 36484
rect 57988 36428 57998 36484
rect 8866 36316 8876 36372
rect 8932 36316 11564 36372
rect 11620 36316 11900 36372
rect 11956 36316 11966 36372
rect 15698 36316 15708 36372
rect 15764 36316 18844 36372
rect 18900 36316 18910 36372
rect 36082 36316 36092 36372
rect 36148 36316 37996 36372
rect 38052 36316 38062 36372
rect 49970 36316 49980 36372
rect 50036 36316 50316 36372
rect 50372 36316 50382 36372
rect 55570 36316 55580 36372
rect 55636 36316 56700 36372
rect 56756 36316 56766 36372
rect 10770 36204 10780 36260
rect 10836 36204 12684 36260
rect 12740 36204 12750 36260
rect 31154 36204 31164 36260
rect 31220 36204 32060 36260
rect 32116 36204 32126 36260
rect 56018 36204 56028 36260
rect 56084 36204 57148 36260
rect 57204 36204 57214 36260
rect 9874 36092 9884 36148
rect 9940 36092 11004 36148
rect 11060 36092 11070 36148
rect 33282 36092 33292 36148
rect 33348 36092 35084 36148
rect 35140 36092 35980 36148
rect 36036 36092 36046 36148
rect 36530 36092 36540 36148
rect 36596 36092 38220 36148
rect 38276 36092 38286 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 24210 35980 24220 36036
rect 24276 35980 25228 36036
rect 25284 35980 25294 36036
rect 22754 35868 22764 35924
rect 22820 35868 23324 35924
rect 23380 35868 27244 35924
rect 27300 35868 27310 35924
rect 8642 35644 8652 35700
rect 8708 35644 11340 35700
rect 11396 35644 11406 35700
rect 14914 35644 14924 35700
rect 14980 35644 16156 35700
rect 16212 35644 16222 35700
rect 22754 35644 22764 35700
rect 22820 35644 23660 35700
rect 23716 35644 23726 35700
rect 29698 35644 29708 35700
rect 29764 35644 30492 35700
rect 30548 35644 30558 35700
rect 32498 35644 32508 35700
rect 32564 35644 33964 35700
rect 34020 35644 34030 35700
rect 42466 35644 42476 35700
rect 42532 35644 45500 35700
rect 45556 35644 45566 35700
rect 52210 35644 52220 35700
rect 52276 35644 52892 35700
rect 52948 35644 52958 35700
rect 55346 35644 55356 35700
rect 55412 35644 56476 35700
rect 56532 35644 56542 35700
rect 56914 35644 56924 35700
rect 56980 35644 57820 35700
rect 57876 35644 57886 35700
rect 2258 35532 2268 35588
rect 2324 35532 21308 35588
rect 21364 35532 21374 35588
rect 25442 35532 25452 35588
rect 25508 35532 27356 35588
rect 27412 35532 27422 35588
rect 32162 35532 32172 35588
rect 32228 35532 34188 35588
rect 34244 35532 36540 35588
rect 36596 35532 36606 35588
rect 17490 35420 17500 35476
rect 17556 35420 19180 35476
rect 19236 35420 20860 35476
rect 20916 35420 20926 35476
rect 50082 35420 50092 35476
rect 50148 35420 50316 35476
rect 50372 35420 51772 35476
rect 51828 35420 53116 35476
rect 53172 35420 53182 35476
rect 8754 35308 8764 35364
rect 8820 35308 9436 35364
rect 9492 35308 9502 35364
rect 23314 35308 23324 35364
rect 23380 35308 25676 35364
rect 25732 35308 25742 35364
rect 35858 35308 35868 35364
rect 35924 35308 36988 35364
rect 37044 35308 38332 35364
rect 38388 35308 38398 35364
rect 54002 35308 54012 35364
rect 54068 35308 56812 35364
rect 56868 35308 57708 35364
rect 57764 35308 57774 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 37538 35084 37548 35140
rect 37604 35084 38332 35140
rect 38388 35084 38398 35140
rect 0 35028 800 35056
rect 0 34972 1820 35028
rect 1876 34972 1886 35028
rect 27906 34972 27916 35028
rect 27972 34972 29148 35028
rect 29204 34972 29214 35028
rect 30930 34972 30940 35028
rect 30996 34972 31612 35028
rect 31668 34972 34748 35028
rect 34804 34972 35756 35028
rect 35812 34972 35822 35028
rect 36194 34972 36204 35028
rect 36260 34972 38220 35028
rect 38276 34972 38286 35028
rect 45042 34972 45052 35028
rect 45108 34972 45500 35028
rect 45556 34972 45566 35028
rect 48850 34972 48860 35028
rect 48916 34972 49980 35028
rect 50036 34972 50046 35028
rect 0 34944 800 34972
rect 7858 34860 7868 34916
rect 7924 34860 8428 34916
rect 8484 34860 8494 34916
rect 9538 34860 9548 34916
rect 9604 34860 9996 34916
rect 10052 34860 10062 34916
rect 11106 34860 11116 34916
rect 11172 34860 13468 34916
rect 13524 34860 13534 34916
rect 16594 34860 16604 34916
rect 16660 34860 17836 34916
rect 17892 34860 17902 34916
rect 29810 34860 29820 34916
rect 29876 34860 30716 34916
rect 30772 34860 30782 34916
rect 12898 34748 12908 34804
rect 12964 34748 13804 34804
rect 13860 34748 13870 34804
rect 17938 34748 17948 34804
rect 18004 34748 18508 34804
rect 18564 34748 18574 34804
rect 31042 34748 31052 34804
rect 31108 34748 35084 34804
rect 35140 34748 37100 34804
rect 37156 34748 37166 34804
rect 42354 34748 42364 34804
rect 42420 34748 43820 34804
rect 43876 34748 44268 34804
rect 44324 34748 44334 34804
rect 10546 34636 10556 34692
rect 10612 34636 11452 34692
rect 11508 34636 12684 34692
rect 12740 34636 12750 34692
rect 29362 34636 29372 34692
rect 29428 34636 30044 34692
rect 30100 34636 30110 34692
rect 53442 34636 53452 34692
rect 53508 34636 54012 34692
rect 54068 34636 54078 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 28354 34412 28364 34468
rect 28420 34412 38780 34468
rect 38836 34412 38846 34468
rect 40226 34412 40236 34468
rect 40292 34412 42700 34468
rect 42756 34412 43596 34468
rect 43652 34412 44492 34468
rect 44548 34412 44558 34468
rect 41458 34300 41468 34356
rect 41524 34300 42364 34356
rect 42420 34300 42430 34356
rect 47730 34300 47740 34356
rect 47796 34300 51100 34356
rect 51156 34300 51166 34356
rect 8754 34188 8764 34244
rect 8820 34188 10780 34244
rect 10836 34188 10846 34244
rect 29586 34188 29596 34244
rect 29652 34188 30268 34244
rect 30324 34188 30940 34244
rect 30996 34188 31006 34244
rect 9874 34076 9884 34132
rect 9940 34076 13916 34132
rect 13972 34076 13982 34132
rect 17602 34076 17612 34132
rect 17668 34076 18284 34132
rect 18340 34076 18350 34132
rect 19170 34076 19180 34132
rect 19236 34076 19516 34132
rect 19572 34076 19582 34132
rect 31826 34076 31836 34132
rect 31892 34076 33628 34132
rect 33684 34076 33694 34132
rect 34962 34076 34972 34132
rect 35028 34076 36764 34132
rect 36820 34076 37996 34132
rect 38052 34076 38062 34132
rect 38210 34076 38220 34132
rect 38276 34076 38332 34132
rect 38388 34076 40348 34132
rect 40404 34076 41020 34132
rect 41076 34076 41086 34132
rect 41234 34076 41244 34132
rect 41300 34076 42028 34132
rect 42084 34076 42094 34132
rect 44594 34076 44604 34132
rect 44660 34076 45052 34132
rect 45108 34076 45724 34132
rect 45780 34076 45790 34132
rect 55570 34076 55580 34132
rect 55636 34076 56924 34132
rect 56980 34076 57260 34132
rect 57316 34076 57326 34132
rect 5842 33964 5852 34020
rect 5908 33964 29820 34020
rect 29876 33964 29886 34020
rect 34402 33964 34412 34020
rect 34468 33964 36876 34020
rect 36932 33964 37436 34020
rect 37492 33964 37502 34020
rect 39666 33964 39676 34020
rect 39732 33964 41916 34020
rect 41972 33964 41982 34020
rect 13122 33852 13132 33908
rect 13188 33852 13692 33908
rect 13748 33852 13758 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 10546 33628 10556 33684
rect 10612 33628 12012 33684
rect 12068 33628 13692 33684
rect 13748 33628 14812 33684
rect 14868 33628 14878 33684
rect 28354 33628 28364 33684
rect 28420 33628 28812 33684
rect 28868 33628 28878 33684
rect 31826 33628 31836 33684
rect 31892 33628 32956 33684
rect 33012 33628 33022 33684
rect 48934 33628 48972 33684
rect 49028 33628 49038 33684
rect 22754 33516 22764 33572
rect 22820 33516 23548 33572
rect 23604 33516 23614 33572
rect 34178 33516 34188 33572
rect 34244 33516 34972 33572
rect 35028 33516 35038 33572
rect 41682 33516 41692 33572
rect 41748 33516 42364 33572
rect 42420 33516 42430 33572
rect 49046 33516 49084 33572
rect 49140 33516 49150 33572
rect 21634 33404 21644 33460
rect 21700 33404 25116 33460
rect 25172 33404 25182 33460
rect 29474 33404 29484 33460
rect 29540 33404 31500 33460
rect 31556 33404 31566 33460
rect 39106 33404 39116 33460
rect 39172 33404 49420 33460
rect 49476 33404 49486 33460
rect 57138 33404 57148 33460
rect 57204 33404 57214 33460
rect 57148 33348 57204 33404
rect 10882 33292 10892 33348
rect 10948 33292 11676 33348
rect 11732 33292 11742 33348
rect 18834 33292 18844 33348
rect 18900 33292 19516 33348
rect 19572 33292 19582 33348
rect 28130 33292 28140 33348
rect 28196 33292 28924 33348
rect 28980 33292 30436 33348
rect 31266 33292 31276 33348
rect 31332 33292 31612 33348
rect 31668 33292 33852 33348
rect 33908 33292 34300 33348
rect 34356 33292 34366 33348
rect 34524 33292 38892 33348
rect 38948 33292 38958 33348
rect 39890 33292 39900 33348
rect 39956 33292 43260 33348
rect 43316 33292 43326 33348
rect 51874 33292 51884 33348
rect 51940 33292 53788 33348
rect 53844 33292 53854 33348
rect 55010 33292 55020 33348
rect 55076 33292 57484 33348
rect 57540 33292 57550 33348
rect 30380 33236 30436 33292
rect 34524 33236 34580 33292
rect 15922 33180 15932 33236
rect 15988 33180 18620 33236
rect 18676 33180 18686 33236
rect 22166 33180 22204 33236
rect 22260 33180 22270 33236
rect 25778 33180 25788 33236
rect 25844 33180 28252 33236
rect 28308 33180 28318 33236
rect 30380 33180 34580 33236
rect 38098 33180 38108 33236
rect 38164 33180 38668 33236
rect 42354 33180 42364 33236
rect 42420 33180 43372 33236
rect 43428 33180 43438 33236
rect 51986 33180 51996 33236
rect 52052 33180 53452 33236
rect 53508 33180 53518 33236
rect 54002 33180 54012 33236
rect 54068 33180 57148 33236
rect 57204 33180 57214 33236
rect 38612 33124 38668 33180
rect 12786 33068 12796 33124
rect 12852 33068 13468 33124
rect 13524 33068 13534 33124
rect 18498 33068 18508 33124
rect 18564 33068 19404 33124
rect 19460 33068 19470 33124
rect 21410 33068 21420 33124
rect 21476 33068 23884 33124
rect 23940 33068 24668 33124
rect 24724 33068 24734 33124
rect 27794 33068 27804 33124
rect 27860 33068 28700 33124
rect 28756 33068 29372 33124
rect 29428 33068 29438 33124
rect 34962 33068 34972 33124
rect 35028 33068 37100 33124
rect 37156 33068 37166 33124
rect 38612 33068 45948 33124
rect 46004 33068 46014 33124
rect 57026 33068 57036 33124
rect 57092 33068 57596 33124
rect 57652 33068 58044 33124
rect 58100 33068 58110 33124
rect 19058 32956 19068 33012
rect 19124 32956 19516 33012
rect 19572 32956 19582 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 37202 32732 37212 32788
rect 37268 32732 38108 32788
rect 38164 32732 39452 32788
rect 39508 32732 39518 32788
rect 53890 32732 53900 32788
rect 53956 32732 54908 32788
rect 54964 32732 55580 32788
rect 55636 32732 55646 32788
rect 8530 32620 8540 32676
rect 8596 32620 12460 32676
rect 12516 32620 12526 32676
rect 31826 32620 31836 32676
rect 31892 32620 32284 32676
rect 32340 32620 32350 32676
rect 34850 32620 34860 32676
rect 34916 32620 36988 32676
rect 37044 32620 37054 32676
rect 52210 32620 52220 32676
rect 52276 32620 52668 32676
rect 52724 32620 54796 32676
rect 54852 32620 54862 32676
rect 33628 32508 37436 32564
rect 37492 32508 37502 32564
rect 37650 32508 37660 32564
rect 37716 32508 46732 32564
rect 46788 32508 46798 32564
rect 47394 32508 47404 32564
rect 47460 32508 48972 32564
rect 49028 32508 49038 32564
rect 49634 32508 49644 32564
rect 49700 32508 50428 32564
rect 50484 32508 50494 32564
rect 33628 32452 33684 32508
rect 8754 32396 8764 32452
rect 8820 32396 9884 32452
rect 9940 32396 9950 32452
rect 19394 32396 19404 32452
rect 19460 32396 20748 32452
rect 20804 32396 20814 32452
rect 31714 32396 31724 32452
rect 31780 32396 33628 32452
rect 33684 32396 33694 32452
rect 34738 32396 34748 32452
rect 34804 32396 36204 32452
rect 36260 32396 36270 32452
rect 39340 32396 39900 32452
rect 39956 32396 39966 32452
rect 43586 32396 43596 32452
rect 43652 32396 44044 32452
rect 44100 32396 44110 32452
rect 39340 32340 39396 32396
rect 20178 32284 20188 32340
rect 20244 32284 39396 32340
rect 39554 32284 39564 32340
rect 39620 32284 42028 32340
rect 42084 32284 42094 32340
rect 36194 32172 36204 32228
rect 36260 32172 38892 32228
rect 38948 32172 49084 32228
rect 49140 32172 49532 32228
rect 49588 32172 49598 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 32274 32060 32284 32116
rect 32340 32060 34076 32116
rect 34132 32060 34860 32116
rect 34916 32060 34926 32116
rect 51426 32060 51436 32116
rect 51492 32060 52780 32116
rect 52836 32060 55244 32116
rect 55300 32060 56028 32116
rect 56084 32060 58156 32116
rect 58212 32060 58222 32116
rect 17938 31948 17948 32004
rect 18004 31948 20188 32004
rect 20244 31948 20254 32004
rect 34290 31948 34300 32004
rect 34356 31948 35308 32004
rect 35364 31948 35374 32004
rect 35746 31948 35756 32004
rect 35812 31948 37212 32004
rect 37268 31948 37278 32004
rect 7970 31836 7980 31892
rect 8036 31836 8876 31892
rect 8932 31836 8942 31892
rect 13010 31836 13020 31892
rect 13076 31836 13916 31892
rect 13972 31836 13982 31892
rect 17490 31836 17500 31892
rect 17556 31836 18956 31892
rect 19012 31836 19022 31892
rect 24098 31836 24108 31892
rect 24164 31836 26796 31892
rect 26852 31836 26862 31892
rect 31490 31836 31500 31892
rect 31556 31836 33068 31892
rect 33124 31836 34748 31892
rect 34804 31836 34814 31892
rect 37874 31836 37884 31892
rect 37940 31836 45388 31892
rect 45444 31836 45454 31892
rect 50082 31836 50092 31892
rect 50148 31836 50876 31892
rect 50932 31836 51772 31892
rect 51828 31836 51838 31892
rect 30482 31724 30492 31780
rect 30548 31724 32060 31780
rect 32116 31724 34300 31780
rect 34356 31724 34366 31780
rect 35410 31724 35420 31780
rect 35476 31724 35868 31780
rect 35924 31724 37996 31780
rect 38052 31724 38444 31780
rect 38500 31724 38510 31780
rect 44258 31724 44268 31780
rect 44324 31724 45164 31780
rect 45220 31724 45230 31780
rect 49298 31724 49308 31780
rect 49364 31724 50428 31780
rect 50484 31724 50494 31780
rect 8082 31612 8092 31668
rect 8148 31612 8988 31668
rect 9044 31612 9772 31668
rect 9828 31612 9838 31668
rect 12562 31612 12572 31668
rect 12628 31612 14252 31668
rect 14308 31612 14318 31668
rect 35186 31612 35196 31668
rect 35252 31612 38556 31668
rect 38612 31612 38622 31668
rect 47506 31612 47516 31668
rect 47572 31612 49420 31668
rect 49476 31612 49486 31668
rect 50754 31500 50764 31556
rect 50820 31500 53116 31556
rect 53172 31500 53182 31556
rect 59200 31444 60000 31472
rect 15026 31388 15036 31444
rect 15092 31388 16716 31444
rect 16772 31388 16782 31444
rect 58146 31388 58156 31444
rect 58212 31388 60000 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 59200 31360 60000 31388
rect 31042 31164 31052 31220
rect 31108 31164 32060 31220
rect 32116 31164 32126 31220
rect 38612 31164 52332 31220
rect 52388 31164 52398 31220
rect 38612 31108 38668 31164
rect 22166 31052 22204 31108
rect 22260 31052 22270 31108
rect 29922 31052 29932 31108
rect 29988 31052 38668 31108
rect 7634 30940 7644 30996
rect 7700 30940 8540 30996
rect 8596 30940 8606 30996
rect 8866 30940 8876 30996
rect 8932 30940 11788 30996
rect 11844 30940 12908 30996
rect 12964 30940 12974 30996
rect 21970 30940 21980 30996
rect 22036 30940 22540 30996
rect 22596 30940 22606 30996
rect 22866 30940 22876 30996
rect 22932 30940 23436 30996
rect 23492 30940 23996 30996
rect 24052 30940 24062 30996
rect 55346 30940 55356 30996
rect 55412 30940 56588 30996
rect 56644 30940 56924 30996
rect 56980 30940 56990 30996
rect 10210 30828 10220 30884
rect 10276 30828 11452 30884
rect 11508 30828 12684 30884
rect 12740 30828 12750 30884
rect 20290 30828 20300 30884
rect 20356 30828 21196 30884
rect 21252 30828 22092 30884
rect 22148 30828 29708 30884
rect 29764 30828 29774 30884
rect 50194 30828 50204 30884
rect 50260 30828 50876 30884
rect 50932 30828 50942 30884
rect 9314 30716 9324 30772
rect 9380 30716 10444 30772
rect 10500 30716 11116 30772
rect 11172 30716 11182 30772
rect 28578 30716 28588 30772
rect 28644 30716 30156 30772
rect 30212 30716 34860 30772
rect 34916 30716 34926 30772
rect 48402 30604 48412 30660
rect 48468 30604 49868 30660
rect 49924 30604 49934 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 8194 30380 8204 30436
rect 8260 30380 8988 30436
rect 9044 30380 11004 30436
rect 11060 30380 11070 30436
rect 13570 30380 13580 30436
rect 13636 30380 13860 30436
rect 22194 30380 22204 30436
rect 22260 30380 22988 30436
rect 23044 30380 23054 30436
rect 51538 30380 51548 30436
rect 51604 30380 55132 30436
rect 55188 30380 55198 30436
rect 8082 30268 8092 30324
rect 8148 30268 8428 30324
rect 8484 30268 9212 30324
rect 9268 30268 9772 30324
rect 9828 30268 11116 30324
rect 11172 30268 11182 30324
rect 13804 30212 13860 30380
rect 29586 30268 29596 30324
rect 29652 30268 30156 30324
rect 30212 30268 30222 30324
rect 46946 30268 46956 30324
rect 47012 30268 49980 30324
rect 50036 30268 50316 30324
rect 50372 30268 50382 30324
rect 51762 30268 51772 30324
rect 51828 30268 52668 30324
rect 52724 30268 52734 30324
rect 11890 30156 11900 30212
rect 11956 30156 13580 30212
rect 13636 30156 13646 30212
rect 13804 30156 13972 30212
rect 14802 30156 14812 30212
rect 14868 30156 15708 30212
rect 15764 30156 15774 30212
rect 16258 30156 16268 30212
rect 16324 30156 19180 30212
rect 19236 30156 19246 30212
rect 21858 30156 21868 30212
rect 21924 30156 22316 30212
rect 22372 30156 22382 30212
rect 23986 30156 23996 30212
rect 24052 30156 25900 30212
rect 25956 30156 28140 30212
rect 28196 30156 28206 30212
rect 32274 30156 32284 30212
rect 32340 30156 33180 30212
rect 33236 30156 33246 30212
rect 42354 30156 42364 30212
rect 42420 30156 45276 30212
rect 45332 30156 45612 30212
rect 45668 30156 45678 30212
rect 49858 30156 49868 30212
rect 49924 30156 50876 30212
rect 50932 30156 50942 30212
rect 13916 29988 13972 30156
rect 22316 30100 22372 30156
rect 22316 30044 24220 30100
rect 24276 30044 24286 30100
rect 30482 30044 30492 30100
rect 30548 30044 31276 30100
rect 31332 30044 31342 30100
rect 35410 30044 35420 30100
rect 35476 30044 48972 30100
rect 49028 30044 49038 30100
rect 13906 29932 13916 29988
rect 13972 29932 13982 29988
rect 15586 29932 15596 29988
rect 15652 29932 16604 29988
rect 16660 29932 18060 29988
rect 18116 29932 20244 29988
rect 22194 29932 22204 29988
rect 22260 29932 22764 29988
rect 22820 29932 22830 29988
rect 24434 29932 24444 29988
rect 24500 29932 25452 29988
rect 25508 29932 25518 29988
rect 29922 29932 29932 29988
rect 29988 29932 30604 29988
rect 30660 29932 30670 29988
rect 31378 29932 31388 29988
rect 31444 29932 34524 29988
rect 34580 29932 34590 29988
rect 38882 29932 38892 29988
rect 38948 29932 40348 29988
rect 40404 29932 41916 29988
rect 41972 29932 41982 29988
rect 53218 29932 53228 29988
rect 53284 29932 54572 29988
rect 54628 29932 54638 29988
rect 54898 29932 54908 29988
rect 54964 29932 57036 29988
rect 57092 29932 57708 29988
rect 57764 29932 57774 29988
rect 20188 29876 20244 29932
rect 24444 29876 24500 29932
rect 20188 29820 24500 29876
rect 37762 29820 37772 29876
rect 37828 29820 39788 29876
rect 39844 29820 39854 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 10658 29708 10668 29764
rect 10724 29708 17948 29764
rect 18004 29708 18014 29764
rect 21298 29708 21308 29764
rect 21364 29708 35084 29764
rect 35140 29708 35150 29764
rect 8978 29596 8988 29652
rect 9044 29596 10332 29652
rect 10388 29596 10398 29652
rect 15362 29596 15372 29652
rect 15428 29596 21084 29652
rect 21140 29596 21756 29652
rect 21812 29596 22876 29652
rect 22932 29596 22942 29652
rect 23202 29596 23212 29652
rect 23268 29596 25564 29652
rect 25620 29596 25630 29652
rect 26898 29596 26908 29652
rect 26964 29596 27804 29652
rect 27860 29596 27870 29652
rect 30818 29596 30828 29652
rect 30884 29596 31836 29652
rect 31892 29596 36428 29652
rect 36484 29596 36988 29652
rect 37044 29596 37054 29652
rect 49074 29596 49084 29652
rect 49140 29596 51100 29652
rect 51156 29596 51166 29652
rect 56914 29596 56924 29652
rect 56980 29596 57372 29652
rect 57428 29596 58156 29652
rect 58212 29596 58222 29652
rect 16482 29484 16492 29540
rect 16548 29484 17276 29540
rect 17332 29484 17342 29540
rect 21522 29484 21532 29540
rect 21588 29484 22092 29540
rect 22148 29484 22158 29540
rect 22418 29484 22428 29540
rect 22484 29484 23660 29540
rect 23716 29484 23726 29540
rect 27682 29484 27692 29540
rect 27748 29484 28476 29540
rect 28532 29484 28542 29540
rect 29474 29484 29484 29540
rect 29540 29484 31164 29540
rect 31220 29484 31230 29540
rect 51538 29484 51548 29540
rect 51604 29484 53004 29540
rect 53060 29484 53070 29540
rect 29484 29428 29540 29484
rect 9986 29372 9996 29428
rect 10052 29372 12012 29428
rect 12068 29372 12078 29428
rect 16034 29372 16044 29428
rect 16100 29372 18844 29428
rect 18900 29372 18910 29428
rect 24770 29372 24780 29428
rect 24836 29372 25228 29428
rect 25284 29372 27580 29428
rect 27636 29372 29540 29428
rect 36866 29372 36876 29428
rect 36932 29372 37884 29428
rect 37940 29372 37950 29428
rect 50978 29372 50988 29428
rect 51044 29372 53228 29428
rect 53284 29372 53294 29428
rect 5058 29260 5068 29316
rect 5124 29260 14700 29316
rect 14756 29260 14766 29316
rect 14802 29036 14812 29092
rect 14868 29036 15596 29092
rect 15652 29036 15662 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 16044 28980 16100 29372
rect 20402 29260 20412 29316
rect 20468 29260 21532 29316
rect 21588 29260 21598 29316
rect 26450 29260 26460 29316
rect 26516 29260 27692 29316
rect 27748 29260 27758 29316
rect 28130 29260 28140 29316
rect 28196 29260 29708 29316
rect 29764 29260 29774 29316
rect 40226 29260 40236 29316
rect 40292 29260 41468 29316
rect 41524 29260 46508 29316
rect 46564 29260 46574 29316
rect 20738 29148 20748 29204
rect 20804 29148 21644 29204
rect 21700 29148 26908 29204
rect 26964 29148 26974 29204
rect 28690 29148 28700 29204
rect 28756 29148 35868 29204
rect 35924 29148 35934 29204
rect 41794 29148 41804 29204
rect 41860 29148 42812 29204
rect 42868 29148 42878 29204
rect 25442 29036 25452 29092
rect 25508 29036 31276 29092
rect 31332 29036 31342 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14130 28924 14140 28980
rect 14196 28924 14206 28980
rect 15092 28924 16100 28980
rect 26852 28924 34524 28980
rect 34580 28924 34590 28980
rect 38612 28924 49084 28980
rect 49140 28924 49150 28980
rect 11218 28812 11228 28868
rect 11284 28812 12012 28868
rect 12068 28812 12078 28868
rect 14140 28644 14196 28924
rect 15092 28644 15148 28924
rect 26852 28868 26908 28924
rect 25554 28812 25564 28868
rect 25620 28812 26908 28868
rect 28466 28812 28476 28868
rect 28532 28812 30604 28868
rect 30660 28812 30670 28868
rect 38612 28756 38668 28924
rect 49522 28812 49532 28868
rect 49588 28812 50652 28868
rect 50708 28812 50718 28868
rect 28812 28700 30380 28756
rect 30436 28700 30446 28756
rect 35858 28700 35868 28756
rect 35924 28700 36988 28756
rect 37044 28700 38668 28756
rect 44370 28700 44380 28756
rect 44436 28700 45276 28756
rect 45332 28700 45342 28756
rect 48514 28700 48524 28756
rect 48580 28700 49756 28756
rect 49812 28700 49822 28756
rect 51426 28700 51436 28756
rect 51492 28700 55356 28756
rect 55412 28700 56588 28756
rect 56644 28700 58044 28756
rect 58100 28700 58110 28756
rect 28812 28644 28868 28700
rect 13916 28588 14196 28644
rect 14662 28588 14700 28644
rect 14756 28588 15148 28644
rect 28354 28588 28364 28644
rect 28420 28588 28812 28644
rect 28868 28588 28878 28644
rect 29698 28588 29708 28644
rect 29764 28588 30268 28644
rect 30324 28588 31164 28644
rect 31220 28588 31230 28644
rect 31612 28588 33516 28644
rect 33572 28588 34860 28644
rect 34916 28588 34926 28644
rect 37090 28588 37100 28644
rect 37156 28588 38668 28644
rect 38724 28588 38734 28644
rect 13916 28532 13972 28588
rect 31612 28532 31668 28588
rect 12562 28476 12572 28532
rect 12628 28476 13972 28532
rect 14130 28476 14140 28532
rect 14196 28476 15148 28532
rect 15204 28476 15214 28532
rect 16146 28476 16156 28532
rect 16212 28476 17612 28532
rect 17668 28476 17678 28532
rect 30706 28476 30716 28532
rect 30772 28476 31668 28532
rect 31826 28476 31836 28532
rect 31892 28476 50428 28532
rect 52770 28476 52780 28532
rect 52836 28476 53004 28532
rect 53060 28476 53564 28532
rect 53620 28476 53630 28532
rect 55122 28476 55132 28532
rect 55188 28476 56588 28532
rect 56644 28476 56654 28532
rect 58258 28476 58268 28532
rect 58324 28476 58334 28532
rect 50372 28420 50428 28476
rect 58268 28420 58324 28476
rect 5506 28364 5516 28420
rect 5572 28364 14028 28420
rect 14084 28364 14094 28420
rect 16482 28364 16492 28420
rect 16548 28364 17724 28420
rect 17780 28364 17790 28420
rect 43362 28364 43372 28420
rect 43428 28364 44044 28420
rect 44100 28364 44110 28420
rect 50372 28364 58324 28420
rect 10994 28252 11004 28308
rect 11060 28252 14924 28308
rect 14980 28252 14990 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 34514 28140 34524 28196
rect 34580 28140 36092 28196
rect 36148 28140 37100 28196
rect 37156 28140 37166 28196
rect 37426 28140 37436 28196
rect 37492 28140 38108 28196
rect 38164 28140 38174 28196
rect 8306 28028 8316 28084
rect 8372 28028 11452 28084
rect 11508 28028 11788 28084
rect 11844 28028 12348 28084
rect 12404 28028 12684 28084
rect 12740 28028 12750 28084
rect 19170 28028 19180 28084
rect 19236 28028 19516 28084
rect 19572 28028 28700 28084
rect 28756 28028 28766 28084
rect 28914 28028 28924 28084
rect 28980 28028 29708 28084
rect 29764 28028 33852 28084
rect 33908 28028 40012 28084
rect 40068 28028 40078 28084
rect 50082 28028 50092 28084
rect 50148 28028 51660 28084
rect 51716 28028 51726 28084
rect 17602 27916 17612 27972
rect 17668 27916 18620 27972
rect 18676 27916 18686 27972
rect 4834 27804 4844 27860
rect 4900 27804 6076 27860
rect 6132 27804 7196 27860
rect 7252 27804 8092 27860
rect 8148 27804 9660 27860
rect 9716 27804 9726 27860
rect 19618 27804 19628 27860
rect 19684 27804 22876 27860
rect 22932 27804 22942 27860
rect 28924 27748 28980 28028
rect 31042 27916 31052 27972
rect 31108 27916 31388 27972
rect 31444 27916 32060 27972
rect 32116 27916 32126 27972
rect 38434 27916 38444 27972
rect 38500 27916 39004 27972
rect 39060 27916 39070 27972
rect 52658 27916 52668 27972
rect 52724 27916 55188 27972
rect 55458 27916 55468 27972
rect 55524 27916 57260 27972
rect 57316 27916 57326 27972
rect 57922 27916 57932 27972
rect 57988 27916 58156 27972
rect 58212 27916 58222 27972
rect 55132 27860 55188 27916
rect 31490 27804 31500 27860
rect 31556 27804 32508 27860
rect 32564 27804 34972 27860
rect 35028 27804 35038 27860
rect 38098 27804 38108 27860
rect 38164 27804 38668 27860
rect 38724 27804 38734 27860
rect 41122 27804 41132 27860
rect 41188 27804 41916 27860
rect 41972 27804 41982 27860
rect 50306 27804 50316 27860
rect 50372 27804 51436 27860
rect 51492 27804 51502 27860
rect 53330 27804 53340 27860
rect 53396 27804 53676 27860
rect 53732 27804 53742 27860
rect 55122 27804 55132 27860
rect 55188 27804 55198 27860
rect 7634 27692 7644 27748
rect 7700 27692 8652 27748
rect 8708 27692 9548 27748
rect 9604 27692 9614 27748
rect 9986 27692 9996 27748
rect 10052 27692 13468 27748
rect 13524 27692 14364 27748
rect 14420 27692 14430 27748
rect 23426 27692 23436 27748
rect 23492 27692 25788 27748
rect 25844 27692 28980 27748
rect 53442 27692 53452 27748
rect 53508 27692 54236 27748
rect 54292 27692 54302 27748
rect 18162 27580 18172 27636
rect 18228 27580 18956 27636
rect 19012 27580 35308 27636
rect 35364 27580 37772 27636
rect 37828 27580 39116 27636
rect 39172 27580 39182 27636
rect 56914 27580 56924 27636
rect 56980 27580 57932 27636
rect 57988 27580 57998 27636
rect 15138 27468 15148 27524
rect 15204 27468 17836 27524
rect 17892 27468 17902 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 26674 27244 26684 27300
rect 26740 27244 28140 27300
rect 28196 27244 28206 27300
rect 38210 27244 38220 27300
rect 38276 27244 38286 27300
rect 12562 27132 12572 27188
rect 12628 27132 14588 27188
rect 14644 27132 14654 27188
rect 12226 27020 12236 27076
rect 12292 27020 13580 27076
rect 13636 27020 14252 27076
rect 14308 27020 14318 27076
rect 38220 26964 38276 27244
rect 56802 27132 56812 27188
rect 56868 27132 58156 27188
rect 58212 27132 58222 27188
rect 40002 27020 40012 27076
rect 40068 27020 40908 27076
rect 40964 27020 54460 27076
rect 54516 27020 54526 27076
rect 8876 26908 10892 26964
rect 10948 26908 10958 26964
rect 13458 26908 13468 26964
rect 13524 26908 15988 26964
rect 22866 26908 22876 26964
rect 22932 26908 23996 26964
rect 24052 26908 26348 26964
rect 26404 26908 26414 26964
rect 38220 26908 38668 26964
rect 38724 26908 39676 26964
rect 39732 26908 39742 26964
rect 41906 26908 41916 26964
rect 41972 26908 42644 26964
rect 44258 26908 44268 26964
rect 44324 26908 45052 26964
rect 45108 26908 45118 26964
rect 52994 26908 53004 26964
rect 53060 26908 53452 26964
rect 53508 26908 53518 26964
rect 53676 26908 54236 26964
rect 54292 26908 54302 26964
rect 8866 26852 8876 26908
rect 8932 26852 8942 26908
rect 15932 26852 15988 26908
rect 38444 26852 38500 26908
rect 42578 26852 42588 26908
rect 42644 26852 42654 26908
rect 53676 26852 53732 26908
rect 15922 26796 15932 26852
rect 15988 26796 15998 26852
rect 24546 26796 24556 26852
rect 24612 26796 25340 26852
rect 25396 26796 26684 26852
rect 26740 26796 26750 26852
rect 26852 26796 27020 26852
rect 27076 26796 27086 26852
rect 34402 26796 34412 26852
rect 34468 26796 38500 26852
rect 43922 26796 43932 26852
rect 43988 26796 44828 26852
rect 44884 26796 44894 26852
rect 53666 26796 53676 26852
rect 53732 26796 53742 26852
rect 26852 26740 26908 26796
rect 25890 26684 25900 26740
rect 25956 26684 26908 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 14466 26572 14476 26628
rect 14532 26572 14700 26628
rect 14756 26572 14766 26628
rect 25526 26572 25564 26628
rect 25620 26572 25630 26628
rect 2258 26460 2268 26516
rect 2324 26460 22316 26516
rect 22372 26460 23324 26516
rect 23380 26460 23772 26516
rect 23828 26460 23838 26516
rect 28578 26460 28588 26516
rect 28644 26460 29596 26516
rect 29652 26460 30268 26516
rect 30324 26460 30828 26516
rect 30884 26460 31836 26516
rect 31892 26460 31902 26516
rect 37986 26460 37996 26516
rect 38052 26460 38444 26516
rect 38500 26460 39228 26516
rect 39284 26460 39294 26516
rect 56018 26460 56028 26516
rect 56084 26460 57036 26516
rect 57092 26460 57102 26516
rect 13682 26348 13692 26404
rect 13748 26348 15596 26404
rect 15652 26348 15662 26404
rect 15922 26348 15932 26404
rect 15988 26348 25116 26404
rect 25172 26348 25182 26404
rect 26002 26348 26012 26404
rect 26068 26348 27468 26404
rect 27524 26348 28812 26404
rect 28868 26348 28878 26404
rect 33282 26348 33292 26404
rect 33348 26348 39788 26404
rect 39844 26348 39854 26404
rect 41458 26348 41468 26404
rect 41524 26348 46396 26404
rect 46452 26348 46462 26404
rect 17378 26236 17388 26292
rect 17444 26236 18060 26292
rect 18116 26236 18126 26292
rect 26562 26236 26572 26292
rect 26628 26236 28252 26292
rect 28308 26236 28318 26292
rect 28578 26236 28588 26292
rect 28644 26236 29148 26292
rect 29204 26236 29372 26292
rect 29428 26236 29438 26292
rect 39442 26236 39452 26292
rect 39508 26236 40684 26292
rect 40740 26236 41132 26292
rect 41188 26236 41198 26292
rect 45826 26236 45836 26292
rect 45892 26236 58380 26292
rect 58436 26236 58446 26292
rect 8978 26124 8988 26180
rect 9044 26124 9548 26180
rect 9604 26124 11004 26180
rect 11060 26124 11070 26180
rect 16818 26124 16828 26180
rect 16884 26124 17724 26180
rect 17780 26124 17790 26180
rect 24210 26124 24220 26180
rect 24276 26124 26908 26180
rect 26964 26124 26974 26180
rect 39330 26124 39340 26180
rect 39396 26124 40124 26180
rect 40180 26124 41916 26180
rect 41972 26124 57596 26180
rect 57652 26124 57662 26180
rect 24658 26012 24668 26068
rect 24724 26012 26236 26068
rect 26292 26012 26302 26068
rect 30258 26012 30268 26068
rect 30324 26012 39116 26068
rect 39172 26012 39788 26068
rect 39844 26012 41020 26068
rect 41076 26012 41086 26068
rect 43922 26012 43932 26068
rect 43988 26012 44940 26068
rect 44996 26012 45006 26068
rect 47618 26012 47628 26068
rect 47684 26012 49084 26068
rect 49140 26012 49150 26068
rect 8866 25900 8876 25956
rect 8932 25900 9660 25956
rect 9716 25900 9726 25956
rect 15474 25900 15484 25956
rect 15540 25900 23436 25956
rect 23492 25900 23502 25956
rect 24434 25900 24444 25956
rect 24500 25900 24510 25956
rect 25554 25900 25564 25956
rect 25620 25900 26124 25956
rect 26180 25900 26190 25956
rect 26338 25900 26348 25956
rect 26404 25900 32396 25956
rect 32452 25900 32462 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 24444 25844 24500 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 24444 25788 27580 25844
rect 27636 25788 27646 25844
rect 44370 25788 44380 25844
rect 44436 25788 49980 25844
rect 50036 25788 50046 25844
rect 24098 25676 24108 25732
rect 24164 25676 24556 25732
rect 24612 25676 24622 25732
rect 25890 25676 25900 25732
rect 25956 25676 26740 25732
rect 26898 25676 26908 25732
rect 26964 25676 27692 25732
rect 27748 25676 27758 25732
rect 33842 25676 33852 25732
rect 33908 25676 34188 25732
rect 34244 25676 34972 25732
rect 35028 25676 36204 25732
rect 36260 25676 57484 25732
rect 57540 25676 57550 25732
rect 26684 25620 26740 25676
rect 9426 25564 9436 25620
rect 9492 25564 11788 25620
rect 11844 25564 11854 25620
rect 13234 25564 13244 25620
rect 13300 25564 15484 25620
rect 15540 25564 15550 25620
rect 15922 25564 15932 25620
rect 15988 25564 15998 25620
rect 26002 25564 26012 25620
rect 26068 25564 26460 25620
rect 26516 25564 26526 25620
rect 26684 25564 27132 25620
rect 27188 25564 27198 25620
rect 27794 25564 27804 25620
rect 27860 25564 28140 25620
rect 28196 25564 28588 25620
rect 28644 25564 28654 25620
rect 28914 25564 28924 25620
rect 28980 25564 35420 25620
rect 35476 25564 35486 25620
rect 37202 25564 37212 25620
rect 37268 25564 40012 25620
rect 40068 25564 40078 25620
rect 46610 25564 46620 25620
rect 46676 25564 47292 25620
rect 47348 25564 47358 25620
rect 52322 25564 52332 25620
rect 52388 25564 53564 25620
rect 53620 25564 53630 25620
rect 15932 25508 15988 25564
rect 9986 25452 9996 25508
rect 10052 25452 12236 25508
rect 12292 25452 12796 25508
rect 12852 25452 13356 25508
rect 13412 25452 13916 25508
rect 13972 25452 14700 25508
rect 14756 25452 15988 25508
rect 16258 25452 16268 25508
rect 16324 25452 17388 25508
rect 17444 25452 17454 25508
rect 17714 25452 17724 25508
rect 17780 25452 23884 25508
rect 23940 25452 23950 25508
rect 24210 25452 24220 25508
rect 24276 25452 26740 25508
rect 26684 25396 26740 25452
rect 26796 25452 27244 25508
rect 27300 25452 27310 25508
rect 27682 25452 27692 25508
rect 27748 25452 29148 25508
rect 29204 25452 30156 25508
rect 30212 25452 30222 25508
rect 32610 25452 32620 25508
rect 32676 25452 33516 25508
rect 33572 25452 34636 25508
rect 34692 25452 40124 25508
rect 40180 25452 40684 25508
rect 40740 25452 40750 25508
rect 45154 25452 45164 25508
rect 45220 25452 45948 25508
rect 46004 25452 46956 25508
rect 47012 25452 47022 25508
rect 52994 25452 53004 25508
rect 53060 25452 53452 25508
rect 53508 25452 53518 25508
rect 26796 25396 26852 25452
rect 8194 25340 8204 25396
rect 8260 25340 8988 25396
rect 9044 25340 9054 25396
rect 11554 25340 11564 25396
rect 11620 25340 14028 25396
rect 14084 25340 14094 25396
rect 23202 25340 23212 25396
rect 23268 25340 24556 25396
rect 24612 25340 26348 25396
rect 26404 25340 26414 25396
rect 26684 25340 26852 25396
rect 28018 25340 28028 25396
rect 28084 25340 32956 25396
rect 33012 25340 33022 25396
rect 35410 25340 35420 25396
rect 35476 25340 37436 25396
rect 37492 25340 37828 25396
rect 39218 25340 39228 25396
rect 39284 25340 40572 25396
rect 40628 25340 40638 25396
rect 41458 25340 41468 25396
rect 41524 25340 41916 25396
rect 41972 25340 44828 25396
rect 44884 25340 45836 25396
rect 45892 25340 45902 25396
rect 52434 25340 52444 25396
rect 52500 25340 53564 25396
rect 53620 25340 53630 25396
rect 28028 25284 28084 25340
rect 37772 25284 37828 25340
rect 21746 25228 21756 25284
rect 21812 25228 22540 25284
rect 22596 25228 22606 25284
rect 23426 25228 23436 25284
rect 23492 25228 26068 25284
rect 26226 25228 26236 25284
rect 26292 25228 28084 25284
rect 28140 25228 28924 25284
rect 28980 25228 28990 25284
rect 33170 25228 33180 25284
rect 33236 25228 33628 25284
rect 33684 25228 34076 25284
rect 34132 25228 34142 25284
rect 36082 25228 36092 25284
rect 36148 25228 37100 25284
rect 37156 25228 37166 25284
rect 37772 25228 37996 25284
rect 38052 25228 38062 25284
rect 41346 25228 41356 25284
rect 41412 25228 42476 25284
rect 42532 25228 43260 25284
rect 43316 25228 43708 25284
rect 43764 25228 44380 25284
rect 44436 25228 44446 25284
rect 50194 25228 50204 25284
rect 50260 25228 52780 25284
rect 52836 25228 52846 25284
rect 57586 25228 57596 25284
rect 57652 25228 58156 25284
rect 58212 25228 58222 25284
rect 26012 25172 26068 25228
rect 28140 25172 28196 25228
rect 14130 25116 14140 25172
rect 14196 25116 15148 25172
rect 15204 25116 18732 25172
rect 18788 25116 18798 25172
rect 20738 25116 20748 25172
rect 20804 25116 20814 25172
rect 26012 25116 28196 25172
rect 29474 25116 29484 25172
rect 29540 25116 29932 25172
rect 29988 25116 32284 25172
rect 32340 25116 42140 25172
rect 42196 25116 42206 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 20748 24948 20804 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 25442 25004 25452 25060
rect 25508 25004 26684 25060
rect 26740 25004 26750 25060
rect 16034 24892 16044 24948
rect 16100 24892 16716 24948
rect 16772 24892 17388 24948
rect 17444 24892 17454 24948
rect 18050 24892 18060 24948
rect 18116 24892 18956 24948
rect 19012 24892 19022 24948
rect 19394 24892 19404 24948
rect 19460 24892 20804 24948
rect 25526 24892 25564 24948
rect 25620 24892 25630 24948
rect 26310 24892 26348 24948
rect 26404 24892 26414 24948
rect 17602 24780 17612 24836
rect 17668 24780 18620 24836
rect 18676 24780 22764 24836
rect 22820 24780 23212 24836
rect 23268 24780 23278 24836
rect 27682 24780 27692 24836
rect 27748 24780 28924 24836
rect 28980 24780 28990 24836
rect 31892 24780 34188 24836
rect 34244 24780 41132 24836
rect 41188 24780 41198 24836
rect 52882 24780 52892 24836
rect 52948 24780 52958 24836
rect 13906 24668 13916 24724
rect 13972 24668 15820 24724
rect 15876 24668 16380 24724
rect 16436 24668 16446 24724
rect 17826 24668 17836 24724
rect 17892 24668 18172 24724
rect 18228 24668 18238 24724
rect 22642 24668 22652 24724
rect 22708 24668 23436 24724
rect 23492 24668 25228 24724
rect 25284 24668 25294 24724
rect 27458 24668 27468 24724
rect 27524 24668 28140 24724
rect 28196 24668 28206 24724
rect 31892 24612 31948 24780
rect 52892 24724 52948 24780
rect 35410 24668 35420 24724
rect 35476 24668 37884 24724
rect 37940 24668 38444 24724
rect 38500 24668 38510 24724
rect 41234 24668 41244 24724
rect 41300 24668 45164 24724
rect 45220 24668 45230 24724
rect 52892 24668 53340 24724
rect 53396 24668 53406 24724
rect 56578 24668 56588 24724
rect 56644 24668 57148 24724
rect 57204 24668 57214 24724
rect 10770 24556 10780 24612
rect 10836 24556 14028 24612
rect 14084 24556 14094 24612
rect 14242 24556 14252 24612
rect 14308 24556 15596 24612
rect 15652 24556 16268 24612
rect 16324 24556 16334 24612
rect 29138 24556 29148 24612
rect 29204 24556 29708 24612
rect 29764 24556 31948 24612
rect 35970 24556 35980 24612
rect 36036 24556 41804 24612
rect 41860 24556 42700 24612
rect 42756 24556 42766 24612
rect 43138 24556 43148 24612
rect 43204 24556 43484 24612
rect 43540 24556 45276 24612
rect 45332 24556 45724 24612
rect 45780 24556 45790 24612
rect 59200 24500 60000 24528
rect 16706 24444 16716 24500
rect 16772 24444 17836 24500
rect 17892 24444 17902 24500
rect 26338 24444 26348 24500
rect 26404 24444 27132 24500
rect 27188 24444 27198 24500
rect 31714 24444 31724 24500
rect 31780 24444 36876 24500
rect 36932 24444 36942 24500
rect 43026 24444 43036 24500
rect 43092 24444 44828 24500
rect 44884 24444 55916 24500
rect 55972 24444 55982 24500
rect 58146 24444 58156 24500
rect 58212 24444 60000 24500
rect 59200 24416 60000 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 40226 23996 40236 24052
rect 40292 23996 44604 24052
rect 44660 23996 45500 24052
rect 45556 23996 45566 24052
rect 21634 23884 21644 23940
rect 21700 23884 22204 23940
rect 22260 23884 28252 23940
rect 28308 23884 28318 23940
rect 45154 23884 45164 23940
rect 45220 23884 46060 23940
rect 46116 23884 46126 23940
rect 16258 23772 16268 23828
rect 16324 23772 17276 23828
rect 17332 23772 18956 23828
rect 19012 23772 19022 23828
rect 25116 23772 25340 23828
rect 25396 23772 25406 23828
rect 31602 23772 31612 23828
rect 31668 23772 32060 23828
rect 32116 23772 32126 23828
rect 52658 23772 52668 23828
rect 52724 23772 53732 23828
rect 25116 23716 25172 23772
rect 53676 23716 53732 23772
rect 18722 23660 18732 23716
rect 18788 23660 19852 23716
rect 19908 23660 20748 23716
rect 20804 23660 20814 23716
rect 25106 23660 25116 23716
rect 25172 23660 25182 23716
rect 29250 23660 29260 23716
rect 29316 23660 29932 23716
rect 29988 23660 29998 23716
rect 51426 23660 51436 23716
rect 51492 23660 53004 23716
rect 53060 23660 53070 23716
rect 53666 23660 53676 23716
rect 53732 23660 53742 23716
rect 22418 23548 22428 23604
rect 22484 23548 22764 23604
rect 22820 23548 24892 23604
rect 24948 23548 26908 23604
rect 26964 23548 26974 23604
rect 42690 23548 42700 23604
rect 42756 23548 43596 23604
rect 43652 23548 43662 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 21970 23436 21980 23492
rect 22036 23436 22652 23492
rect 22708 23436 23324 23492
rect 23380 23436 23390 23492
rect 24322 23436 24332 23492
rect 24388 23436 25340 23492
rect 25396 23436 25788 23492
rect 25844 23436 25854 23492
rect 26786 23436 26796 23492
rect 26852 23436 27916 23492
rect 27972 23436 27982 23492
rect 30940 23436 31948 23492
rect 32004 23436 33404 23492
rect 33460 23436 33470 23492
rect 41906 23436 41916 23492
rect 41972 23436 42476 23492
rect 42532 23436 42542 23492
rect 43362 23436 43372 23492
rect 43428 23436 44156 23492
rect 44212 23436 50428 23492
rect 23986 23324 23996 23380
rect 24052 23324 27580 23380
rect 27636 23324 30716 23380
rect 30772 23324 30782 23380
rect 30940 23268 30996 23436
rect 50372 23380 50428 23436
rect 51100 23436 57484 23492
rect 57540 23436 57550 23492
rect 51100 23380 51156 23436
rect 37874 23324 37884 23380
rect 37940 23324 41020 23380
rect 41076 23324 42924 23380
rect 42980 23324 45052 23380
rect 45108 23324 45118 23380
rect 45826 23324 45836 23380
rect 45892 23324 46844 23380
rect 46900 23324 46910 23380
rect 50372 23324 51156 23380
rect 55122 23324 55132 23380
rect 55188 23324 56700 23380
rect 56756 23324 56766 23380
rect 22754 23212 22764 23268
rect 22820 23212 30996 23268
rect 31892 23212 38108 23268
rect 38164 23212 39228 23268
rect 39284 23212 39294 23268
rect 44930 23212 44940 23268
rect 44996 23212 45612 23268
rect 45668 23212 45678 23268
rect 52210 23212 52220 23268
rect 52276 23212 53564 23268
rect 53620 23212 54124 23268
rect 54180 23212 54190 23268
rect 56578 23212 56588 23268
rect 56644 23212 57932 23268
rect 57988 23212 57998 23268
rect 31892 23156 31948 23212
rect 22978 23100 22988 23156
rect 23044 23100 24220 23156
rect 24276 23100 24286 23156
rect 28802 23100 28812 23156
rect 28868 23100 31948 23156
rect 36418 23100 36428 23156
rect 36484 23100 38444 23156
rect 38500 23100 38510 23156
rect 47954 23100 47964 23156
rect 48020 23100 50428 23156
rect 50484 23100 50494 23156
rect 50372 23044 50428 23100
rect 30706 22988 30716 23044
rect 30772 22988 33180 23044
rect 33236 22988 33246 23044
rect 46498 22988 46508 23044
rect 46564 22988 48188 23044
rect 48244 22988 48254 23044
rect 50372 22988 50764 23044
rect 50820 22988 51212 23044
rect 51268 22988 53900 23044
rect 53956 22988 54684 23044
rect 54740 22988 54750 23044
rect 33842 22876 33852 22932
rect 33908 22876 35084 22932
rect 35140 22876 35588 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 35532 22708 35588 22876
rect 20738 22652 20748 22708
rect 20804 22652 33628 22708
rect 33684 22652 33694 22708
rect 35532 22652 46172 22708
rect 46228 22652 47180 22708
rect 47236 22652 47246 22708
rect 18946 22540 18956 22596
rect 19012 22540 19740 22596
rect 19796 22540 43372 22596
rect 43428 22540 43438 22596
rect 35522 22428 35532 22484
rect 35588 22428 36428 22484
rect 36484 22428 36494 22484
rect 38770 22428 38780 22484
rect 38836 22428 40684 22484
rect 40740 22428 40750 22484
rect 42242 22428 42252 22484
rect 42308 22428 44156 22484
rect 44212 22428 44222 22484
rect 48178 22428 48188 22484
rect 48244 22428 50204 22484
rect 50260 22428 50270 22484
rect 24434 22316 24444 22372
rect 24500 22316 25900 22372
rect 25956 22316 25966 22372
rect 37174 22316 37212 22372
rect 37268 22316 37278 22372
rect 45602 22316 45612 22372
rect 45668 22316 46732 22372
rect 46788 22316 46798 22372
rect 56802 22316 56812 22372
rect 56868 22316 57372 22372
rect 57428 22316 57438 22372
rect 23874 22204 23884 22260
rect 23940 22204 24108 22260
rect 24164 22204 25228 22260
rect 25284 22204 27804 22260
rect 27860 22204 27870 22260
rect 37314 22204 37324 22260
rect 37380 22204 38444 22260
rect 38500 22204 38510 22260
rect 41458 22204 41468 22260
rect 41524 22204 42028 22260
rect 42084 22204 42094 22260
rect 43698 22204 43708 22260
rect 43764 22204 45388 22260
rect 45444 22204 45948 22260
rect 46004 22204 46014 22260
rect 54562 22204 54572 22260
rect 54628 22204 57036 22260
rect 57092 22204 57102 22260
rect 56914 22092 56924 22148
rect 56980 22092 57596 22148
rect 57652 22092 57662 22148
rect 55122 21980 55132 22036
rect 55188 21980 57148 22036
rect 57204 21980 57214 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 18610 21756 18620 21812
rect 18676 21756 19292 21812
rect 19348 21756 19964 21812
rect 20020 21756 25340 21812
rect 25396 21756 25406 21812
rect 28466 21756 28476 21812
rect 28532 21756 33628 21812
rect 33684 21756 36316 21812
rect 36372 21756 36764 21812
rect 36820 21756 36830 21812
rect 40870 21756 40908 21812
rect 40964 21756 40974 21812
rect 46946 21756 46956 21812
rect 47012 21756 49644 21812
rect 49700 21756 49710 21812
rect 18946 21644 18956 21700
rect 19012 21644 20076 21700
rect 20132 21644 20142 21700
rect 20514 21644 20524 21700
rect 20580 21644 22764 21700
rect 22820 21644 22830 21700
rect 31938 21644 31948 21700
rect 32004 21644 34524 21700
rect 34580 21644 34590 21700
rect 49746 21644 49756 21700
rect 49812 21644 50876 21700
rect 50932 21644 50942 21700
rect 21746 21532 21756 21588
rect 21812 21532 23996 21588
rect 24052 21532 24892 21588
rect 24948 21532 24958 21588
rect 34850 21532 34860 21588
rect 34916 21532 35644 21588
rect 35700 21532 35710 21588
rect 40338 21532 40348 21588
rect 40404 21532 41468 21588
rect 41524 21532 41534 21588
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 18610 20860 18620 20916
rect 18676 20860 19292 20916
rect 19348 20860 20300 20916
rect 20356 20860 29372 20916
rect 29428 20860 30156 20916
rect 30212 20860 30222 20916
rect 30930 20748 30940 20804
rect 30996 20748 33964 20804
rect 34020 20748 34030 20804
rect 15810 20636 15820 20692
rect 15876 20636 18396 20692
rect 18452 20636 18462 20692
rect 20738 20636 20748 20692
rect 20804 20636 21980 20692
rect 22036 20636 22046 20692
rect 18498 20524 18508 20580
rect 18564 20524 19628 20580
rect 19684 20524 21868 20580
rect 21924 20524 21934 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 36418 20188 36428 20244
rect 36484 20188 40460 20244
rect 40516 20188 40526 20244
rect 29026 20132 29036 20188
rect 29092 20132 29102 20188
rect 15026 20076 15036 20132
rect 15092 20076 16716 20132
rect 16772 20076 18060 20132
rect 18116 20076 19404 20132
rect 19460 20076 19470 20132
rect 26786 20076 26796 20132
rect 26852 20076 27692 20132
rect 27748 20076 29092 20132
rect 31602 20076 31612 20132
rect 31668 20076 32060 20132
rect 32116 20076 32126 20132
rect 38882 20076 38892 20132
rect 38948 20076 40348 20132
rect 40404 20076 41244 20132
rect 41300 20076 46340 20132
rect 46284 20020 46340 20076
rect 17714 19964 17724 20020
rect 17780 19964 18620 20020
rect 18676 19964 18686 20020
rect 26562 19964 26572 20020
rect 26628 19964 27244 20020
rect 27300 19964 27310 20020
rect 28242 19964 28252 20020
rect 28308 19964 30492 20020
rect 30548 19964 31052 20020
rect 31108 19964 31118 20020
rect 31378 19964 31388 20020
rect 31444 19964 31836 20020
rect 31892 19964 31902 20020
rect 41458 19964 41468 20020
rect 41524 19964 42140 20020
rect 42196 19964 42206 20020
rect 46274 19964 46284 20020
rect 46340 19964 46844 20020
rect 46900 19964 46910 20020
rect 47282 19964 47292 20020
rect 47348 19964 47964 20020
rect 48020 19964 48030 20020
rect 37762 19852 37772 19908
rect 37828 19852 38668 19908
rect 38724 19852 38734 19908
rect 41010 19852 41020 19908
rect 41076 19852 42588 19908
rect 42644 19852 42654 19908
rect 44370 19852 44380 19908
rect 44436 19852 45164 19908
rect 45220 19852 45230 19908
rect 46722 19852 46732 19908
rect 46788 19852 47852 19908
rect 47908 19852 47918 19908
rect 38770 19740 38780 19796
rect 38836 19740 40908 19796
rect 40964 19740 41916 19796
rect 41972 19740 41982 19796
rect 46946 19740 46956 19796
rect 47012 19740 47516 19796
rect 47572 19740 47582 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 23202 19404 23212 19460
rect 23268 19404 33740 19460
rect 33796 19404 33806 19460
rect 34178 19404 34188 19460
rect 34244 19404 36988 19460
rect 37044 19404 42364 19460
rect 42420 19404 42430 19460
rect 46162 19404 46172 19460
rect 46228 19404 47628 19460
rect 47684 19404 47694 19460
rect 19282 19292 19292 19348
rect 19348 19292 26236 19348
rect 26292 19292 26796 19348
rect 26852 19292 26862 19348
rect 34514 19292 34524 19348
rect 34580 19292 38892 19348
rect 38948 19292 38958 19348
rect 39106 19292 39116 19348
rect 39172 19292 39788 19348
rect 39844 19292 44380 19348
rect 44436 19292 44446 19348
rect 47730 19292 47740 19348
rect 47796 19292 50764 19348
rect 50820 19292 50830 19348
rect 23202 19180 23212 19236
rect 23268 19180 23660 19236
rect 23716 19180 24332 19236
rect 24388 19180 25004 19236
rect 25060 19180 25070 19236
rect 37090 19180 37100 19236
rect 37156 19180 38780 19236
rect 38836 19180 38846 19236
rect 47170 19180 47180 19236
rect 47236 19180 50316 19236
rect 50372 19180 54908 19236
rect 54964 19180 54974 19236
rect 29932 19068 31500 19124
rect 31556 19068 31948 19124
rect 32004 19068 32014 19124
rect 34178 19068 34188 19124
rect 34244 19068 35420 19124
rect 35476 19068 35486 19124
rect 17266 18956 17276 19012
rect 17332 18956 18508 19012
rect 18564 18956 18574 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 29932 18788 29988 19068
rect 30258 18956 30268 19012
rect 30324 18956 30716 19012
rect 30772 18956 30782 19012
rect 33618 18956 33628 19012
rect 33684 18956 34636 19012
rect 34692 18956 34702 19012
rect 34962 18956 34972 19012
rect 35028 18956 38332 19012
rect 38388 18956 38398 19012
rect 42018 18956 42028 19012
rect 42084 18956 44716 19012
rect 44772 18956 44782 19012
rect 50754 18956 50764 19012
rect 50820 18956 52108 19012
rect 52164 18956 53788 19012
rect 53844 18956 53854 19012
rect 38332 18900 38388 18956
rect 36082 18844 36092 18900
rect 36148 18844 37884 18900
rect 37940 18844 37950 18900
rect 38332 18844 40236 18900
rect 40292 18844 40302 18900
rect 37884 18788 37940 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 28476 18732 29932 18788
rect 29988 18732 29998 18788
rect 31938 18732 31948 18788
rect 32004 18732 33068 18788
rect 33124 18732 37828 18788
rect 37884 18732 39564 18788
rect 39620 18732 41244 18788
rect 41300 18732 41310 18788
rect 50306 18732 50316 18788
rect 28476 18676 28532 18732
rect 37772 18676 37828 18732
rect 19058 18620 19068 18676
rect 19124 18620 19292 18676
rect 19348 18620 19358 18676
rect 27458 18620 27468 18676
rect 27524 18620 28476 18676
rect 28532 18620 28542 18676
rect 29362 18620 29372 18676
rect 29428 18620 30380 18676
rect 30436 18620 33852 18676
rect 33908 18620 35084 18676
rect 35140 18620 35150 18676
rect 37772 18620 42364 18676
rect 42420 18620 43148 18676
rect 43204 18620 45276 18676
rect 45332 18620 45948 18676
rect 46004 18620 46014 18676
rect 50372 18620 50428 18788
rect 50484 18620 50494 18676
rect 24210 18508 24220 18564
rect 24276 18508 33628 18564
rect 33684 18508 33694 18564
rect 35970 18508 35980 18564
rect 36036 18508 37100 18564
rect 37156 18508 37166 18564
rect 44706 18508 44716 18564
rect 44772 18508 46732 18564
rect 46788 18508 46798 18564
rect 24220 18452 24276 18508
rect 15138 18396 15148 18452
rect 15204 18396 18060 18452
rect 18116 18396 18126 18452
rect 18274 18396 18284 18452
rect 18340 18396 19068 18452
rect 19124 18396 19134 18452
rect 23090 18396 23100 18452
rect 23156 18396 24276 18452
rect 27122 18396 27132 18452
rect 27188 18396 28588 18452
rect 28644 18396 28654 18452
rect 32162 18396 32172 18452
rect 32228 18396 33516 18452
rect 33572 18396 33582 18452
rect 34738 18396 34748 18452
rect 34804 18396 35868 18452
rect 35924 18396 35934 18452
rect 41346 18396 41356 18452
rect 41412 18396 42588 18452
rect 42644 18396 42654 18452
rect 44482 18396 44492 18452
rect 44548 18396 50428 18452
rect 51538 18396 51548 18452
rect 51604 18396 52220 18452
rect 52276 18396 52286 18452
rect 50372 18340 50428 18396
rect 22530 18284 22540 18340
rect 22596 18284 22606 18340
rect 23762 18284 23772 18340
rect 23828 18284 23838 18340
rect 24434 18284 24444 18340
rect 24500 18284 28924 18340
rect 28980 18284 28990 18340
rect 31378 18284 31388 18340
rect 31444 18284 37212 18340
rect 37268 18284 37278 18340
rect 40226 18284 40236 18340
rect 40292 18284 41804 18340
rect 41860 18284 41870 18340
rect 50372 18284 52444 18340
rect 52500 18284 52668 18340
rect 52724 18284 52734 18340
rect 53218 18284 53228 18340
rect 53284 18284 54460 18340
rect 54516 18284 54526 18340
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 22540 17780 22596 18284
rect 23772 18116 23828 18284
rect 28924 18228 28980 18284
rect 28924 18172 32284 18228
rect 32340 18172 32350 18228
rect 34972 18172 42364 18228
rect 42420 18172 43596 18228
rect 43652 18172 43932 18228
rect 43988 18172 43998 18228
rect 52322 18172 52332 18228
rect 52388 18172 53564 18228
rect 53620 18172 53630 18228
rect 54562 18172 54572 18228
rect 54628 18172 56476 18228
rect 56532 18172 56542 18228
rect 34972 18116 35028 18172
rect 23772 18060 25004 18116
rect 25060 18060 35028 18116
rect 37090 18060 37100 18116
rect 37156 18060 40572 18116
rect 40628 18060 40638 18116
rect 51286 18060 51324 18116
rect 51380 18060 51390 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 40002 17948 40012 18004
rect 40068 17948 57820 18004
rect 57876 17948 57886 18004
rect 35522 17836 35532 17892
rect 35588 17836 37772 17892
rect 37828 17836 38556 17892
rect 38612 17836 38622 17892
rect 41458 17836 41468 17892
rect 41524 17836 44268 17892
rect 44324 17836 45276 17892
rect 45332 17836 45342 17892
rect 52070 17836 52108 17892
rect 52164 17836 52174 17892
rect 52322 17836 52332 17892
rect 52388 17836 52780 17892
rect 52836 17836 54124 17892
rect 54180 17836 54190 17892
rect 21634 17724 21644 17780
rect 21700 17724 22316 17780
rect 22372 17724 30940 17780
rect 30996 17724 31388 17780
rect 31444 17724 31454 17780
rect 39778 17724 39788 17780
rect 39844 17724 40684 17780
rect 40740 17724 40750 17780
rect 50978 17724 50988 17780
rect 51044 17724 53340 17780
rect 53396 17724 54348 17780
rect 54404 17724 54414 17780
rect 19842 17612 19852 17668
rect 19908 17612 24444 17668
rect 24500 17612 24510 17668
rect 28802 17612 28812 17668
rect 28868 17612 30492 17668
rect 30548 17612 30558 17668
rect 31154 17612 31164 17668
rect 31220 17612 31612 17668
rect 31668 17612 31678 17668
rect 40562 17612 40572 17668
rect 40628 17612 40908 17668
rect 40964 17612 40974 17668
rect 41682 17612 41692 17668
rect 41748 17612 44940 17668
rect 44996 17612 45006 17668
rect 47170 17612 47180 17668
rect 47236 17612 49980 17668
rect 50036 17612 50652 17668
rect 50708 17612 50718 17668
rect 50866 17612 50876 17668
rect 50932 17612 50942 17668
rect 54898 17612 54908 17668
rect 54964 17612 57148 17668
rect 57204 17612 57214 17668
rect 50876 17556 50932 17612
rect 59200 17556 60000 17584
rect 18946 17500 18956 17556
rect 19012 17500 22764 17556
rect 22820 17500 22830 17556
rect 50876 17500 53564 17556
rect 53620 17500 53630 17556
rect 58146 17500 58156 17556
rect 58212 17500 60000 17556
rect 53564 17444 53620 17500
rect 59200 17472 60000 17500
rect 14690 17388 14700 17444
rect 14756 17388 17500 17444
rect 17556 17388 17566 17444
rect 18274 17388 18284 17444
rect 18340 17388 19180 17444
rect 19236 17388 21196 17444
rect 21252 17388 21262 17444
rect 25330 17388 25340 17444
rect 25396 17388 27916 17444
rect 27972 17388 28364 17444
rect 28420 17388 29708 17444
rect 29764 17388 30828 17444
rect 30884 17388 33180 17444
rect 33236 17388 33246 17444
rect 35074 17388 35084 17444
rect 35140 17388 35980 17444
rect 36036 17388 36046 17444
rect 44482 17388 44492 17444
rect 44548 17388 46620 17444
rect 46676 17388 47404 17444
rect 47460 17388 47470 17444
rect 52434 17388 52444 17444
rect 52500 17388 52780 17444
rect 52836 17388 53116 17444
rect 53172 17388 53182 17444
rect 53564 17388 53788 17444
rect 53844 17388 53854 17444
rect 17378 17276 17388 17332
rect 17444 17276 18396 17332
rect 18452 17276 18462 17332
rect 53330 17276 53340 17332
rect 53396 17276 55132 17332
rect 55188 17276 55198 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 17714 17164 17724 17220
rect 17780 17164 18284 17220
rect 18340 17164 19684 17220
rect 28690 17164 28700 17220
rect 28756 17164 31500 17220
rect 31556 17164 31566 17220
rect 19628 17108 19684 17164
rect 16818 17052 16828 17108
rect 16884 17052 18060 17108
rect 18116 17052 18508 17108
rect 18564 17052 18574 17108
rect 19628 17052 27580 17108
rect 27636 17052 28140 17108
rect 28196 17052 35420 17108
rect 35476 17052 35486 17108
rect 51202 17052 51212 17108
rect 51268 17052 51660 17108
rect 51716 17052 51726 17108
rect 51986 17052 51996 17108
rect 52052 17052 52668 17108
rect 52724 17052 52734 17108
rect 16594 16940 16604 16996
rect 16660 16940 18620 16996
rect 18676 16940 18686 16996
rect 16828 16828 17612 16884
rect 17668 16828 19628 16884
rect 19684 16828 19694 16884
rect 49298 16828 49308 16884
rect 49364 16828 50316 16884
rect 50372 16828 50382 16884
rect 51650 16828 51660 16884
rect 51716 16828 52892 16884
rect 52948 16828 52958 16884
rect 53778 16828 53788 16884
rect 53844 16828 55020 16884
rect 55076 16828 55086 16884
rect 16828 16772 16884 16828
rect 15810 16716 15820 16772
rect 15876 16716 16884 16772
rect 28242 16716 28252 16772
rect 28308 16716 28812 16772
rect 28868 16716 28878 16772
rect 31892 16716 32508 16772
rect 32564 16716 34188 16772
rect 34244 16716 34254 16772
rect 44146 16716 44156 16772
rect 44212 16716 49084 16772
rect 49140 16716 49150 16772
rect 51314 16716 51324 16772
rect 51380 16716 52220 16772
rect 52276 16716 53340 16772
rect 53396 16716 53406 16772
rect 55234 16716 55244 16772
rect 55300 16716 57372 16772
rect 57428 16716 57438 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 31892 16324 31948 16716
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 10994 16268 11004 16324
rect 11060 16268 26908 16324
rect 31714 16268 31724 16324
rect 31780 16268 31948 16324
rect 38322 16268 38332 16324
rect 38388 16268 41020 16324
rect 41076 16268 41086 16324
rect 18722 16156 18732 16212
rect 18788 16156 19404 16212
rect 19460 16156 19470 16212
rect 20402 16156 20412 16212
rect 20468 16156 21868 16212
rect 21924 16156 22428 16212
rect 22484 16156 22764 16212
rect 22820 16156 22830 16212
rect 26852 16100 26908 16268
rect 32162 16156 32172 16212
rect 32228 16156 33628 16212
rect 33684 16156 33694 16212
rect 35522 16156 35532 16212
rect 35588 16156 36092 16212
rect 36148 16156 36158 16212
rect 32172 16100 32228 16156
rect 14018 16044 14028 16100
rect 14084 16044 15820 16100
rect 15876 16044 15886 16100
rect 26852 16044 32228 16100
rect 19282 15932 19292 15988
rect 19348 15932 27468 15988
rect 27524 15932 28140 15988
rect 28196 15932 28206 15988
rect 28354 15932 28364 15988
rect 28420 15932 29372 15988
rect 29428 15932 29438 15988
rect 34290 15932 34300 15988
rect 34356 15932 37772 15988
rect 37828 15932 37838 15988
rect 40674 15932 40684 15988
rect 40740 15932 47852 15988
rect 47908 15932 47918 15988
rect 50372 15932 50540 15988
rect 50596 15932 50606 15988
rect 28140 15876 28196 15932
rect 50372 15876 50428 15932
rect 22978 15820 22988 15876
rect 23044 15820 23660 15876
rect 23716 15820 23726 15876
rect 28140 15820 31724 15876
rect 31780 15820 31790 15876
rect 32722 15820 32732 15876
rect 32788 15820 33180 15876
rect 33236 15820 37604 15876
rect 39666 15820 39676 15876
rect 39732 15820 41132 15876
rect 41188 15820 45052 15876
rect 45108 15820 45388 15876
rect 45444 15820 45454 15876
rect 45714 15820 45724 15876
rect 45780 15820 47180 15876
rect 47236 15820 47246 15876
rect 47730 15820 47740 15876
rect 47796 15820 50428 15876
rect 37548 15764 37604 15820
rect 24770 15708 24780 15764
rect 24836 15708 25228 15764
rect 25284 15708 35532 15764
rect 35588 15708 35598 15764
rect 37538 15708 37548 15764
rect 37604 15708 40908 15764
rect 40964 15708 40974 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 47282 15484 47292 15540
rect 47348 15484 48972 15540
rect 49028 15484 50428 15540
rect 51650 15484 51660 15540
rect 51716 15484 52332 15540
rect 52388 15484 52398 15540
rect 34626 15372 34636 15428
rect 34692 15372 35308 15428
rect 35364 15372 35374 15428
rect 38098 15372 38108 15428
rect 38164 15372 39228 15428
rect 39284 15372 39294 15428
rect 47170 15372 47180 15428
rect 47236 15372 48860 15428
rect 48916 15372 49420 15428
rect 49476 15372 49980 15428
rect 50036 15372 50046 15428
rect 50372 15316 50428 15484
rect 38546 15260 38556 15316
rect 38612 15260 39676 15316
rect 39732 15260 39742 15316
rect 41010 15260 41020 15316
rect 41076 15260 41916 15316
rect 41972 15260 41982 15316
rect 45714 15260 45724 15316
rect 45780 15260 46844 15316
rect 46900 15260 46910 15316
rect 50372 15260 52108 15316
rect 52164 15260 52174 15316
rect 31714 15148 31724 15204
rect 31780 15148 32508 15204
rect 32564 15148 33852 15204
rect 33908 15148 33918 15204
rect 43652 15148 44716 15204
rect 44772 15148 46620 15204
rect 46676 15148 46686 15204
rect 50194 15148 50204 15204
rect 50260 15148 51436 15204
rect 51492 15148 52556 15204
rect 52612 15148 52622 15204
rect 43652 15092 43708 15148
rect 32050 15036 32060 15092
rect 32116 15036 33404 15092
rect 33460 15036 33470 15092
rect 41682 15036 41692 15092
rect 41748 15036 42812 15092
rect 42868 15036 43708 15092
rect 50642 15036 50652 15092
rect 50708 15036 53564 15092
rect 53620 15036 53630 15092
rect 54226 15036 54236 15092
rect 54292 15036 56476 15092
rect 56532 15036 56542 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 22642 14812 22652 14868
rect 22708 14812 26796 14868
rect 26852 14644 26908 14868
rect 38612 14812 51212 14868
rect 51268 14812 51884 14868
rect 51940 14812 51950 14868
rect 38612 14756 38668 14812
rect 28466 14700 28476 14756
rect 28532 14700 38332 14756
rect 38388 14700 38668 14756
rect 40002 14700 40012 14756
rect 40068 14700 43036 14756
rect 43092 14700 43102 14756
rect 49298 14700 49308 14756
rect 49364 14700 50540 14756
rect 50596 14700 50606 14756
rect 17266 14588 17276 14644
rect 17332 14588 18284 14644
rect 18340 14588 18350 14644
rect 23202 14588 23212 14644
rect 23268 14588 26460 14644
rect 26516 14588 26526 14644
rect 26852 14588 27580 14644
rect 27636 14588 32732 14644
rect 32788 14588 32798 14644
rect 41458 14588 41468 14644
rect 41524 14588 42588 14644
rect 42644 14588 42654 14644
rect 50418 14588 50428 14644
rect 50484 14588 50764 14644
rect 50820 14588 52780 14644
rect 52836 14588 52846 14644
rect 53554 14588 53564 14644
rect 53620 14588 54348 14644
rect 54404 14588 54414 14644
rect 18498 14476 18508 14532
rect 18564 14476 19068 14532
rect 19124 14476 22428 14532
rect 22484 14476 22494 14532
rect 41906 14476 41916 14532
rect 41972 14476 43036 14532
rect 43092 14476 43708 14532
rect 43652 14420 43708 14476
rect 47628 14476 48076 14532
rect 48132 14476 50204 14532
rect 50260 14476 51212 14532
rect 51268 14476 51278 14532
rect 52098 14476 52108 14532
rect 52164 14476 53004 14532
rect 53060 14476 53070 14532
rect 47628 14420 47684 14476
rect 39554 14364 39564 14420
rect 39620 14364 40908 14420
rect 40964 14364 40974 14420
rect 43652 14364 44044 14420
rect 44100 14364 44716 14420
rect 44772 14364 44782 14420
rect 47618 14364 47628 14420
rect 47684 14364 47694 14420
rect 48290 14364 48300 14420
rect 48356 14364 51604 14420
rect 51762 14364 51772 14420
rect 51828 14364 53340 14420
rect 53396 14364 53406 14420
rect 51548 14308 51604 14364
rect 24322 14252 24332 14308
rect 24388 14252 27132 14308
rect 27188 14252 28140 14308
rect 28196 14252 28206 14308
rect 33730 14252 33740 14308
rect 33796 14252 41132 14308
rect 41188 14252 41198 14308
rect 41458 14252 41468 14308
rect 41524 14252 42700 14308
rect 42756 14252 42766 14308
rect 50530 14252 50540 14308
rect 50596 14252 50988 14308
rect 51044 14252 51054 14308
rect 51538 14252 51548 14308
rect 51604 14252 53116 14308
rect 53172 14252 53182 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 14690 13916 14700 13972
rect 14756 13916 20748 13972
rect 20804 13916 20814 13972
rect 34178 13916 34188 13972
rect 34244 13916 34524 13972
rect 34580 13916 34590 13972
rect 39106 13916 39116 13972
rect 39172 13916 39182 13972
rect 41906 13916 41916 13972
rect 41972 13916 43260 13972
rect 43316 13916 43326 13972
rect 44482 13916 44492 13972
rect 44548 13916 44558 13972
rect 39116 13860 39172 13916
rect 44492 13860 44548 13916
rect 16818 13804 16828 13860
rect 16884 13804 18508 13860
rect 18564 13804 18732 13860
rect 18788 13804 19852 13860
rect 19908 13804 19918 13860
rect 21074 13804 21084 13860
rect 21140 13804 22092 13860
rect 22148 13804 22158 13860
rect 22642 13804 22652 13860
rect 22708 13804 23324 13860
rect 23380 13804 23390 13860
rect 28914 13804 28924 13860
rect 28980 13804 30044 13860
rect 30100 13804 35588 13860
rect 35746 13804 35756 13860
rect 35812 13804 37212 13860
rect 37268 13804 37548 13860
rect 37604 13804 37884 13860
rect 37940 13804 38444 13860
rect 38500 13804 39172 13860
rect 44156 13804 44548 13860
rect 44930 13804 44940 13860
rect 44996 13804 47516 13860
rect 47572 13804 47582 13860
rect 18834 13692 18844 13748
rect 18900 13692 21756 13748
rect 21812 13692 21822 13748
rect 22194 13692 22204 13748
rect 22260 13692 23100 13748
rect 23156 13692 23166 13748
rect 32162 13692 32172 13748
rect 32228 13692 33068 13748
rect 33124 13692 33740 13748
rect 33796 13692 33806 13748
rect 35532 13636 35588 13804
rect 44156 13748 44212 13804
rect 44146 13692 44156 13748
rect 44212 13692 44222 13748
rect 47394 13692 47404 13748
rect 47460 13692 50204 13748
rect 50260 13692 50270 13748
rect 51874 13692 51884 13748
rect 51940 13692 52668 13748
rect 52724 13692 52734 13748
rect 55346 13692 55356 13748
rect 55412 13692 56028 13748
rect 56084 13692 56700 13748
rect 56756 13692 56766 13748
rect 14018 13580 14028 13636
rect 14084 13580 17500 13636
rect 17556 13580 23212 13636
rect 23268 13580 23278 13636
rect 29922 13580 29932 13636
rect 29988 13580 30492 13636
rect 30548 13580 31836 13636
rect 31892 13580 31902 13636
rect 35522 13580 35532 13636
rect 35588 13580 35598 13636
rect 42130 13580 42140 13636
rect 42196 13580 43708 13636
rect 43764 13580 50316 13636
rect 50372 13580 50382 13636
rect 52770 13580 52780 13636
rect 52836 13580 55244 13636
rect 55300 13580 55310 13636
rect 18946 13468 18956 13524
rect 19012 13468 19404 13524
rect 19460 13468 19470 13524
rect 20402 13468 20412 13524
rect 20468 13468 21196 13524
rect 21252 13468 23548 13524
rect 23604 13468 23614 13524
rect 24658 13468 24668 13524
rect 24724 13468 35308 13524
rect 35364 13468 35374 13524
rect 39106 13468 39116 13524
rect 39172 13468 40012 13524
rect 40068 13468 40078 13524
rect 39116 13412 39172 13468
rect 19842 13356 19852 13412
rect 19908 13356 20300 13412
rect 20356 13356 20366 13412
rect 33394 13356 33404 13412
rect 33460 13356 33796 13412
rect 34066 13356 34076 13412
rect 34132 13356 34972 13412
rect 35028 13356 35038 13412
rect 36428 13356 39172 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 33740 13300 33796 13356
rect 33740 13244 34020 13300
rect 33964 13188 34020 13244
rect 34972 13188 35028 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 17826 13132 17836 13188
rect 17892 13132 18284 13188
rect 18340 13132 20076 13188
rect 20132 13132 20142 13188
rect 23762 13132 23772 13188
rect 23828 13132 24556 13188
rect 24612 13132 33236 13188
rect 33954 13132 33964 13188
rect 34020 13132 34748 13188
rect 34804 13132 34814 13188
rect 34972 13132 35644 13188
rect 35700 13132 35710 13188
rect 33180 13076 33236 13132
rect 36428 13076 36484 13356
rect 20178 13020 20188 13076
rect 20244 13020 20860 13076
rect 20916 13020 28476 13076
rect 28532 13020 28542 13076
rect 33180 13020 34972 13076
rect 35028 13020 36428 13076
rect 36484 13020 36494 13076
rect 42914 13020 42924 13076
rect 42980 13020 49756 13076
rect 49812 13020 49822 13076
rect 22530 12908 22540 12964
rect 22596 12908 24220 12964
rect 24276 12908 24286 12964
rect 24770 12908 24780 12964
rect 24836 12908 25228 12964
rect 25284 12908 25294 12964
rect 29474 12908 29484 12964
rect 29540 12908 29932 12964
rect 29988 12908 29998 12964
rect 32050 12908 32060 12964
rect 32116 12908 32620 12964
rect 32676 12908 32686 12964
rect 32946 12908 32956 12964
rect 33012 12908 38780 12964
rect 38836 12908 39676 12964
rect 39732 12908 52892 12964
rect 52948 12908 52958 12964
rect 17938 12796 17948 12852
rect 18004 12796 18732 12852
rect 18788 12796 19180 12852
rect 19236 12796 19246 12852
rect 21634 12796 21644 12852
rect 21700 12796 22428 12852
rect 22484 12796 32172 12852
rect 32228 12796 32238 12852
rect 32386 12796 32396 12852
rect 32452 12796 33292 12852
rect 33348 12796 33358 12852
rect 34514 12796 34524 12852
rect 34580 12796 35420 12852
rect 35476 12796 35486 12852
rect 35970 12796 35980 12852
rect 36036 12796 37100 12852
rect 37156 12796 37166 12852
rect 41122 12796 41132 12852
rect 41188 12796 42028 12852
rect 42084 12796 42588 12852
rect 42644 12796 42654 12852
rect 44034 12796 44044 12852
rect 44100 12796 45276 12852
rect 45332 12796 47852 12852
rect 47908 12796 47918 12852
rect 17826 12684 17836 12740
rect 17892 12684 19404 12740
rect 19460 12684 19470 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 23324 12516 23380 12796
rect 35980 12740 36036 12796
rect 25218 12684 25228 12740
rect 25284 12684 26684 12740
rect 26740 12684 27468 12740
rect 27524 12684 36036 12740
rect 44706 12684 44716 12740
rect 44772 12684 45612 12740
rect 45668 12684 45678 12740
rect 31602 12572 31612 12628
rect 31668 12572 32508 12628
rect 32564 12572 32574 12628
rect 45490 12572 45500 12628
rect 45556 12572 47516 12628
rect 47572 12572 50204 12628
rect 50260 12572 50270 12628
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 23314 12460 23324 12516
rect 23380 12460 23390 12516
rect 43652 12460 49532 12516
rect 49588 12460 49598 12516
rect 40226 12348 40236 12404
rect 40292 12348 40302 12404
rect 40236 12292 40292 12348
rect 43652 12292 43708 12460
rect 49746 12348 49756 12404
rect 49812 12348 50652 12404
rect 50708 12348 51436 12404
rect 51492 12348 51502 12404
rect 39116 12236 42364 12292
rect 42420 12236 43708 12292
rect 50306 12236 50316 12292
rect 50372 12236 52220 12292
rect 52276 12236 52668 12292
rect 52724 12236 52734 12292
rect 39116 12180 39172 12236
rect 26852 12124 30156 12180
rect 30212 12124 32956 12180
rect 33012 12124 33022 12180
rect 39106 12124 39116 12180
rect 39172 12124 39182 12180
rect 26852 11956 26908 12124
rect 27010 12012 27020 12068
rect 27076 12012 27468 12068
rect 27524 12012 27534 12068
rect 27794 12012 27804 12068
rect 27860 12012 28252 12068
rect 28308 12012 34300 12068
rect 34356 12012 35084 12068
rect 35140 12012 38668 12068
rect 40226 12012 40236 12068
rect 40292 12012 42140 12068
rect 42196 12012 42206 12068
rect 38612 11956 38668 12012
rect 18274 11900 18284 11956
rect 18340 11900 21196 11956
rect 21252 11900 26908 11956
rect 34626 11900 34636 11956
rect 34692 11900 37660 11956
rect 37716 11900 38108 11956
rect 38164 11900 38174 11956
rect 38612 11900 38780 11956
rect 38836 11900 41692 11956
rect 41748 11900 50988 11956
rect 51044 11900 51660 11956
rect 51716 11900 51726 11956
rect 30594 11788 30604 11844
rect 30660 11788 31500 11844
rect 31556 11788 31566 11844
rect 0 11732 800 11760
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 0 11676 2996 11732
rect 5842 11676 5852 11732
rect 5908 11676 5918 11732
rect 18946 11676 18956 11732
rect 19012 11676 21308 11732
rect 21364 11676 21374 11732
rect 22642 11676 22652 11732
rect 22708 11676 31836 11732
rect 31892 11676 33516 11732
rect 33572 11676 33582 11732
rect 36194 11676 36204 11732
rect 36260 11676 57260 11732
rect 57316 11676 57326 11732
rect 0 11648 800 11676
rect 2940 11620 2996 11676
rect 5852 11620 5908 11676
rect 2940 11564 5908 11620
rect 28242 11564 28252 11620
rect 28308 11564 29708 11620
rect 29764 11564 37884 11620
rect 37940 11564 38668 11620
rect 38724 11564 38734 11620
rect 46946 11564 46956 11620
rect 47012 11564 48412 11620
rect 48468 11564 48478 11620
rect 49858 11564 49868 11620
rect 49924 11564 51100 11620
rect 51156 11564 51324 11620
rect 51380 11564 51390 11620
rect 55346 11564 55356 11620
rect 55412 11508 55468 11620
rect 17266 11452 17276 11508
rect 17332 11452 18284 11508
rect 18340 11452 18732 11508
rect 18788 11452 18798 11508
rect 27122 11452 27132 11508
rect 27188 11452 27468 11508
rect 27524 11452 29260 11508
rect 29316 11452 30156 11508
rect 30212 11452 30222 11508
rect 35522 11452 35532 11508
rect 35588 11452 38332 11508
rect 38388 11452 39452 11508
rect 39508 11452 39518 11508
rect 41010 11452 41020 11508
rect 41076 11452 43036 11508
rect 43092 11452 43102 11508
rect 47842 11452 47852 11508
rect 47908 11452 48860 11508
rect 48916 11452 48926 11508
rect 49634 11452 49644 11508
rect 49700 11452 50092 11508
rect 50148 11452 55580 11508
rect 55636 11452 56028 11508
rect 56084 11452 56094 11508
rect 17714 11340 17724 11396
rect 17780 11340 18844 11396
rect 18900 11340 18910 11396
rect 33506 11340 33516 11396
rect 33572 11340 42028 11396
rect 42084 11340 42094 11396
rect 52098 11340 52108 11396
rect 52164 11340 52780 11396
rect 52836 11340 52846 11396
rect 18946 11228 18956 11284
rect 19012 11228 20244 11284
rect 21970 11228 21980 11284
rect 22036 11228 32060 11284
rect 32116 11228 33964 11284
rect 34020 11228 34030 11284
rect 51762 11228 51772 11284
rect 51828 11228 54796 11284
rect 54852 11228 54862 11284
rect 20188 11172 20244 11228
rect 15922 11116 15932 11172
rect 15988 11116 18844 11172
rect 18900 11116 18910 11172
rect 20178 11116 20188 11172
rect 20244 11116 42252 11172
rect 42308 11116 42318 11172
rect 33282 11004 33292 11060
rect 33348 11004 35532 11060
rect 35588 11004 35598 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 31154 10892 31164 10948
rect 31220 10892 31724 10948
rect 31780 10892 46956 10948
rect 47012 10892 47022 10948
rect 18946 10780 18956 10836
rect 19012 10780 19292 10836
rect 19348 10780 19358 10836
rect 38994 10780 39004 10836
rect 39060 10780 40236 10836
rect 40292 10780 41692 10836
rect 41748 10780 41758 10836
rect 42130 10780 42140 10836
rect 42196 10780 51996 10836
rect 52052 10780 52062 10836
rect 41692 10724 41748 10780
rect 18386 10668 18396 10724
rect 18452 10668 21532 10724
rect 21588 10668 21598 10724
rect 41692 10668 42924 10724
rect 42980 10668 42990 10724
rect 43922 10668 43932 10724
rect 43988 10668 44604 10724
rect 44660 10668 44670 10724
rect 59200 10612 60000 10640
rect 19142 10556 19180 10612
rect 19236 10556 19246 10612
rect 24546 10556 24556 10612
rect 24612 10556 25340 10612
rect 25396 10556 27132 10612
rect 27188 10556 27198 10612
rect 42242 10556 42252 10612
rect 42308 10556 42318 10612
rect 43138 10556 43148 10612
rect 43204 10556 44380 10612
rect 44436 10556 44446 10612
rect 58146 10556 58156 10612
rect 58212 10556 60000 10612
rect 42252 10500 42308 10556
rect 59200 10528 60000 10556
rect 42252 10444 50652 10500
rect 50708 10444 50718 10500
rect 21634 10332 21644 10388
rect 21700 10332 22764 10388
rect 22820 10332 25340 10388
rect 25396 10332 25406 10388
rect 40450 10332 40460 10388
rect 40516 10332 49532 10388
rect 49588 10332 49598 10388
rect 27010 10220 27020 10276
rect 27076 10220 32900 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 14354 10108 14364 10164
rect 14420 10108 17500 10164
rect 17556 10108 17724 10164
rect 17780 10108 17790 10164
rect 18844 10108 19964 10164
rect 20020 10108 20030 10164
rect 24658 10108 24668 10164
rect 24724 10108 27580 10164
rect 27636 10108 27646 10164
rect 18844 10052 18900 10108
rect 32844 10052 32900 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 42914 10108 42924 10164
rect 42980 10108 46844 10164
rect 46900 10108 46910 10164
rect 52098 10108 52108 10164
rect 52164 10108 53228 10164
rect 53284 10108 53294 10164
rect 18834 9996 18844 10052
rect 18900 9996 18910 10052
rect 32834 9996 32844 10052
rect 32900 9996 38668 10052
rect 50194 9996 50204 10052
rect 50260 9996 51212 10052
rect 51268 9996 51278 10052
rect 38612 9940 38668 9996
rect 15922 9884 15932 9940
rect 15988 9884 18620 9940
rect 18676 9884 18686 9940
rect 21746 9884 21756 9940
rect 21812 9884 22204 9940
rect 22260 9884 25004 9940
rect 25060 9884 25070 9940
rect 27458 9884 27468 9940
rect 27524 9884 28644 9940
rect 29586 9884 29596 9940
rect 29652 9884 30492 9940
rect 30548 9884 30558 9940
rect 31154 9884 31164 9940
rect 31220 9884 32284 9940
rect 32340 9884 32350 9940
rect 33842 9884 33852 9940
rect 33908 9884 34692 9940
rect 38612 9884 43484 9940
rect 43540 9884 43550 9940
rect 51426 9884 51436 9940
rect 51492 9884 52332 9940
rect 52388 9884 52398 9940
rect 17602 9772 17612 9828
rect 17668 9772 19404 9828
rect 19460 9772 19470 9828
rect 26674 9772 26684 9828
rect 26740 9772 28028 9828
rect 28084 9772 28094 9828
rect 28588 9716 28644 9884
rect 34636 9828 34692 9884
rect 31378 9772 31388 9828
rect 31444 9772 31836 9828
rect 31892 9772 32172 9828
rect 32228 9772 32238 9828
rect 33282 9772 33292 9828
rect 33348 9772 34020 9828
rect 34626 9772 34636 9828
rect 34692 9772 35644 9828
rect 35700 9772 35710 9828
rect 36082 9772 36092 9828
rect 36148 9772 37100 9828
rect 37156 9772 37166 9828
rect 42578 9772 42588 9828
rect 42644 9772 43820 9828
rect 43876 9772 43886 9828
rect 51650 9772 51660 9828
rect 51716 9772 52892 9828
rect 52948 9772 52958 9828
rect 33964 9716 34020 9772
rect 16818 9660 16828 9716
rect 16884 9660 17948 9716
rect 18004 9660 18620 9716
rect 18676 9660 18956 9716
rect 19012 9660 19022 9716
rect 19842 9660 19852 9716
rect 19908 9660 23436 9716
rect 23492 9660 23502 9716
rect 28578 9660 28588 9716
rect 28644 9660 29932 9716
rect 29988 9660 29998 9716
rect 31042 9660 31052 9716
rect 31108 9660 33404 9716
rect 33460 9660 33470 9716
rect 33954 9660 33964 9716
rect 34020 9660 34188 9716
rect 34244 9660 34254 9716
rect 36530 9660 36540 9716
rect 36596 9660 40348 9716
rect 40404 9660 40414 9716
rect 51090 9660 51100 9716
rect 51156 9660 52556 9716
rect 52612 9660 52622 9716
rect 14690 9548 14700 9604
rect 14756 9548 15820 9604
rect 15876 9548 15886 9604
rect 19058 9548 19068 9604
rect 19124 9548 19180 9604
rect 19236 9548 21420 9604
rect 21476 9548 21486 9604
rect 30034 9548 30044 9604
rect 30100 9548 30604 9604
rect 30660 9548 30670 9604
rect 52882 9548 52892 9604
rect 52948 9548 54460 9604
rect 54516 9548 54526 9604
rect 29698 9436 29708 9492
rect 29764 9436 37324 9492
rect 37380 9436 37390 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 19058 9324 19068 9380
rect 19124 9324 19516 9380
rect 19572 9324 19582 9380
rect 37660 9212 39228 9268
rect 39284 9212 39844 9268
rect 40562 9212 40572 9268
rect 40628 9212 42812 9268
rect 42868 9212 43484 9268
rect 43540 9212 43550 9268
rect 47282 9212 47292 9268
rect 47348 9212 49756 9268
rect 49812 9212 49822 9268
rect 37660 9156 37716 9212
rect 39788 9156 39844 9212
rect 18162 9100 18172 9156
rect 18228 9100 18956 9156
rect 19012 9100 19404 9156
rect 19460 9100 19470 9156
rect 34514 9100 34524 9156
rect 34580 9100 35532 9156
rect 35588 9100 37660 9156
rect 37716 9100 37726 9156
rect 39778 9100 39788 9156
rect 39844 9100 39854 9156
rect 35074 8988 35084 9044
rect 35140 8988 35868 9044
rect 35924 8988 35934 9044
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 22418 8428 22428 8484
rect 22484 8428 25452 8484
rect 25508 8428 26572 8484
rect 26628 8428 26638 8484
rect 30930 8316 30940 8372
rect 30996 8316 34076 8372
rect 34132 8316 34142 8372
rect 47394 8316 47404 8372
rect 47460 8316 48636 8372
rect 48692 8316 49644 8372
rect 49700 8316 49710 8372
rect 50194 8316 50204 8372
rect 50260 8316 51100 8372
rect 51156 8316 51166 8372
rect 27346 8204 27356 8260
rect 27412 8204 36316 8260
rect 36372 8204 36382 8260
rect 39676 8204 40460 8260
rect 40516 8204 40526 8260
rect 44930 8204 44940 8260
rect 44996 8204 45612 8260
rect 45668 8204 45678 8260
rect 46386 8204 46396 8260
rect 46452 8204 47628 8260
rect 47684 8204 47694 8260
rect 48962 8204 48972 8260
rect 49028 8204 50764 8260
rect 50820 8204 51996 8260
rect 52052 8204 52062 8260
rect 39676 8148 39732 8204
rect 28018 8092 28028 8148
rect 28084 8092 39004 8148
rect 39060 8092 39676 8148
rect 39732 8092 39742 8148
rect 40002 8092 40012 8148
rect 40068 8092 47292 8148
rect 47348 8092 47358 8148
rect 47506 8092 47516 8148
rect 47572 8092 50428 8148
rect 50484 8092 51324 8148
rect 51380 8092 51390 8148
rect 18834 7868 18844 7924
rect 18900 7868 19628 7924
rect 19684 7868 19694 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 19282 7532 19292 7588
rect 19348 7532 21532 7588
rect 21588 7532 21598 7588
rect 26852 7476 26908 8036
rect 26964 7980 26974 8036
rect 29810 7980 29820 8036
rect 29876 7980 30716 8036
rect 30772 7980 30782 8036
rect 31154 7980 31164 8036
rect 31220 7980 31612 8036
rect 31668 7980 31678 8036
rect 33954 7980 33964 8036
rect 34020 7980 34972 8036
rect 35028 7980 35038 8036
rect 35522 7980 35532 8036
rect 35588 7980 36092 8036
rect 36148 7980 36158 8036
rect 41906 7980 41916 8036
rect 41972 7980 49420 8036
rect 49476 7980 49486 8036
rect 36306 7868 36316 7924
rect 36372 7868 38892 7924
rect 38948 7868 39900 7924
rect 39956 7868 40796 7924
rect 40852 7868 40862 7924
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 32498 7756 32508 7812
rect 32564 7756 42140 7812
rect 42196 7756 45836 7812
rect 45892 7756 46620 7812
rect 46676 7756 46686 7812
rect 30930 7644 30940 7700
rect 30996 7644 31500 7700
rect 31556 7644 31566 7700
rect 40002 7644 40012 7700
rect 40068 7644 41468 7700
rect 41524 7644 41534 7700
rect 43698 7644 43708 7700
rect 43764 7644 46172 7700
rect 46228 7644 46238 7700
rect 47954 7644 47964 7700
rect 48020 7644 48748 7700
rect 48804 7644 51436 7700
rect 51492 7644 51502 7700
rect 33954 7532 33964 7588
rect 34020 7532 35644 7588
rect 35700 7532 36428 7588
rect 36484 7532 36494 7588
rect 40114 7532 40124 7588
rect 40180 7532 41580 7588
rect 41636 7532 41860 7588
rect 43250 7532 43260 7588
rect 43316 7532 50876 7588
rect 50932 7532 50942 7588
rect 41804 7476 41860 7532
rect 18918 7420 18956 7476
rect 19012 7420 19022 7476
rect 26338 7420 26348 7476
rect 26404 7420 26908 7476
rect 27234 7420 27244 7476
rect 27300 7420 28140 7476
rect 28196 7420 28206 7476
rect 32610 7420 32620 7476
rect 32676 7420 33628 7476
rect 33684 7420 33694 7476
rect 34290 7420 34300 7476
rect 34356 7420 35420 7476
rect 35476 7420 35486 7476
rect 38098 7420 38108 7476
rect 38164 7420 38668 7476
rect 38724 7420 40684 7476
rect 40740 7420 40750 7476
rect 41804 7420 43820 7476
rect 43876 7420 43886 7476
rect 49858 7420 49868 7476
rect 49924 7420 50652 7476
rect 50708 7420 51660 7476
rect 51716 7420 51726 7476
rect 35420 7364 35476 7420
rect 21074 7308 21084 7364
rect 21140 7308 21644 7364
rect 21700 7308 21710 7364
rect 23762 7308 23772 7364
rect 23828 7308 25788 7364
rect 25844 7308 26796 7364
rect 26852 7308 26862 7364
rect 27010 7308 27020 7364
rect 27076 7308 27692 7364
rect 27748 7308 31724 7364
rect 31780 7308 31790 7364
rect 35420 7308 38220 7364
rect 38276 7308 39340 7364
rect 39396 7308 39406 7364
rect 49746 7308 49756 7364
rect 49812 7308 50092 7364
rect 50148 7308 50158 7364
rect 51538 7308 51548 7364
rect 51604 7308 52444 7364
rect 52500 7308 52510 7364
rect 18834 7196 18844 7252
rect 18900 7196 19964 7252
rect 20020 7196 20030 7252
rect 20738 7196 20748 7252
rect 20804 7196 21420 7252
rect 21476 7196 21486 7252
rect 24098 7196 24108 7252
rect 24164 7196 25900 7252
rect 25956 7196 25966 7252
rect 34962 7196 34972 7252
rect 35028 7196 35980 7252
rect 36036 7196 36046 7252
rect 36194 7196 36204 7252
rect 36260 7196 36764 7252
rect 36820 7196 42588 7252
rect 42644 7196 42654 7252
rect 20524 7084 21308 7140
rect 21364 7084 22764 7140
rect 22820 7084 23548 7140
rect 23604 7084 23614 7140
rect 36418 7084 36428 7140
rect 36484 7084 37548 7140
rect 37604 7084 38668 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 20524 7028 20580 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 38612 7028 38668 7084
rect 19058 6972 19068 7028
rect 19124 6972 20188 7028
rect 20244 6972 20254 7028
rect 20514 6972 20524 7028
rect 20580 6972 20590 7028
rect 23874 6972 23884 7028
rect 23940 6972 24444 7028
rect 24500 6972 24510 7028
rect 38612 6972 38780 7028
rect 38836 6972 38846 7028
rect 25890 6860 25900 6916
rect 25956 6860 27244 6916
rect 27300 6860 27310 6916
rect 17714 6748 17724 6804
rect 17780 6748 18620 6804
rect 18676 6748 18686 6804
rect 20178 6748 20188 6804
rect 20244 6748 22204 6804
rect 22260 6748 22270 6804
rect 23202 6748 23212 6804
rect 23268 6748 24332 6804
rect 24388 6748 24398 6804
rect 41580 6748 43260 6804
rect 43316 6748 43326 6804
rect 50194 6748 50204 6804
rect 50260 6748 50652 6804
rect 50708 6748 50718 6804
rect 51538 6748 51548 6804
rect 51604 6748 52668 6804
rect 52724 6748 52734 6804
rect 41580 6692 41636 6748
rect 15474 6636 15484 6692
rect 15540 6636 17500 6692
rect 17556 6636 18508 6692
rect 18564 6636 18574 6692
rect 19394 6636 19404 6692
rect 19460 6636 20300 6692
rect 20356 6636 20366 6692
rect 20626 6636 20636 6692
rect 20692 6636 21308 6692
rect 21364 6636 21374 6692
rect 23314 6636 23324 6692
rect 23380 6636 25116 6692
rect 25172 6636 25182 6692
rect 26226 6636 26236 6692
rect 26292 6636 27244 6692
rect 27300 6636 27310 6692
rect 30482 6636 30492 6692
rect 30548 6636 31836 6692
rect 31892 6636 32508 6692
rect 32564 6636 32574 6692
rect 38546 6636 38556 6692
rect 38612 6636 40460 6692
rect 40516 6636 41636 6692
rect 41794 6636 41804 6692
rect 41860 6636 50428 6692
rect 50484 6636 50494 6692
rect 52546 6636 52556 6692
rect 52612 6636 54796 6692
rect 54852 6636 54862 6692
rect 49420 6580 49476 6636
rect 16146 6524 16156 6580
rect 16212 6524 17388 6580
rect 17444 6524 17454 6580
rect 18946 6524 18956 6580
rect 19012 6524 21980 6580
rect 22036 6524 24108 6580
rect 24164 6524 24174 6580
rect 24994 6524 25004 6580
rect 25060 6524 26908 6580
rect 29362 6524 29372 6580
rect 29428 6524 31500 6580
rect 31556 6524 31566 6580
rect 39330 6524 39340 6580
rect 39396 6524 40236 6580
rect 40292 6524 40302 6580
rect 42914 6524 42924 6580
rect 42980 6524 45052 6580
rect 45108 6524 45118 6580
rect 46386 6524 46396 6580
rect 46452 6524 47180 6580
rect 47236 6524 47246 6580
rect 49410 6524 49420 6580
rect 49476 6524 49486 6580
rect 26852 6468 26908 6524
rect 19282 6412 19292 6468
rect 19348 6412 21196 6468
rect 21252 6412 21756 6468
rect 21812 6412 21822 6468
rect 22306 6412 22316 6468
rect 22372 6412 23660 6468
rect 23716 6412 23726 6468
rect 23874 6412 23884 6468
rect 23940 6412 26460 6468
rect 26516 6412 26526 6468
rect 26852 6412 27692 6468
rect 27748 6412 30716 6468
rect 30772 6412 30782 6468
rect 32162 6412 32172 6468
rect 32228 6412 43260 6468
rect 43316 6412 43932 6468
rect 43988 6412 43998 6468
rect 48402 6412 48412 6468
rect 48468 6412 50428 6468
rect 50484 6412 51212 6468
rect 51268 6412 51278 6468
rect 26460 6356 26516 6412
rect 20290 6300 20300 6356
rect 20356 6300 23996 6356
rect 24052 6300 24062 6356
rect 26460 6300 33628 6356
rect 33684 6300 33694 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 24098 6188 24108 6244
rect 24164 6188 26236 6244
rect 26292 6188 26302 6244
rect 30146 6188 30156 6244
rect 30212 6188 30492 6244
rect 30548 6188 31948 6244
rect 32004 6188 32014 6244
rect 20738 6076 20748 6132
rect 20804 6076 21644 6132
rect 21700 6076 21710 6132
rect 40002 6076 40012 6132
rect 40068 6076 43820 6132
rect 43876 6076 48300 6132
rect 48356 6076 48366 6132
rect 46498 5964 46508 6020
rect 46564 5964 47068 6020
rect 47124 5964 47134 6020
rect 21746 5852 21756 5908
rect 21812 5852 29372 5908
rect 29428 5852 29438 5908
rect 31378 5852 31388 5908
rect 31444 5852 32172 5908
rect 32228 5852 32238 5908
rect 45042 5852 45052 5908
rect 45108 5852 46732 5908
rect 46788 5852 46798 5908
rect 21298 5740 21308 5796
rect 21364 5740 22092 5796
rect 22148 5740 22158 5796
rect 30594 5740 30604 5796
rect 30660 5740 30940 5796
rect 30996 5740 31006 5796
rect 32050 5628 32060 5684
rect 32116 5628 44940 5684
rect 44996 5628 45276 5684
rect 45332 5628 45342 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 29698 5292 29708 5348
rect 29764 5292 30940 5348
rect 30996 5292 31006 5348
rect 37650 5292 37660 5348
rect 37716 5292 39564 5348
rect 39620 5292 39630 5348
rect 18498 5180 18508 5236
rect 18564 5180 21420 5236
rect 21476 5180 21486 5236
rect 34626 5180 34636 5236
rect 34692 5180 35644 5236
rect 35700 5180 35710 5236
rect 40338 5180 40348 5236
rect 40404 5180 40908 5236
rect 40964 5180 41244 5236
rect 41300 5180 41310 5236
rect 30930 5068 30940 5124
rect 30996 5068 32060 5124
rect 32116 5068 32126 5124
rect 38210 5068 38220 5124
rect 38276 5068 39116 5124
rect 39172 5068 39182 5124
rect 44594 5068 44604 5124
rect 44660 5068 45500 5124
rect 45556 5068 46396 5124
rect 46452 5068 46462 5124
rect 47058 5068 47068 5124
rect 47124 5068 50316 5124
rect 50372 5068 50382 5124
rect 50316 5012 50372 5068
rect 50316 4956 53340 5012
rect 53396 4956 55468 5012
rect 55524 4956 55534 5012
rect 51314 4844 51324 4900
rect 51380 4844 52668 4900
rect 52724 4844 52734 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 26852 4508 28588 4564
rect 28644 4508 30380 4564
rect 30436 4508 30446 4564
rect 46946 4508 46956 4564
rect 47012 4508 48748 4564
rect 48804 4508 48814 4564
rect 26852 4340 26908 4508
rect 40786 4396 40796 4452
rect 40852 4396 41692 4452
rect 41748 4396 41758 4452
rect 25330 4284 25340 4340
rect 25396 4284 26908 4340
rect 46946 4284 46956 4340
rect 47012 4284 57596 4340
rect 57652 4284 57662 4340
rect 46050 4172 46060 4228
rect 46116 4172 47068 4228
rect 47124 4172 48524 4228
rect 48580 4172 48590 4228
rect 57362 4172 57372 4228
rect 57428 4172 58156 4228
rect 58212 4172 58222 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 59200 3668 60000 3696
rect 58146 3612 58156 3668
rect 58212 3612 60000 3668
rect 59200 3584 60000 3612
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 49084 63084 49140 63140
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 49084 60956 49140 61012
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4284 51324 4340 51380
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 4284 50316 4340 50372
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 31500 46732 31556 46788
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 37212 45836 37268 45892
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 38220 43820 38276 43876
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 57484 41804 57540 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 20300 40348 20356 40404
rect 57484 40348 57540 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 31500 39676 31556 39732
rect 20188 39564 20244 39620
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 46060 38780 46116 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 46060 37996 46116 38052
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 20188 37436 20244 37492
rect 20300 37324 20356 37380
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 38220 34076 38276 34132
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 48972 33628 49028 33684
rect 49084 33516 49140 33572
rect 22204 33180 22260 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 22204 31052 22260 31108
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 48972 30044 49028 30100
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 49084 28924 49140 28980
rect 14700 28588 14756 28644
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 14700 26572 14756 26628
rect 25564 26572 25620 26628
rect 25564 25900 25620 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 26348 25340 26404 25396
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 25564 24892 25620 24948
rect 26348 24892 26404 24948
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 40684 22428 40740 22484
rect 37212 22316 37268 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 40908 21756 40964 21812
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 38892 20076 38948 20132
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 38892 19292 38948 19348
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 52108 18956 52164 19012
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 51324 18060 51380 18116
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 52108 17836 52164 17892
rect 40908 17612 40964 17668
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 51324 16716 51380 16772
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 40684 15932 40740 15988
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 18956 10780 19012 10836
rect 19180 10556 19236 10612
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19180 9548 19236 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 18956 7420 19012 7476
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 66668 4768 66700
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4284 51380 4340 51390
rect 4284 50372 4340 51324
rect 4284 50306 4340 50316
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 19808 65884 20128 66700
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 35168 66668 35488 66700
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 50528 65884 50848 66700
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 49084 63140 49140 63150
rect 49084 61012 49140 63084
rect 49084 60946 49140 60956
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 31500 46788 31556 46798
rect 20300 40404 20356 40414
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 20188 39620 20244 39630
rect 20188 37492 20244 39564
rect 20188 37426 20244 37436
rect 20300 37380 20356 40348
rect 31500 39732 31556 46732
rect 31500 39666 31556 39676
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 20300 37314 20356 37324
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 22204 33236 22260 33246
rect 22204 31108 22260 33180
rect 22204 31042 22260 31052
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 14700 28644 14756 28654
rect 14700 26628 14756 28588
rect 14700 26562 14756 26572
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 25564 26628 25620 26638
rect 25564 25956 25620 26572
rect 25564 24948 25620 25900
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 25564 24882 25620 24892
rect 26348 25396 26404 25406
rect 26348 24948 26404 25340
rect 26348 24882 26404 24892
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 18956 10836 19012 10846
rect 18956 7476 19012 10780
rect 19180 10612 19236 10622
rect 19180 9604 19236 10556
rect 19180 9538 19236 9548
rect 18956 7410 19012 7420
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 37212 45892 37268 45902
rect 37212 22372 37268 45836
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 38220 43876 38276 43886
rect 38220 34132 38276 43820
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 57484 41860 57540 41870
rect 57484 40404 57540 41804
rect 57484 40338 57540 40348
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 46060 38836 46116 38846
rect 46060 38052 46116 38780
rect 46060 37986 46116 37996
rect 38220 34066 38276 34076
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 48972 33684 49028 33694
rect 48972 30100 49028 33628
rect 48972 30034 49028 30044
rect 49084 33572 49140 33582
rect 49084 28980 49140 33516
rect 49084 28914 49140 28924
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 37212 22306 37268 22316
rect 40684 22484 40740 22494
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 38892 20132 38948 20142
rect 38892 19348 38948 20076
rect 38892 19282 38948 19292
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 40684 15988 40740 22428
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 40908 21812 40964 21822
rect 40908 17668 40964 21756
rect 40908 17602 40964 17612
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 40684 15922 40740 15932
rect 50528 17276 50848 18788
rect 52108 19012 52164 19022
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 15708 50848 17220
rect 51324 18116 51380 18126
rect 51324 16772 51380 18060
rect 52108 17892 52164 18956
rect 52108 17826 52164 17836
rect 51324 16706 51380 16716
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 27552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 26544 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1261_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 25088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23744 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1263_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 25872 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1264_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1265_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 26992 0 -1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1266_
timestamp 1694700623
transform -1 0 24192 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1267_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 25088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1268_
timestamp 1694700623
transform -1 0 23520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1269_
timestamp 1694700623
transform -1 0 22848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1270_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 25760 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22400 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1272_
timestamp 1694700623
transform 1 0 27328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1273_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 28336 0 -1 40768
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1274_
timestamp 1694700623
transform 1 0 23968 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1275_
timestamp 1694700623
transform -1 0 24864 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1276_
timestamp 1694700623
transform -1 0 24864 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1277_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 22512 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1278_
timestamp 1694700623
transform 1 0 23184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1279_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 28336 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1280_
timestamp 1694700623
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1281_
timestamp 1694700623
transform -1 0 36064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1282_
timestamp 1694700623
transform -1 0 34384 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1283_
timestamp 1694700623
transform -1 0 32256 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1284_
timestamp 1694700623
transform 1 0 33936 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1285_
timestamp 1694700623
transform 1 0 38304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1286_
timestamp 1694700623
transform -1 0 35840 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1287_
timestamp 1694700623
transform 1 0 38080 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1288_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1289_
timestamp 1694700623
transform -1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1694700623
transform -1 0 38304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1291_
timestamp 1694700623
transform -1 0 36288 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1292_
timestamp 1694700623
transform 1 0 35056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1293_
timestamp 1694700623
transform 1 0 36960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1294_
timestamp 1694700623
transform 1 0 32928 0 -1 37632
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1295_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 33824 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1296_
timestamp 1694700623
transform -1 0 33824 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1694700623
transform 1 0 37856 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1298_
timestamp 1694700623
transform -1 0 36512 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1299_
timestamp 1694700623
transform -1 0 35280 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1300_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 33936 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1301_
timestamp 1694700623
transform -1 0 20160 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1302_
timestamp 1694700623
transform 1 0 20496 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1303_
timestamp 1694700623
transform 1 0 18368 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1304_
timestamp 1694700623
transform -1 0 20496 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1305_
timestamp 1694700623
transform 1 0 18480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1306_
timestamp 1694700623
transform -1 0 18144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1307_
timestamp 1694700623
transform -1 0 16464 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1308_
timestamp 1694700623
transform 1 0 15344 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1309_
timestamp 1694700623
transform 1 0 20160 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1310_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 16464 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1311_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 16352 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1312_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15120 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1313_
timestamp 1694700623
transform 1 0 18480 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1314_
timestamp 1694700623
transform 1 0 17584 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1315_
timestamp 1694700623
transform 1 0 18032 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1316_
timestamp 1694700623
transform 1 0 16464 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1317_
timestamp 1694700623
transform -1 0 16576 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1318_
timestamp 1694700623
transform 1 0 7504 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1319_
timestamp 1694700623
transform 1 0 11200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1320_
timestamp 1694700623
transform -1 0 8512 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1321_
timestamp 1694700623
transform 1 0 8848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1322_
timestamp 1694700623
transform 1 0 7392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1323_
timestamp 1694700623
transform 1 0 9408 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1324_
timestamp 1694700623
transform -1 0 11648 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1325_
timestamp 1694700623
transform 1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1326_
timestamp 1694700623
transform -1 0 11200 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1327_
timestamp 1694700623
transform -1 0 11648 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1328_
timestamp 1694700623
transform -1 0 13104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1329_
timestamp 1694700623
transform -1 0 12768 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1330_
timestamp 1694700623
transform -1 0 11536 0 -1 32928
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1331_
timestamp 1694700623
transform 1 0 8400 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1332_
timestamp 1694700623
transform 1 0 11648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1333_
timestamp 1694700623
transform -1 0 14672 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1334_
timestamp 1694700623
transform 1 0 12544 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1335_
timestamp 1694700623
transform -1 0 13104 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1336_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 11872 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 11312 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1338_
timestamp 1694700623
transform 1 0 33264 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 35392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1340_
timestamp 1694700623
transform 1 0 34496 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1341_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 38192 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 37408 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1343_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 24416 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1344_
timestamp 1694700623
transform 1 0 23856 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 27664 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1346_
timestamp 1694700623
transform 1 0 34272 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1347_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 38192 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1348_
timestamp 1694700623
transform -1 0 39536 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1349_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 38976 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1350_
timestamp 1694700623
transform 1 0 36848 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1351_
timestamp 1694700623
transform -1 0 35840 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 35504 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 37520 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1354_
timestamp 1694700623
transform -1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1355_
timestamp 1694700623
transform -1 0 19376 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1356_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 19824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1357_
timestamp 1694700623
transform 1 0 18032 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1358_
timestamp 1694700623
transform -1 0 21056 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1359_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 17024 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1360_
timestamp 1694700623
transform 1 0 16128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1361_
timestamp 1694700623
transform 1 0 17360 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1362_
timestamp 1694700623
transform -1 0 12656 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1363_
timestamp 1694700623
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1364_
timestamp 1694700623
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1365_
timestamp 1694700623
transform -1 0 13104 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1366_
timestamp 1694700623
transform 1 0 11648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1367_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13328 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1694700623
transform -1 0 12768 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 15568 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1370_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 10752 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1371_
timestamp 1694700623
transform 1 0 38304 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1372_
timestamp 1694700623
transform -1 0 37968 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 37408 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 38080 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1375_
timestamp 1694700623
transform 1 0 37408 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1376_
timestamp 1694700623
transform -1 0 11200 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1377_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 14448 0 -1 29792
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1378_
timestamp 1694700623
transform 1 0 13328 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1379_
timestamp 1694700623
transform -1 0 14896 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1380_
timestamp 1694700623
transform -1 0 14784 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1381_
timestamp 1694700623
transform 1 0 14560 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1382_
timestamp 1694700623
transform -1 0 8848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1383_
timestamp 1694700623
transform 1 0 8288 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1694700623
transform 1 0 8736 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1385_
timestamp 1694700623
transform 1 0 7280 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1386_
timestamp 1694700623
transform -1 0 9744 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1387_
timestamp 1694700623
transform -1 0 11536 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1388_
timestamp 1694700623
transform -1 0 11312 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1389_
timestamp 1694700623
transform 1 0 11424 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1390_
timestamp 1694700623
transform -1 0 13104 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1391_
timestamp 1694700623
transform -1 0 19824 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1392_
timestamp 1694700623
transform 1 0 17920 0 1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1694700623
transform 1 0 18480 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1394_
timestamp 1694700623
transform 1 0 17360 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1395_
timestamp 1694700623
transform -1 0 15344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1396_
timestamp 1694700623
transform 1 0 17248 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1397_
timestamp 1694700623
transform 1 0 15792 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1398_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 15344 0 1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1399_
timestamp 1694700623
transform 1 0 15120 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1400_
timestamp 1694700623
transform -1 0 36960 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1401_
timestamp 1694700623
transform 1 0 34384 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1402_
timestamp 1694700623
transform -1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1403_
timestamp 1694700623
transform 1 0 36848 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1404_
timestamp 1694700623
transform -1 0 32704 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1405_
timestamp 1694700623
transform 1 0 31360 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1406_
timestamp 1694700623
transform 1 0 30800 0 1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1407_
timestamp 1694700623
transform 1 0 22848 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1408_
timestamp 1694700623
transform -1 0 28000 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1409_
timestamp 1694700623
transform 1 0 25760 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1410_
timestamp 1694700623
transform -1 0 25984 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1411_
timestamp 1694700623
transform -1 0 28784 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1412_
timestamp 1694700623
transform -1 0 27888 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1413_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 24640 0 1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1414_
timestamp 1694700623
transform -1 0 26432 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1415_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 17360 0 -1 47040
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1694700623
transform 1 0 35616 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1417_
timestamp 1694700623
transform 1 0 36176 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1418_
timestamp 1694700623
transform 1 0 38304 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1419_
timestamp 1694700623
transform 1 0 17136 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_
timestamp 1694700623
transform -1 0 26096 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1421_
timestamp 1694700623
transform -1 0 24976 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1422_
timestamp 1694700623
transform -1 0 24864 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1423_
timestamp 1694700623
transform -1 0 24864 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1424_
timestamp 1694700623
transform -1 0 38080 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1694700623
transform -1 0 32704 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1426_
timestamp 1694700623
transform -1 0 36176 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1427_
timestamp 1694700623
transform 1 0 31472 0 1 32928
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1428_
timestamp 1694700623
transform -1 0 24416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1429_
timestamp 1694700623
transform 1 0 23520 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1694700623
transform -1 0 26320 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1694700623
transform -1 0 28224 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1432_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 26208 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1433_
timestamp 1694700623
transform -1 0 28336 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1434_
timestamp 1694700623
transform 1 0 12432 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1694700623
transform 1 0 12432 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1436_
timestamp 1694700623
transform 1 0 13328 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1437_
timestamp 1694700623
transform 1 0 15008 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1438_
timestamp 1694700623
transform 1 0 17248 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1439_
timestamp 1694700623
transform 1 0 17248 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1440_
timestamp 1694700623
transform 1 0 16128 0 1 42336
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1441_
timestamp 1694700623
transform 1 0 14224 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1442_
timestamp 1694700623
transform -1 0 14000 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1443_
timestamp 1694700623
transform -1 0 15344 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1444_
timestamp 1694700623
transform 1 0 15344 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1445_
timestamp 1694700623
transform 1 0 17024 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1446_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 25536 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1447_
timestamp 1694700623
transform 1 0 34272 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1448_
timestamp 1694700623
transform 1 0 34608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1449_
timestamp 1694700623
transform 1 0 35952 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1450_
timestamp 1694700623
transform 1 0 25648 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1694700623
transform 1 0 28224 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1694700623
transform -1 0 27776 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1694700623
transform 1 0 28112 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 27104 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1694700623
transform 1 0 26768 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1456_
timestamp 1694700623
transform 1 0 29568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1457_
timestamp 1694700623
transform -1 0 31360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1458_
timestamp 1694700623
transform -1 0 33264 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1459_
timestamp 1694700623
transform 1 0 31136 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1460_
timestamp 1694700623
transform 1 0 14112 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1461_
timestamp 1694700623
transform -1 0 11424 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1462_
timestamp 1694700623
transform 1 0 13552 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1463_
timestamp 1694700623
transform 1 0 14224 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1694700623
transform -1 0 14224 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1465_
timestamp 1694700623
transform -1 0 14336 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1466_
timestamp 1694700623
transform -1 0 14336 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1694700623
transform 1 0 15232 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1468_
timestamp 1694700623
transform 1 0 15120 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1694700623
transform 1 0 32928 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1470_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 34496 0 1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1471_
timestamp 1694700623
transform 1 0 37520 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1472_
timestamp 1694700623
transform 1 0 38752 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1473_
timestamp 1694700623
transform 1 0 34720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1474_
timestamp 1694700623
transform 1 0 36064 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1475_
timestamp 1694700623
transform -1 0 31808 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1476_
timestamp 1694700623
transform 1 0 31808 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1477_
timestamp 1694700623
transform 1 0 32592 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1478_
timestamp 1694700623
transform -1 0 33712 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 28336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_
timestamp 1694700623
transform 1 0 29232 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1481_
timestamp 1694700623
transform 1 0 29680 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1482_
timestamp 1694700623
transform 1 0 31024 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_
timestamp 1694700623
transform 1 0 31248 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1694700623
transform 1 0 13888 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1485_
timestamp 1694700623
transform 1 0 14336 0 -1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1486_
timestamp 1694700623
transform 1 0 15232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1487_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 13440 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1488_
timestamp 1694700623
transform 1 0 8512 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1489_
timestamp 1694700623
transform 1 0 9408 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1694700623
transform 1 0 8624 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1491_
timestamp 1694700623
transform -1 0 10192 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1492_
timestamp 1694700623
transform 1 0 13328 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1694700623
transform -1 0 15456 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 14672 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1495_
timestamp 1694700623
transform 1 0 15792 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1496_
timestamp 1694700623
transform 1 0 33264 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1497_
timestamp 1694700623
transform 1 0 35056 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1498_
timestamp 1694700623
transform 1 0 36848 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1694700623
transform -1 0 42672 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1694700623
transform -1 0 31472 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1694700623
transform -1 0 30576 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1694700623
transform -1 0 30016 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1503_
timestamp 1694700623
transform 1 0 30576 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1504_
timestamp 1694700623
transform -1 0 31808 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1505_
timestamp 1694700623
transform 1 0 26320 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1506_
timestamp 1694700623
transform -1 0 29568 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1507_
timestamp 1694700623
transform -1 0 29568 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1508_
timestamp 1694700623
transform 1 0 28336 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1694700623
transform 1 0 28224 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1510_
timestamp 1694700623
transform 1 0 29008 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1511_
timestamp 1694700623
transform 1 0 30352 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1512_
timestamp 1694700623
transform -1 0 20944 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1694700623
transform 1 0 20160 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1514_
timestamp 1694700623
transform 1 0 20272 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1515_
timestamp 1694700623
transform -1 0 18032 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1516_
timestamp 1694700623
transform -1 0 10080 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1694700623
transform 1 0 7728 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 9184 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1519_
timestamp 1694700623
transform 1 0 9408 0 -1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1520_
timestamp 1694700623
transform 1 0 10864 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1521_
timestamp 1694700623
transform -1 0 13552 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1522_
timestamp 1694700623
transform -1 0 15120 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1523_
timestamp 1694700623
transform 1 0 14896 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1524_
timestamp 1694700623
transform 1 0 32592 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1694700623
transform -1 0 31248 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1694700623
transform -1 0 31808 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1527_
timestamp 1694700623
transform 1 0 31808 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1528_
timestamp 1694700623
transform 1 0 32592 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1529_
timestamp 1694700623
transform 1 0 33376 0 -1 56448
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1530_
timestamp 1694700623
transform 1 0 35280 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1694700623
transform -1 0 36960 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1532_
timestamp 1694700623
transform -1 0 36624 0 1 53312
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1533_
timestamp 1694700623
transform 1 0 36848 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1534_
timestamp 1694700623
transform 1 0 41888 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1535_
timestamp 1694700623
transform 1 0 34384 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1694700623
transform -1 0 36624 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1694700623
transform -1 0 31248 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1538_
timestamp 1694700623
transform 1 0 29904 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1694700623
transform 1 0 31248 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1694700623
transform -1 0 32592 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1541_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 31696 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1694700623
transform 1 0 11312 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1543_
timestamp 1694700623
transform -1 0 12096 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1544_
timestamp 1694700623
transform 1 0 14672 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1545_
timestamp 1694700623
transform 1 0 14896 0 -1 40768
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1694700623
transform 1 0 12656 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1694700623
transform -1 0 11760 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1548_
timestamp 1694700623
transform -1 0 12656 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1694700623
transform 1 0 11872 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1550_
timestamp 1694700623
transform 1 0 13776 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1551_
timestamp 1694700623
transform -1 0 11536 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1694700623
transform -1 0 10864 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1694700623
transform 1 0 10864 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1554_
timestamp 1694700623
transform 1 0 14336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1555_
timestamp 1694700623
transform -1 0 14896 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1556_
timestamp 1694700623
transform 1 0 14784 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1694700623
transform 1 0 24304 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1558_
timestamp 1694700623
transform 1 0 25088 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1694700623
transform -1 0 30800 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1560_
timestamp 1694700623
transform 1 0 30576 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1561_
timestamp 1694700623
transform 1 0 25648 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1694700623
transform 1 0 26992 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1563_
timestamp 1694700623
transform 1 0 26432 0 -1 58016
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1564_
timestamp 1694700623
transform 1 0 35952 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1565_
timestamp 1694700623
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1694700623
transform 1 0 35840 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1567_
timestamp 1694700623
transform 1 0 35392 0 -1 56448
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1694700623
transform -1 0 36624 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1694700623
transform -1 0 25648 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1694700623
transform -1 0 26432 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1694700623
transform -1 0 25760 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1572_
timestamp 1694700623
transform 1 0 26656 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1573_
timestamp 1694700623
transform -1 0 31472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1574_
timestamp 1694700623
transform -1 0 30240 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1694700623
transform -1 0 28112 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1576_
timestamp 1694700623
transform 1 0 27664 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1694700623
transform -1 0 27552 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1694700623
transform 1 0 26992 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1694700623
transform -1 0 29568 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1694700623
transform -1 0 15904 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1694700623
transform -1 0 14000 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1582_
timestamp 1694700623
transform -1 0 13216 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1694700623
transform -1 0 11984 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1694700623
transform -1 0 10528 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1585_
timestamp 1694700623
transform 1 0 9968 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1694700623
transform -1 0 13440 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1587_
timestamp 1694700623
transform 1 0 10976 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1588_
timestamp 1694700623
transform 1 0 12096 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1589_
timestamp 1694700623
transform 1 0 12208 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1590_
timestamp 1694700623
transform 1 0 13216 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1591_
timestamp 1694700623
transform -1 0 15344 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1592_
timestamp 1694700623
transform 1 0 13328 0 1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1593_
timestamp 1694700623
transform 1 0 28448 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1594_
timestamp 1694700623
transform 1 0 35616 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1595_
timestamp 1694700623
transform 1 0 40768 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1694700623
transform 1 0 42784 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1694700623
transform 1 0 35056 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1694700623
transform 1 0 34496 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1599_
timestamp 1694700623
transform 1 0 35392 0 -1 59584
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1600_
timestamp 1694700623
transform 1 0 27552 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1601_
timestamp 1694700623
transform -1 0 34384 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1602_
timestamp 1694700623
transform -1 0 31472 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1603_
timestamp 1694700623
transform 1 0 30912 0 1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1604_
timestamp 1694700623
transform -1 0 14896 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1694700623
transform 1 0 16016 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1606_
timestamp 1694700623
transform 1 0 16016 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1694700623
transform 1 0 16240 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1694700623
transform -1 0 16240 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1694700623
transform 1 0 17808 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1694700623
transform 1 0 16016 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1611_
timestamp 1694700623
transform 1 0 12208 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1694700623
transform -1 0 14112 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1613_
timestamp 1694700623
transform -1 0 14448 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1694700623
transform -1 0 15344 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1615_
timestamp 1694700623
transform 1 0 16576 0 1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1616_
timestamp 1694700623
transform 1 0 32928 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1617_
timestamp 1694700623
transform 1 0 34272 0 -1 61152
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1618_
timestamp 1694700623
transform 1 0 36736 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1619_
timestamp 1694700623
transform 1 0 47040 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1694700623
transform 1 0 31808 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1694700623
transform -1 0 30912 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1694700623
transform 1 0 32256 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1694700623
transform -1 0 33376 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1694700623
transform -1 0 32928 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1694700623
transform 1 0 17248 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1626_
timestamp 1694700623
transform 1 0 17248 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1627_
timestamp 1694700623
transform 1 0 37408 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1628_
timestamp 1694700623
transform 1 0 34048 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1629_
timestamp 1694700623
transform -1 0 37744 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1694700623
transform 1 0 38304 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1631_
timestamp 1694700623
transform 1 0 52304 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1694700623
transform 1 0 38080 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1633_
timestamp 1694700623
transform -1 0 40320 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1634_
timestamp 1694700623
transform 1 0 52864 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1635_
timestamp 1694700623
transform -1 0 53424 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1636_
timestamp 1694700623
transform -1 0 55104 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1694700623
transform 1 0 50624 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1638_
timestamp 1694700623
transform 1 0 51632 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1639_
timestamp 1694700623
transform -1 0 50512 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1640_
timestamp 1694700623
transform 1 0 29792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1694700623
transform -1 0 35168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1694700623
transform -1 0 40320 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1643_
timestamp 1694700623
transform -1 0 29792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1694700623
transform -1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1645_
timestamp 1694700623
transform 1 0 23408 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1646_
timestamp 1694700623
transform 1 0 29008 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1647_
timestamp 1694700623
transform 1 0 32928 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1694700623
transform -1 0 31584 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1649_
timestamp 1694700623
transform -1 0 32032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1694700623
transform -1 0 31472 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1694700623
transform 1 0 35280 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1652_
timestamp 1694700623
transform 1 0 35616 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1653_
timestamp 1694700623
transform 1 0 34384 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1654_
timestamp 1694700623
transform 1 0 30240 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1655_
timestamp 1694700623
transform -1 0 57568 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1656_
timestamp 1694700623
transform -1 0 34944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1657_
timestamp 1694700623
transform 1 0 33600 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1694700623
transform 1 0 21168 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1659_
timestamp 1694700623
transform 1 0 23072 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1660_
timestamp 1694700623
transform -1 0 42672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1661_
timestamp 1694700623
transform 1 0 31360 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1662_
timestamp 1694700623
transform 1 0 30464 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1663_
timestamp 1694700623
transform -1 0 34160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1664_
timestamp 1694700623
transform -1 0 33824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1665_
timestamp 1694700623
transform -1 0 31136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1666_
timestamp 1694700623
transform -1 0 31360 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1667_
timestamp 1694700623
transform -1 0 58016 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1694700623
transform -1 0 44352 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1694700623
transform 1 0 31136 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1694700623
transform 1 0 30912 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1671_
timestamp 1694700623
transform -1 0 49056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1694700623
transform -1 0 39536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1673_
timestamp 1694700623
transform 1 0 40432 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1694700623
transform 1 0 40768 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1675_
timestamp 1694700623
transform 1 0 42672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1694700623
transform 1 0 43344 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1694700623
transform 1 0 46032 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1678_
timestamp 1694700623
transform 1 0 46592 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1679_
timestamp 1694700623
transform 1 0 46032 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1694700623
transform 1 0 45136 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1681_
timestamp 1694700623
transform 1 0 43680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1682_
timestamp 1694700623
transform 1 0 45696 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1683_
timestamp 1694700623
transform 1 0 44912 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1694700623
transform 1 0 43456 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1685_
timestamp 1694700623
transform 1 0 42784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1686_
timestamp 1694700623
transform -1 0 49952 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1694700623
transform 1 0 30016 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1688_
timestamp 1694700623
transform 1 0 39536 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1694700623
transform 1 0 44464 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1694700623
transform 1 0 45360 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1694700623
transform -1 0 47600 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1692_
timestamp 1694700623
transform 1 0 46592 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1693_
timestamp 1694700623
transform 1 0 46816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1694_
timestamp 1694700623
transform 1 0 46480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1694700623
transform 1 0 47376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1696_
timestamp 1694700623
transform 1 0 45472 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1697_
timestamp 1694700623
transform -1 0 21840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1698_
timestamp 1694700623
transform 1 0 20048 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1699_
timestamp 1694700623
transform -1 0 46928 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1700_
timestamp 1694700623
transform 1 0 45584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1701_
timestamp 1694700623
transform 1 0 40992 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1702_
timestamp 1694700623
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1703_
timestamp 1694700623
transform 1 0 49952 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1694700623
transform -1 0 49504 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1705_
timestamp 1694700623
transform -1 0 42336 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1694700623
transform -1 0 40544 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1707_
timestamp 1694700623
transform 1 0 38528 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1694700623
transform 1 0 40768 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1709_
timestamp 1694700623
transform 1 0 38752 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1710_
timestamp 1694700623
transform 1 0 39424 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1711_
timestamp 1694700623
transform -1 0 40544 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1712_
timestamp 1694700623
transform 1 0 21168 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1713_
timestamp 1694700623
transform 1 0 22512 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1714_
timestamp 1694700623
transform 1 0 22064 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1694700623
transform 1 0 49056 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1716_
timestamp 1694700623
transform -1 0 49504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1717_
timestamp 1694700623
transform -1 0 24528 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1694700623
transform 1 0 21504 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1694700623
transform 1 0 22064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1720_
timestamp 1694700623
transform 1 0 22960 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1721_
timestamp 1694700623
transform -1 0 24192 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1694700623
transform 1 0 23296 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1694700623
transform -1 0 24864 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1724_
timestamp 1694700623
transform -1 0 25088 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1725_
timestamp 1694700623
transform -1 0 23856 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1726_
timestamp 1694700623
transform 1 0 19488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1694700623
transform 1 0 19264 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1694700623
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1694700623
transform 1 0 19824 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1694700623
transform 1 0 19040 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1694700623
transform 1 0 21280 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1732_
timestamp 1694700623
transform -1 0 21280 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1733_
timestamp 1694700623
transform -1 0 19712 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1734_
timestamp 1694700623
transform 1 0 6832 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1735_
timestamp 1694700623
transform 1 0 18480 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1694700623
transform -1 0 18480 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1694700623
transform -1 0 20832 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1738_
timestamp 1694700623
transform -1 0 20272 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1739_
timestamp 1694700623
transform 1 0 20048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1740_
timestamp 1694700623
transform -1 0 24864 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1694700623
transform -1 0 22848 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1694700623
transform -1 0 23520 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1743_
timestamp 1694700623
transform 1 0 23744 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1744_
timestamp 1694700623
transform 1 0 23520 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1745_
timestamp 1694700623
transform -1 0 24752 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1746_
timestamp 1694700623
transform 1 0 22512 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1694700623
transform 1 0 23408 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1694700623
transform -1 0 24976 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1749_
timestamp 1694700623
transform -1 0 24864 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1750_
timestamp 1694700623
transform -1 0 25760 0 1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1694700623
transform -1 0 23184 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1752_
timestamp 1694700623
transform -1 0 22064 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1753_
timestamp 1694700623
transform 1 0 24752 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1754_
timestamp 1694700623
transform 1 0 25760 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1755_
timestamp 1694700623
transform 1 0 25088 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1756_
timestamp 1694700623
transform 1 0 25760 0 1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1757_
timestamp 1694700623
transform -1 0 21168 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1694700623
transform -1 0 18368 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1694700623
transform -1 0 19936 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1760_
timestamp 1694700623
transform -1 0 20496 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1761_
timestamp 1694700623
transform -1 0 20832 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1694700623
transform -1 0 11872 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1763_
timestamp 1694700623
transform 1 0 3472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1694700623
transform 1 0 2576 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1694700623
transform -1 0 4256 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1766_
timestamp 1694700623
transform -1 0 4816 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1694700623
transform -1 0 3248 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1768_
timestamp 1694700623
transform -1 0 5488 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1694700623
transform -1 0 6048 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1770_
timestamp 1694700623
transform -1 0 5264 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1771_
timestamp 1694700623
transform -1 0 6384 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1694700623
transform -1 0 5264 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1773_
timestamp 1694700623
transform -1 0 3808 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1774_
timestamp 1694700623
transform -1 0 4144 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1775_
timestamp 1694700623
transform -1 0 3024 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1694700623
transform -1 0 5264 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1777_
timestamp 1694700623
transform -1 0 5264 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1778_
timestamp 1694700623
transform -1 0 5824 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1779_
timestamp 1694700623
transform -1 0 2912 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1694700623
transform -1 0 6160 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1694700623
transform -1 0 6384 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1782_
timestamp 1694700623
transform -1 0 5824 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1783_
timestamp 1694700623
transform 1 0 4816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1694700623
transform 1 0 2912 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1785_
timestamp 1694700623
transform -1 0 4592 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1694700623
transform 1 0 4256 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1694700623
transform 1 0 3136 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1694700623
transform 1 0 5488 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1789_
timestamp 1694700623
transform -1 0 6272 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1790_
timestamp 1694700623
transform -1 0 4144 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1791_
timestamp 1694700623
transform -1 0 7504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1694700623
transform 1 0 3584 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1694700623
transform 1 0 2688 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1794_
timestamp 1694700623
transform 1 0 4144 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1694700623
transform 1 0 4816 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1694700623
transform -1 0 5040 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1797_
timestamp 1694700623
transform -1 0 6160 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1694700623
transform 1 0 4144 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1694700623
transform 1 0 3696 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1800_
timestamp 1694700623
transform -1 0 48608 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1801_
timestamp 1694700623
transform -1 0 20944 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1694700623
transform 1 0 5488 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1803_
timestamp 1694700623
transform -1 0 6384 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1694700623
transform 1 0 6160 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1805_
timestamp 1694700623
transform 1 0 5824 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1806_
timestamp 1694700623
transform -1 0 7952 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1807_
timestamp 1694700623
transform -1 0 6608 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1694700623
transform 1 0 6608 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1809_
timestamp 1694700623
transform -1 0 7952 0 1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1810_
timestamp 1694700623
transform 1 0 8736 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1811_
timestamp 1694700623
transform -1 0 8848 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1694700623
transform -1 0 7504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1813_
timestamp 1694700623
transform 1 0 6384 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1694700623
transform 1 0 7728 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1694700623
transform 1 0 8288 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1816_
timestamp 1694700623
transform 1 0 9408 0 -1 62720
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1817_
timestamp 1694700623
transform -1 0 20944 0 1 59584
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1818_
timestamp 1694700623
transform 1 0 19824 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1819_
timestamp 1694700623
transform -1 0 19712 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1820_
timestamp 1694700623
transform 1 0 35504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1821_
timestamp 1694700623
transform -1 0 42896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1822_
timestamp 1694700623
transform 1 0 19712 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1823_
timestamp 1694700623
transform -1 0 20160 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1824_
timestamp 1694700623
transform -1 0 12992 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1694700623
transform -1 0 6832 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1694700623
transform 1 0 5712 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1827_
timestamp 1694700623
transform 1 0 7728 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1828_
timestamp 1694700623
transform -1 0 10416 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1694700623
transform -1 0 9296 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1694700623
transform -1 0 9184 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1694700623
transform 1 0 9408 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1832_
timestamp 1694700623
transform -1 0 11088 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1694700623
transform -1 0 9296 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1694700623
transform 1 0 7616 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1835_
timestamp 1694700623
transform 1 0 7840 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1694700623
transform 1 0 7056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1694700623
transform 1 0 8624 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1694700623
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1839_
timestamp 1694700623
transform 1 0 8960 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1840_
timestamp 1694700623
transform 1 0 10080 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1841_
timestamp 1694700623
transform 1 0 12320 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1694700623
transform 1 0 10976 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1694700623
transform -1 0 13104 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1844_
timestamp 1694700623
transform -1 0 12320 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1845_
timestamp 1694700623
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1694700623
transform -1 0 9184 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1694700623
transform -1 0 8736 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1848_
timestamp 1694700623
transform 1 0 9072 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1849_
timestamp 1694700623
transform -1 0 10528 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1694700623
transform -1 0 9968 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1851_
timestamp 1694700623
transform -1 0 10304 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1852_
timestamp 1694700623
transform -1 0 8512 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1694700623
transform 1 0 8288 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1694700623
transform 1 0 6944 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1694700623
transform 1 0 8512 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1856_
timestamp 1694700623
transform -1 0 8736 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1694700623
transform 1 0 8736 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1858_
timestamp 1694700623
transform -1 0 11088 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1859_
timestamp 1694700623
transform -1 0 8960 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1860_
timestamp 1694700623
transform 1 0 7840 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1861_
timestamp 1694700623
transform -1 0 48384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1862_
timestamp 1694700623
transform -1 0 10864 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1694700623
transform -1 0 10304 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1864_
timestamp 1694700623
transform 1 0 10080 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1865_
timestamp 1694700623
transform 1 0 9968 0 1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1866_
timestamp 1694700623
transform -1 0 12208 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1694700623
transform 1 0 10640 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1694700623
transform -1 0 13552 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1869_
timestamp 1694700623
transform -1 0 12992 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1870_
timestamp 1694700623
transform -1 0 13440 0 -1 64288
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1694700623
transform 1 0 12432 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1872_
timestamp 1694700623
transform -1 0 14448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1694700623
transform -1 0 14000 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1874_
timestamp 1694700623
transform 1 0 12432 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1875_
timestamp 1694700623
transform 1 0 12768 0 -1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1876_
timestamp 1694700623
transform -1 0 17248 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1694700623
transform 1 0 14672 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1694700623
transform 1 0 16240 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1879_
timestamp 1694700623
transform 1 0 25312 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1880_
timestamp 1694700623
transform -1 0 38976 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1881_
timestamp 1694700623
transform 1 0 17248 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1882_
timestamp 1694700623
transform 1 0 17248 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1694700623
transform -1 0 57344 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1884_
timestamp 1694700623
transform 1 0 48720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1885_
timestamp 1694700623
transform 1 0 53760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1886_
timestamp 1694700623
transform -1 0 55440 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1887_
timestamp 1694700623
transform -1 0 53872 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1888_
timestamp 1694700623
transform 1 0 50400 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1694700623
transform -1 0 56224 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1890_
timestamp 1694700623
transform -1 0 57120 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1891_
timestamp 1694700623
transform 1 0 56448 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1892_
timestamp 1694700623
transform -1 0 54768 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1694700623
transform -1 0 55664 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1894_
timestamp 1694700623
transform 1 0 53312 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1694700623
transform 1 0 48608 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1896_
timestamp 1694700623
transform -1 0 52304 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1694700623
transform -1 0 51408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1694700623
transform 1 0 51408 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1694700623
transform 1 0 35392 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1900_
timestamp 1694700623
transform 1 0 49056 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1694700623
transform 1 0 51408 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1694700623
transform -1 0 50400 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1694700623
transform 1 0 50176 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1904_
timestamp 1694700623
transform -1 0 52192 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1694700623
transform -1 0 51520 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1906_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 37968 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1907_
timestamp 1694700623
transform 1 0 49280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1908_
timestamp 1694700623
transform 1 0 52752 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1909_
timestamp 1694700623
transform -1 0 53424 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1910_
timestamp 1694700623
transform -1 0 50960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1911_
timestamp 1694700623
transform -1 0 50400 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1912_
timestamp 1694700623
transform 1 0 49392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1913_
timestamp 1694700623
transform 1 0 51296 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1914_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 49168 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1694700623
transform 1 0 50064 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1694700623
transform 1 0 51632 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1917_
timestamp 1694700623
transform 1 0 52528 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1694700623
transform -1 0 53760 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1919_
timestamp 1694700623
transform 1 0 52528 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1920_
timestamp 1694700623
transform 1 0 50848 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1921_
timestamp 1694700623
transform 1 0 52976 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1922_
timestamp 1694700623
transform -1 0 53984 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1694700623
transform -1 0 52864 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1924_
timestamp 1694700623
transform 1 0 52528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1925_
timestamp 1694700623
transform -1 0 53984 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1694700623
transform -1 0 53088 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1694700623
transform 1 0 52528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1694700623
transform -1 0 53984 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1694700623
transform -1 0 53648 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1694700623
transform -1 0 53424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1694700623
transform 1 0 53872 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1694700623
transform 1 0 54992 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1933_
timestamp 1694700623
transform -1 0 57568 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1934_
timestamp 1694700623
transform 1 0 56448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1935_
timestamp 1694700623
transform 1 0 54432 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1936_
timestamp 1694700623
transform 1 0 54432 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1694700623
transform -1 0 58128 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1694700623
transform -1 0 57008 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1939_
timestamp 1694700623
transform 1 0 56448 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1694700623
transform 1 0 56448 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1694700623
transform -1 0 56896 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1942_
timestamp 1694700623
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1694700623
transform 1 0 57680 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1694700623
transform 1 0 57120 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1694700623
transform -1 0 57344 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1694700623
transform -1 0 57232 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1947_
timestamp 1694700623
transform 1 0 54656 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1694700623
transform 1 0 57344 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1949_
timestamp 1694700623
transform 1 0 54880 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1694700623
transform -1 0 57344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1694700623
transform 1 0 52976 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1694700623
transform -1 0 57344 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1694700623
transform -1 0 57232 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1954_
timestamp 1694700623
transform 1 0 56560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1694700623
transform 1 0 57568 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1694700623
transform 1 0 57008 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1694700623
transform -1 0 57456 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1694700623
transform -1 0 57008 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1694700623
transform -1 0 55216 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1960_
timestamp 1694700623
transform 1 0 54880 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1694700623
transform -1 0 54208 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1694700623
transform -1 0 52304 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1963_
timestamp 1694700623
transform -1 0 52304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1964_
timestamp 1694700623
transform -1 0 46816 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1694700623
transform 1 0 46256 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1966_
timestamp 1694700623
transform 1 0 50176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1967_
timestamp 1694700623
transform 1 0 48832 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1968_
timestamp 1694700623
transform -1 0 57568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1969_
timestamp 1694700623
transform 1 0 52528 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1694700623
transform -1 0 58016 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1694700623
transform -1 0 56224 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1972_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 54208 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1973_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 54768 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1974_
timestamp 1694700623
transform 1 0 42896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1975_
timestamp 1694700623
transform 1 0 45472 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1694700623
transform 1 0 47152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1977_
timestamp 1694700623
transform 1 0 49504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1978_
timestamp 1694700623
transform -1 0 57792 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1979_
timestamp 1694700623
transform -1 0 57904 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1980_
timestamp 1694700623
transform -1 0 42224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1981_
timestamp 1694700623
transform 1 0 26656 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1694700623
transform 1 0 38528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1983_
timestamp 1694700623
transform 1 0 42784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1984_
timestamp 1694700623
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1985_
timestamp 1694700623
transform 1 0 44688 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1986_
timestamp 1694700623
transform -1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1987_
timestamp 1694700623
transform -1 0 44352 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1988_
timestamp 1694700623
transform -1 0 44240 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1694700623
transform -1 0 43792 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1694700623
transform -1 0 43344 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1991_
timestamp 1694700623
transform -1 0 44464 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1992_
timestamp 1694700623
transform -1 0 44240 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1993_
timestamp 1694700623
transform 1 0 43792 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1694700623
transform 1 0 43792 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1694700623
transform -1 0 43792 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1996_
timestamp 1694700623
transform 1 0 41888 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1997_
timestamp 1694700623
transform -1 0 41888 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1998_
timestamp 1694700623
transform -1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1694700623
transform -1 0 44352 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2000_
timestamp 1694700623
transform 1 0 43904 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1694700623
transform -1 0 45248 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1694700623
transform -1 0 44240 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2003_
timestamp 1694700623
transform 1 0 45472 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2004_
timestamp 1694700623
transform 1 0 46816 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2005_
timestamp 1694700623
transform 1 0 45808 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2006_
timestamp 1694700623
transform -1 0 46256 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2007_
timestamp 1694700623
transform 1 0 46368 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2008_
timestamp 1694700623
transform -1 0 47712 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1694700623
transform 1 0 43120 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1694700623
transform 1 0 44912 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1694700623
transform 1 0 45584 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1694700623
transform -1 0 44464 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2013_
timestamp 1694700623
transform 1 0 45024 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2014_
timestamp 1694700623
transform -1 0 44912 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2015_
timestamp 1694700623
transform 1 0 31920 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2016_
timestamp 1694700623
transform 1 0 34496 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2017_
timestamp 1694700623
transform 1 0 33600 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2018_
timestamp 1694700623
transform -1 0 38304 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2019_
timestamp 1694700623
transform 1 0 31024 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2020_
timestamp 1694700623
transform 1 0 31696 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2021_
timestamp 1694700623
transform -1 0 32704 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2022_
timestamp 1694700623
transform 1 0 29008 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1694700623
transform 1 0 31584 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1694700623
transform 1 0 29232 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1694700623
transform 1 0 28448 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2026_
timestamp 1694700623
transform 1 0 29008 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2027_
timestamp 1694700623
transform 1 0 28224 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2028_
timestamp 1694700623
transform 1 0 29008 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2029_
timestamp 1694700623
transform -1 0 29680 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1694700623
transform 1 0 30352 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1694700623
transform 1 0 28224 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1694700623
transform 1 0 29680 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2033_
timestamp 1694700623
transform -1 0 30352 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1694700623
transform -1 0 28784 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2035_
timestamp 1694700623
transform -1 0 28560 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1694700623
transform 1 0 27552 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2037_
timestamp 1694700623
transform 1 0 26544 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2038_
timestamp 1694700623
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2039_
timestamp 1694700623
transform 1 0 28784 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2040_
timestamp 1694700623
transform -1 0 30576 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1694700623
transform 1 0 29232 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2042_
timestamp 1694700623
transform 1 0 31920 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1694700623
transform 1 0 29680 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1694700623
transform 1 0 30352 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2045_
timestamp 1694700623
transform -1 0 31024 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1694700623
transform 1 0 25984 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1694700623
transform 1 0 26880 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1694700623
transform 1 0 25984 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1694700623
transform -1 0 28336 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2050_
timestamp 1694700623
transform 1 0 27104 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2051_
timestamp 1694700623
transform 1 0 27328 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1694700623
transform -1 0 30688 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1694700623
transform -1 0 29904 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1694700623
transform 1 0 28784 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1694700623
transform 1 0 31024 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2056_
timestamp 1694700623
transform -1 0 31248 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2057_
timestamp 1694700623
transform 1 0 32816 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2058_
timestamp 1694700623
transform 1 0 32928 0 -1 64288
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2059_
timestamp 1694700623
transform -1 0 35280 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2060_
timestamp 1694700623
transform -1 0 32816 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2061_
timestamp 1694700623
transform -1 0 32704 0 1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2062_
timestamp 1694700623
transform -1 0 32704 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2063_
timestamp 1694700623
transform -1 0 23856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2064_
timestamp 1694700623
transform 1 0 49616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1694700623
transform -1 0 52416 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2066_
timestamp 1694700623
transform 1 0 41552 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2067_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 54208 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2068_
timestamp 1694700623
transform 1 0 46480 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2069_
timestamp 1694700623
transform -1 0 51856 0 1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2070_
timestamp 1694700623
transform -1 0 51744 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2071_
timestamp 1694700623
transform 1 0 50848 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2072_
timestamp 1694700623
transform 1 0 51408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1694700623
transform -1 0 28448 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2074_
timestamp 1694700623
transform 1 0 51184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1694700623
transform 1 0 50288 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2076_
timestamp 1694700623
transform 1 0 51184 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2077_
timestamp 1694700623
transform -1 0 37744 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2078_
timestamp 1694700623
transform 1 0 37744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2079_
timestamp 1694700623
transform 1 0 51296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 52080 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2081_
timestamp 1694700623
transform 1 0 54320 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2082_
timestamp 1694700623
transform 1 0 50400 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2083_
timestamp 1694700623
transform 1 0 53424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1694700623
transform -1 0 52304 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2085_
timestamp 1694700623
transform 1 0 52528 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1694700623
transform 1 0 54992 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2087_
timestamp 1694700623
transform -1 0 49504 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2088_
timestamp 1694700623
transform 1 0 49952 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2089_
timestamp 1694700623
transform -1 0 51856 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1694700623
transform -1 0 52752 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2091_
timestamp 1694700623
transform 1 0 43568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2092_
timestamp 1694700623
transform 1 0 52528 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2093_
timestamp 1694700623
transform 1 0 53984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2094_
timestamp 1694700623
transform -1 0 49616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2095_
timestamp 1694700623
transform -1 0 50960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2096_
timestamp 1694700623
transform 1 0 46704 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1694700623
transform -1 0 51072 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2098_
timestamp 1694700623
transform 1 0 50960 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2099_
timestamp 1694700623
transform 1 0 52528 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2100_
timestamp 1694700623
transform 1 0 49728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1694700623
transform -1 0 47376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2102_
timestamp 1694700623
transform -1 0 48272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2103_
timestamp 1694700623
transform -1 0 48048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2104_
timestamp 1694700623
transform -1 0 48384 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2105_
timestamp 1694700623
transform 1 0 47600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2106_
timestamp 1694700623
transform -1 0 45920 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2107_
timestamp 1694700623
transform 1 0 44912 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2108_
timestamp 1694700623
transform -1 0 45360 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1694700623
transform -1 0 45248 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1694700623
transform 1 0 43904 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2111_
timestamp 1694700623
transform 1 0 44688 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2112_
timestamp 1694700623
transform -1 0 44912 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2113_
timestamp 1694700623
transform -1 0 43008 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2114_
timestamp 1694700623
transform -1 0 42560 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2115_
timestamp 1694700623
transform 1 0 40768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2116_
timestamp 1694700623
transform 1 0 40880 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1694700623
transform 1 0 40768 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1694700623
transform 1 0 42448 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 41328 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2120_
timestamp 1694700623
transform -1 0 40432 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2121_
timestamp 1694700623
transform 1 0 38640 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2122_
timestamp 1694700623
transform 1 0 50512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2123_
timestamp 1694700623
transform -1 0 39760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2124_
timestamp 1694700623
transform 1 0 38640 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2125_
timestamp 1694700623
transform 1 0 39536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2126_
timestamp 1694700623
transform -1 0 38976 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1694700623
transform 1 0 38080 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2128_
timestamp 1694700623
transform -1 0 39424 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2129_
timestamp 1694700623
transform -1 0 37632 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2130_
timestamp 1694700623
transform 1 0 28560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2131_
timestamp 1694700623
transform 1 0 27664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1694700623
transform 1 0 51184 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2133_
timestamp 1694700623
transform 1 0 48160 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2134_
timestamp 1694700623
transform 1 0 35280 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2135_
timestamp 1694700623
transform -1 0 41664 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2136_
timestamp 1694700623
transform -1 0 50960 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2137_
timestamp 1694700623
transform 1 0 50624 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2138_
timestamp 1694700623
transform 1 0 52528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1694700623
transform 1 0 47264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2140_
timestamp 1694700623
transform 1 0 50960 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1694700623
transform -1 0 50624 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2142_
timestamp 1694700623
transform 1 0 42784 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2143_
timestamp 1694700623
transform 1 0 50400 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2144_
timestamp 1694700623
transform 1 0 52304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2145_
timestamp 1694700623
transform -1 0 49056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2146_
timestamp 1694700623
transform -1 0 50176 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1694700623
transform 1 0 49504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2148_
timestamp 1694700623
transform 1 0 50176 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1694700623
transform 1 0 51072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2150_
timestamp 1694700623
transform -1 0 39872 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2151_
timestamp 1694700623
transform -1 0 39760 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2152_
timestamp 1694700623
transform 1 0 39648 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2153_
timestamp 1694700623
transform -1 0 42000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2154_
timestamp 1694700623
transform -1 0 40432 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2155_
timestamp 1694700623
transform -1 0 41664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2156_
timestamp 1694700623
transform -1 0 41104 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2157_
timestamp 1694700623
transform 1 0 40544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1694700623
transform -1 0 37856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2159_
timestamp 1694700623
transform -1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2160_
timestamp 1694700623
transform 1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2161_
timestamp 1694700623
transform -1 0 39088 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2162_
timestamp 1694700623
transform 1 0 37968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1694700623
transform -1 0 35728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2164_
timestamp 1694700623
transform -1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2165_
timestamp 1694700623
transform 1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2166_
timestamp 1694700623
transform -1 0 36960 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2167_
timestamp 1694700623
transform -1 0 36288 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2168_
timestamp 1694700623
transform 1 0 35280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2169_
timestamp 1694700623
transform -1 0 34720 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2170_
timestamp 1694700623
transform 1 0 33152 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2171_
timestamp 1694700623
transform 1 0 33488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1694700623
transform 1 0 33376 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1694700623
transform -1 0 33152 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2174_
timestamp 1694700623
transform 1 0 33488 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2175_
timestamp 1694700623
transform -1 0 34048 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2176_
timestamp 1694700623
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1694700623
transform 1 0 31360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2178_
timestamp 1694700623
transform 1 0 32592 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2179_
timestamp 1694700623
transform -1 0 33600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1694700623
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2181_
timestamp 1694700623
transform -1 0 32704 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2182_
timestamp 1694700623
transform 1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2183_
timestamp 1694700623
transform 1 0 34720 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2184_
timestamp 1694700623
transform 1 0 34384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2185_
timestamp 1694700623
transform 1 0 34160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1694700623
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2187_
timestamp 1694700623
transform -1 0 42448 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2188_
timestamp 1694700623
transform -1 0 32928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2189_
timestamp 1694700623
transform 1 0 33600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2190_
timestamp 1694700623
transform 1 0 33376 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2191_
timestamp 1694700623
transform 1 0 35168 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2192_
timestamp 1694700623
transform 1 0 39200 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1694700623
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2194_
timestamp 1694700623
transform 1 0 8064 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2195_
timestamp 1694700623
transform -1 0 28000 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2196_
timestamp 1694700623
transform 1 0 23520 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2197_
timestamp 1694700623
transform 1 0 18592 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2198_
timestamp 1694700623
transform 1 0 23184 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2199_
timestamp 1694700623
transform 1 0 27328 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1694700623
transform 1 0 26768 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1694700623
transform -1 0 27440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1694700623
transform -1 0 27776 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2203_
timestamp 1694700623
transform 1 0 26544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2204_
timestamp 1694700623
transform -1 0 26544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2205_
timestamp 1694700623
transform 1 0 26544 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2206_
timestamp 1694700623
transform -1 0 27104 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1694700623
transform -1 0 26320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2208_
timestamp 1694700623
transform -1 0 25536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2209_
timestamp 1694700623
transform -1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1694700623
transform -1 0 24528 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2211_
timestamp 1694700623
transform 1 0 23408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2212_
timestamp 1694700623
transform 1 0 23296 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2213_
timestamp 1694700623
transform -1 0 23408 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2214_
timestamp 1694700623
transform -1 0 22624 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2215_
timestamp 1694700623
transform 1 0 21392 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2216_
timestamp 1694700623
transform -1 0 21504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1694700623
transform -1 0 20944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1694700623
transform -1 0 21952 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2219_
timestamp 1694700623
transform 1 0 21168 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2220_
timestamp 1694700623
transform -1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2221_
timestamp 1694700623
transform -1 0 19488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2222_
timestamp 1694700623
transform -1 0 20384 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2223_
timestamp 1694700623
transform 1 0 18704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2224_
timestamp 1694700623
transform -1 0 19824 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2225_
timestamp 1694700623
transform -1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2226_
timestamp 1694700623
transform -1 0 18592 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2227_
timestamp 1694700623
transform -1 0 18368 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2228_
timestamp 1694700623
transform 1 0 18592 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2229_
timestamp 1694700623
transform -1 0 19712 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2230_
timestamp 1694700623
transform -1 0 16128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2231_
timestamp 1694700623
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2232_
timestamp 1694700623
transform -1 0 19040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1694700623
transform 1 0 19040 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1694700623
transform -1 0 18144 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2235_
timestamp 1694700623
transform 1 0 19712 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2236_
timestamp 1694700623
transform -1 0 19824 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2237_
timestamp 1694700623
transform -1 0 16128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2238_
timestamp 1694700623
transform 1 0 20272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2239_
timestamp 1694700623
transform 1 0 18144 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2240_
timestamp 1694700623
transform -1 0 20720 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1694700623
transform 1 0 21168 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2242_
timestamp 1694700623
transform -1 0 19152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2243_
timestamp 1694700623
transform -1 0 21952 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2244_
timestamp 1694700623
transform 1 0 22400 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2245_
timestamp 1694700623
transform 1 0 23296 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2246_
timestamp 1694700623
transform 1 0 23184 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1694700623
transform 1 0 22288 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1694700623
transform 1 0 24080 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2249_
timestamp 1694700623
transform -1 0 22624 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2250_
timestamp 1694700623
transform 1 0 22624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2251_
timestamp 1694700623
transform 1 0 22960 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1694700623
transform 1 0 24304 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1694700623
transform 1 0 19264 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2254_
timestamp 1694700623
transform 1 0 18368 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2255_
timestamp 1694700623
transform 1 0 36288 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2256_
timestamp 1694700623
transform -1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2257_
timestamp 1694700623
transform 1 0 46368 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1694700623
transform -1 0 45920 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 34384 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2260_
timestamp 1694700623
transform -1 0 36064 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2261_
timestamp 1694700623
transform 1 0 37968 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2262_
timestamp 1694700623
transform -1 0 44464 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2263_
timestamp 1694700623
transform -1 0 41888 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2264_
timestamp 1694700623
transform 1 0 43344 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1694700623
transform 1 0 43792 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2266_
timestamp 1694700623
transform 1 0 44688 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2267_
timestamp 1694700623
transform 1 0 36848 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1694700623
transform 1 0 44240 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2269_
timestamp 1694700623
transform 1 0 45584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2270_
timestamp 1694700623
transform -1 0 45696 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1694700623
transform -1 0 43344 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2272_
timestamp 1694700623
transform 1 0 43120 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1694700623
transform 1 0 42224 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2274_
timestamp 1694700623
transform 1 0 36848 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2275_
timestamp 1694700623
transform -1 0 43456 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2276_
timestamp 1694700623
transform -1 0 41440 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2277_
timestamp 1694700623
transform 1 0 41440 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2278_
timestamp 1694700623
transform -1 0 42336 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2279_
timestamp 1694700623
transform 1 0 36960 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2280_
timestamp 1694700623
transform 1 0 41664 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2281_
timestamp 1694700623
transform -1 0 42560 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2282_
timestamp 1694700623
transform -1 0 41664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1694700623
transform 1 0 41440 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2284_
timestamp 1694700623
transform -1 0 41440 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2285_
timestamp 1694700623
transform 1 0 40768 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2286_
timestamp 1694700623
transform -1 0 41888 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2287_
timestamp 1694700623
transform -1 0 42000 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2288_
timestamp 1694700623
transform 1 0 38976 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1694700623
transform 1 0 39648 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2290_
timestamp 1694700623
transform 1 0 39312 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2291_
timestamp 1694700623
transform -1 0 49280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2292_
timestamp 1694700623
transform 1 0 42224 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1694700623
transform 1 0 42672 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2294_
timestamp 1694700623
transform 1 0 41216 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2295_
timestamp 1694700623
transform 1 0 43120 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2296_
timestamp 1694700623
transform 1 0 42784 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2297_
timestamp 1694700623
transform 1 0 44800 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1694700623
transform -1 0 43456 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2299_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 43120 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2300_
timestamp 1694700623
transform 1 0 42784 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2301_
timestamp 1694700623
transform 1 0 41216 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2302_
timestamp 1694700623
transform 1 0 39200 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1694700623
transform -1 0 41104 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2304_
timestamp 1694700623
transform 1 0 40768 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1694700623
transform -1 0 43008 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2306_
timestamp 1694700623
transform -1 0 42784 0 -1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2307_
timestamp 1694700623
transform -1 0 43904 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2308_
timestamp 1694700623
transform 1 0 40208 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2309_
timestamp 1694700623
transform 1 0 42112 0 -1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2310_
timestamp 1694700623
transform 1 0 42896 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1694700623
transform -1 0 47040 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1694700623
transform 1 0 43904 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1694700623
transform -1 0 44352 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1694700623
transform 1 0 44464 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2315_
timestamp 1694700623
transform -1 0 45920 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2316_
timestamp 1694700623
transform 1 0 45920 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2317_
timestamp 1694700623
transform -1 0 45696 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2318_
timestamp 1694700623
transform -1 0 47488 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2319_
timestamp 1694700623
transform -1 0 47264 0 -1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2320_
timestamp 1694700623
transform 1 0 52528 0 1 61152
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1694700623
transform 1 0 55440 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2322_
timestamp 1694700623
transform 1 0 53760 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2323_
timestamp 1694700623
transform 1 0 52864 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2324_
timestamp 1694700623
transform -1 0 54992 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2325_
timestamp 1694700623
transform 1 0 53648 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2326_
timestamp 1694700623
transform 1 0 56448 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1694700623
transform 1 0 56448 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1694700623
transform 1 0 57568 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2329_
timestamp 1694700623
transform 1 0 56448 0 -1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2330_
timestamp 1694700623
transform 1 0 52304 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2331_
timestamp 1694700623
transform -1 0 53200 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2332_
timestamp 1694700623
transform 1 0 51408 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2333_
timestamp 1694700623
transform 1 0 53984 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2334_
timestamp 1694700623
transform -1 0 55104 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2335_
timestamp 1694700623
transform -1 0 56224 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2336_
timestamp 1694700623
transform 1 0 56448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2337_
timestamp 1694700623
transform 1 0 54992 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2338_
timestamp 1694700623
transform -1 0 56560 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2339_
timestamp 1694700623
transform 1 0 54544 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1694700623
transform -1 0 55776 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2341_
timestamp 1694700623
transform 1 0 56448 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2342_
timestamp 1694700623
transform -1 0 56224 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2343_
timestamp 1694700623
transform -1 0 51296 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2344_
timestamp 1694700623
transform 1 0 50736 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2345_
timestamp 1694700623
transform -1 0 52752 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2346_
timestamp 1694700623
transform -1 0 55328 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2347_
timestamp 1694700623
transform -1 0 54768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2348_
timestamp 1694700623
transform -1 0 53424 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2349_
timestamp 1694700623
transform -1 0 49728 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2350_
timestamp 1694700623
transform 1 0 46592 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2351_
timestamp 1694700623
transform 1 0 47152 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2352_
timestamp 1694700623
transform 1 0 38976 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2353_
timestamp 1694700623
transform -1 0 47488 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1694700623
transform 1 0 44688 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1694700623
transform 1 0 51184 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2356_
timestamp 1694700623
transform 1 0 50736 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 46816 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1694700623
transform 1 0 48608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2359_
timestamp 1694700623
transform -1 0 47264 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2360_
timestamp 1694700623
transform 1 0 43008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1694700623
transform -1 0 50512 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2362_
timestamp 1694700623
transform 1 0 45696 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2363_
timestamp 1694700623
transform 1 0 45360 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2364_
timestamp 1694700623
transform 1 0 46704 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2365_
timestamp 1694700623
transform 1 0 48608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2366_
timestamp 1694700623
transform -1 0 51520 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2367_
timestamp 1694700623
transform -1 0 50736 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2368_
timestamp 1694700623
transform 1 0 48608 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2369_
timestamp 1694700623
transform -1 0 48384 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2370_
timestamp 1694700623
transform 1 0 48720 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2371_
timestamp 1694700623
transform 1 0 48944 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2372_
timestamp 1694700623
transform 1 0 49280 0 -1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2373_
timestamp 1694700623
transform -1 0 50512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2374_
timestamp 1694700623
transform 1 0 50400 0 1 62720
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2375_
timestamp 1694700623
transform 1 0 51520 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2376_
timestamp 1694700623
transform 1 0 50736 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2377_
timestamp 1694700623
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1694700623
transform -1 0 53536 0 1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2379_
timestamp 1694700623
transform 1 0 51296 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2380_
timestamp 1694700623
transform 1 0 50176 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2381_
timestamp 1694700623
transform -1 0 31808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2382_
timestamp 1694700623
transform 1 0 31248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2383_
timestamp 1694700623
transform -1 0 24640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2384_
timestamp 1694700623
transform -1 0 23744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2385_
timestamp 1694700623
transform 1 0 22512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2386_
timestamp 1694700623
transform -1 0 27552 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2387_
timestamp 1694700623
transform 1 0 24640 0 1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2388_
timestamp 1694700623
transform 1 0 36624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2389_
timestamp 1694700623
transform 1 0 33488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1694700623
transform 1 0 41888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1694700623
transform 1 0 41104 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2392_
timestamp 1694700623
transform -1 0 24528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2393_
timestamp 1694700623
transform 1 0 34496 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2394_
timestamp 1694700623
transform -1 0 42448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2395_
timestamp 1694700623
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2396_
timestamp 1694700623
transform -1 0 36624 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1694700623
transform 1 0 41104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2398_
timestamp 1694700623
transform 1 0 42000 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1694700623
transform 1 0 39424 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2400_
timestamp 1694700623
transform 1 0 38640 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2401_
timestamp 1694700623
transform -1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2402_
timestamp 1694700623
transform 1 0 37744 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2403_
timestamp 1694700623
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2404_
timestamp 1694700623
transform -1 0 34384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1694700623
transform -1 0 33936 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2406_
timestamp 1694700623
transform 1 0 33376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2407_
timestamp 1694700623
transform -1 0 35952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2408_
timestamp 1694700623
transform 1 0 34160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2409_
timestamp 1694700623
transform -1 0 26096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2410_
timestamp 1694700623
transform -1 0 27888 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2411_
timestamp 1694700623
transform -1 0 27104 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2412_
timestamp 1694700623
transform 1 0 26320 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2413_
timestamp 1694700623
transform 1 0 27776 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2414_
timestamp 1694700623
transform 1 0 29120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1694700623
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2416_
timestamp 1694700623
transform 1 0 34832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2417_
timestamp 1694700623
transform 1 0 28560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1694700623
transform 1 0 27664 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2419_
timestamp 1694700623
transform 1 0 19600 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2420_
timestamp 1694700623
transform 1 0 26992 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2421_
timestamp 1694700623
transform 1 0 29792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2422_
timestamp 1694700623
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2423_
timestamp 1694700623
transform 1 0 18704 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2424_
timestamp 1694700623
transform 1 0 23968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2425_
timestamp 1694700623
transform 1 0 28336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2426_
timestamp 1694700623
transform 1 0 26432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2427_
timestamp 1694700623
transform 1 0 31360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2428_
timestamp 1694700623
transform 1 0 30464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1694700623
transform 1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2430_
timestamp 1694700623
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2431_
timestamp 1694700623
transform 1 0 25088 0 -1 21952
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1694700623
transform -1 0 18816 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2433_
timestamp 1694700623
transform -1 0 19488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2434_
timestamp 1694700623
transform 1 0 19040 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2435_
timestamp 1694700623
transform 1 0 18368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2436_
timestamp 1694700623
transform -1 0 23296 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2437_
timestamp 1694700623
transform 1 0 18144 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2438_
timestamp 1694700623
transform 1 0 17248 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1694700623
transform -1 0 20160 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2440_
timestamp 1694700623
transform 1 0 18256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2441_
timestamp 1694700623
transform 1 0 18144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2442_
timestamp 1694700623
transform 1 0 18144 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2443_
timestamp 1694700623
transform 1 0 17808 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1694700623
transform 1 0 21616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2445_
timestamp 1694700623
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2446_
timestamp 1694700623
transform -1 0 35952 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2447_
timestamp 1694700623
transform 1 0 21728 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2448_
timestamp 1694700623
transform 1 0 20048 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2449_
timestamp 1694700623
transform -1 0 31472 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2450_
timestamp 1694700623
transform 1 0 24416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1694700623
transform -1 0 32928 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1694700623
transform -1 0 28784 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2453_
timestamp 1694700623
transform 1 0 25088 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2454_
timestamp 1694700623
transform 1 0 25760 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1694700623
transform 1 0 26432 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2456_
timestamp 1694700623
transform 1 0 28000 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1694700623
transform 1 0 27888 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2458_
timestamp 1694700623
transform 1 0 30464 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2459_
timestamp 1694700623
transform 1 0 30688 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1694700623
transform 1 0 31136 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1694700623
transform -1 0 25760 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2462_
timestamp 1694700623
transform 1 0 30464 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1694700623
transform -1 0 30688 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2464_
timestamp 1694700623
transform -1 0 30128 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2465_
timestamp 1694700623
transform -1 0 29008 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2466_
timestamp 1694700623
transform -1 0 28224 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1694700623
transform -1 0 33488 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1694700623
transform 1 0 25088 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2469_
timestamp 1694700623
transform 1 0 25424 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1694700623
transform -1 0 24864 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1694700623
transform -1 0 24864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2472_
timestamp 1694700623
transform -1 0 24192 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1694700623
transform 1 0 23856 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2474_
timestamp 1694700623
transform 1 0 24080 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1694700623
transform -1 0 23632 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1694700623
transform -1 0 23408 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2477_
timestamp 1694700623
transform -1 0 22512 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1694700623
transform -1 0 23072 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2479_
timestamp 1694700623
transform -1 0 22512 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1694700623
transform -1 0 22624 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2481_
timestamp 1694700623
transform -1 0 22064 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1694700623
transform -1 0 29344 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2483_
timestamp 1694700623
transform -1 0 26432 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2484_
timestamp 1694700623
transform -1 0 25648 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2485_
timestamp 1694700623
transform -1 0 16128 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2486_
timestamp 1694700623
transform 1 0 13328 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2487_
timestamp 1694700623
transform 1 0 14672 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2488_
timestamp 1694700623
transform 1 0 14448 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2489_
timestamp 1694700623
transform -1 0 14672 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1694700623
transform -1 0 19376 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2491_
timestamp 1694700623
transform 1 0 13776 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2492_
timestamp 1694700623
transform 1 0 14000 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2493_
timestamp 1694700623
transform 1 0 13776 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1694700623
transform -1 0 15120 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2495_
timestamp 1694700623
transform 1 0 13776 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2496_
timestamp 1694700623
transform -1 0 28000 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1694700623
transform -1 0 24416 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1694700623
transform -1 0 17024 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2499_
timestamp 1694700623
transform -1 0 17920 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1694700623
transform -1 0 17808 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2501_
timestamp 1694700623
transform -1 0 17024 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1694700623
transform 1 0 17920 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2503_
timestamp 1694700623
transform -1 0 36064 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2504_
timestamp 1694700623
transform 1 0 17248 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2505_
timestamp 1694700623
transform 1 0 16016 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2506_
timestamp 1694700623
transform 1 0 17248 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1694700623
transform 1 0 16128 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2508_
timestamp 1694700623
transform 1 0 15904 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1694700623
transform 1 0 27776 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1694700623
transform 1 0 22064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1694700623
transform 1 0 21280 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1694700623
transform -1 0 24528 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2513_
timestamp 1694700623
transform 1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2514_
timestamp 1694700623
transform 1 0 28560 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1694700623
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2516_
timestamp 1694700623
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2517_
timestamp 1694700623
transform 1 0 38976 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2518_
timestamp 1694700623
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2519_
timestamp 1694700623
transform -1 0 38640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2520_
timestamp 1694700623
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2521_
timestamp 1694700623
transform -1 0 38192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2522_
timestamp 1694700623
transform -1 0 37520 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2523_
timestamp 1694700623
transform -1 0 40432 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1694700623
transform 1 0 37968 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2525_
timestamp 1694700623
transform 1 0 38528 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2526_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 38304 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2527_
timestamp 1694700623
transform -1 0 30576 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2528_
timestamp 1694700623
transform -1 0 30800 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2529_
timestamp 1694700623
transform -1 0 30688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2530_
timestamp 1694700623
transform -1 0 32480 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2531_
timestamp 1694700623
transform 1 0 46816 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2532_
timestamp 1694700623
transform 1 0 44576 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2533_
timestamp 1694700623
transform 1 0 44016 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2534_
timestamp 1694700623
transform -1 0 44688 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2535_
timestamp 1694700623
transform 1 0 47712 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2536_
timestamp 1694700623
transform 1 0 46928 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2537_
timestamp 1694700623
transform 1 0 44912 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2538_
timestamp 1694700623
transform 1 0 45136 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2539_
timestamp 1694700623
transform -1 0 43232 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2540_
timestamp 1694700623
transform -1 0 44016 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2541_
timestamp 1694700623
transform 1 0 18816 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2542_
timestamp 1694700623
transform 1 0 22736 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2543_
timestamp 1694700623
transform 1 0 16464 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2544_
timestamp 1694700623
transform 1 0 17248 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2545_
timestamp 1694700623
transform 1 0 20496 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2546_
timestamp 1694700623
transform 1 0 21168 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2547_
timestamp 1694700623
transform 1 0 21504 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2548_
timestamp 1694700623
transform 1 0 16352 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2549_
timestamp 1694700623
transform 1 0 19936 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2550_
timestamp 1694700623
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2551_
timestamp 1694700623
transform 1 0 1568 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2552_
timestamp 1694700623
transform 1 0 1568 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2553_
timestamp 1694700623
transform 1 0 1568 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2554_
timestamp 1694700623
transform 1 0 1568 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2555_
timestamp 1694700623
transform 1 0 1568 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2556_
timestamp 1694700623
transform 1 0 1568 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2557_
timestamp 1694700623
transform 1 0 2576 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2558_
timestamp 1694700623
transform 1 0 5488 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2559_
timestamp 1694700623
transform -1 0 21952 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2560_
timestamp 1694700623
transform 1 0 17696 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2561_
timestamp 1694700623
transform 1 0 4368 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2562_
timestamp 1694700623
transform 1 0 5152 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2563_
timestamp 1694700623
transform 1 0 5824 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2564_
timestamp 1694700623
transform -1 0 13104 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2565_
timestamp 1694700623
transform 1 0 5824 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2566_
timestamp 1694700623
transform 1 0 5040 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2567_
timestamp 1694700623
transform 1 0 6496 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2568_
timestamp 1694700623
transform 1 0 8176 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_
timestamp 1694700623
transform 1 0 9184 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1694700623
transform 1 0 13328 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1694700623
transform -1 0 20496 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1694700623
transform 1 0 53424 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 52528 0 1 47040
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1694700623
transform -1 0 58352 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1694700623
transform 1 0 52864 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1694700623
transform 1 0 49840 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1694700623
transform 1 0 48944 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1694700623
transform 1 0 50064 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1694700623
transform -1 0 48496 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1694700623
transform -1 0 50064 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1694700623
transform 1 0 51184 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1694700623
transform 1 0 49280 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1694700623
transform 1 0 50512 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1694700623
transform -1 0 55328 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1694700623
transform 1 0 55104 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1694700623
transform -1 0 58240 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1694700623
transform 1 0 55104 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1694700623
transform 1 0 55104 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1694700623
transform 1 0 55104 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1694700623
transform 1 0 55104 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1694700623
transform 1 0 53088 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1694700623
transform 1 0 52528 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1694700623
transform 1 0 48160 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1694700623
transform -1 0 50064 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1694700623
transform 1 0 42336 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1694700623
transform 1 0 40880 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1694700623
transform 1 0 42112 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1694700623
transform 1 0 38640 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1694700623
transform -1 0 45808 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1694700623
transform -1 0 49168 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1694700623
transform -1 0 49504 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1694700623
transform 1 0 44912 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1694700623
transform -1 0 36400 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1694700623
transform -1 0 34160 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1694700623
transform 1 0 25312 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1694700623
transform 1 0 25088 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1694700623
transform -1 0 34720 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1694700623
transform 1 0 23856 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1694700623
transform 1 0 27888 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1694700623
transform -1 0 36624 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1694700623
transform 1 0 21616 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2612_
timestamp 1694700623
transform -1 0 55776 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1694700623
transform -1 0 57456 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1694700623
transform -1 0 58352 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1694700623
transform -1 0 57456 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1694700623
transform -1 0 56224 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1694700623
transform -1 0 49840 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1694700623
transform 1 0 43008 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1694700623
transform 1 0 41664 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2620_
timestamp 1694700623
transform 1 0 39312 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1694700623
transform 1 0 37632 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1694700623
transform -1 0 28560 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1694700623
transform -1 0 55440 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1694700623
transform -1 0 55776 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1694700623
transform -1 0 53648 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1694700623
transform 1 0 40768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1694700623
transform -1 0 40096 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1694700623
transform -1 0 37408 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1694700623
transform 1 0 32592 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1694700623
transform 1 0 29344 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1694700623
transform 1 0 35056 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1694700623
transform 1 0 34832 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2633_
timestamp 1694700623
transform 1 0 5824 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1694700623
transform -1 0 27776 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1694700623
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2636_
timestamp 1694700623
transform 1 0 21504 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1694700623
transform 1 0 18256 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1694700623
transform 1 0 15232 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1694700623
transform 1 0 13776 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1694700623
transform 1 0 14224 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1694700623
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1694700623
transform -1 0 24752 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1694700623
transform 1 0 23408 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2644_
timestamp 1694700623
transform 1 0 15008 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1694700623
transform 1 0 45136 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1694700623
transform 1 0 40544 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1694700623
transform 1 0 44688 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1694700623
transform 1 0 38640 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1694700623
transform -1 0 41664 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1694700623
transform 1 0 37408 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1694700623
transform -1 0 47936 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1694700623
transform 1 0 38304 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1694700623
transform -1 0 44688 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1694700623
transform 1 0 44688 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1694700623
transform -1 0 58352 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1694700623
transform -1 0 58352 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2657_
timestamp 1694700623
transform -1 0 58352 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1694700623
transform 1 0 50624 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1694700623
transform 1 0 55104 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2660_
timestamp 1694700623
transform 1 0 55104 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1694700623
transform 1 0 54656 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1694700623
transform 1 0 55104 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1694700623
transform 1 0 36512 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1694700623
transform -1 0 53984 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1694700623
transform -1 0 49840 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1694700623
transform 1 0 43456 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1694700623
transform -1 0 50736 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1694700623
transform 1 0 42336 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1694700623
transform 1 0 44688 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1694700623
transform -1 0 50176 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1694700623
transform 1 0 46816 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1694700623
transform 1 0 48608 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1694700623
transform 1 0 48608 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1694700623
transform -1 0 55104 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1694700623
transform 1 0 51184 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1694700623
transform 1 0 50736 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1694700623
transform 1 0 49056 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1694700623
transform 1 0 41104 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1694700623
transform 1 0 41664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1694700623
transform 1 0 41216 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1694700623
transform 1 0 37632 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1694700623
transform 1 0 35056 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1694700623
transform 1 0 33376 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1694700623
transform 1 0 26432 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1694700623
transform 1 0 26992 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1694700623
transform 1 0 27664 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1694700623
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1694700623
transform 1 0 29456 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1694700623
transform 1 0 30464 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2690_
timestamp 1694700623
transform 1 0 15680 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1694700623
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1694700623
transform 1 0 14896 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1694700623
transform 1 0 14224 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1694700623
transform 1 0 19712 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1694700623
transform 1 0 19264 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1694700623
transform 1 0 30800 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1694700623
transform 1 0 31024 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2698_
timestamp 1694700623
transform 1 0 27888 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1694700623
transform 1 0 25536 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1694700623
transform 1 0 23744 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1694700623
transform 1 0 21168 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1694700623
transform 1 0 21168 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1694700623
transform 1 0 19376 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1694700623
transform 1 0 4144 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1694700623
transform 1 0 4592 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2706_
timestamp 1694700623
transform -1 0 12544 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1694700623
transform 1 0 9856 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1694700623
transform 1 0 15232 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2709_
timestamp 1694700623
transform 1 0 16688 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2710_
timestamp 1694700623
transform 1 0 16576 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2711_
timestamp 1694700623
transform -1 0 17024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1694700623
transform 1 0 19600 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1694700623
transform 1 0 21504 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1694700623
transform -1 0 31024 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1694700623
transform 1 0 45472 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1694700623
transform 1 0 35168 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1694700623
transform 1 0 36848 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1694700623
transform 1 0 38416 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A3 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 36176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A1
timestamp 1694700623
transform 1 0 34832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A3
timestamp 1694700623
transform 1 0 34720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__A1
timestamp 1694700623
transform 1 0 38752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A1
timestamp 1694700623
transform -1 0 33264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1694700623
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A1
timestamp 1694700623
transform 1 0 21392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A3
timestamp 1694700623
transform 1 0 14000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A2
timestamp 1694700623
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1694700623
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__A1
timestamp 1694700623
transform -1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A3
timestamp 1694700623
transform -1 0 31136 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A1
timestamp 1694700623
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A1
timestamp 1694700623
transform 1 0 20944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A1
timestamp 1694700623
transform 1 0 21392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I
timestamp 1694700623
transform 1 0 29120 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1694700623
transform 1 0 12320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1694700623
transform 1 0 33712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1694700623
transform -1 0 32592 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1694700623
transform 1 0 13664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1694700623
transform -1 0 13776 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A2
timestamp 1694700623
transform -1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1694700623
transform 1 0 31920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1694700623
transform 1 0 12768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1694700623
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A2
timestamp 1694700623
transform -1 0 32592 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__I
timestamp 1694700623
transform -1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A2
timestamp 1694700623
transform -1 0 32592 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1694700623
transform 1 0 14560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1694700623
transform 1 0 13552 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__I
timestamp 1694700623
transform 1 0 11760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__I
timestamp 1694700623
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A1
timestamp 1694700623
transform -1 0 30240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1694700623
transform 1 0 27664 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__I
timestamp 1694700623
transform -1 0 26656 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__I
timestamp 1694700623
transform 1 0 30464 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1694700623
transform 1 0 27440 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__I
timestamp 1694700623
transform 1 0 27776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1694700623
transform 1 0 10752 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__I
timestamp 1694700623
transform 1 0 10752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A2
timestamp 1694700623
transform -1 0 14000 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1694700623
transform 1 0 32256 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A2
timestamp 1694700623
transform 1 0 33600 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1694700623
transform 1 0 15792 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__I
timestamp 1694700623
transform 1 0 15344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__I
timestamp 1694700623
transform 1 0 14224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A2
timestamp 1694700623
transform 1 0 13328 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1694700623
transform 1 0 31584 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__I
timestamp 1694700623
transform 1 0 30912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1694700623
transform -1 0 37408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1694700623
transform 1 0 38640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A1
timestamp 1694700623
transform 1 0 50400 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1694700623
transform 1 0 36176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1694700623
transform 1 0 41888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1694700623
transform 1 0 29792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1694700623
transform 1 0 28112 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1694700623
transform -1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1694700623
transform 1 0 31696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1694700623
transform 1 0 35056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__C
timestamp 1694700623
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1694700623
transform -1 0 36064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1694700623
transform 1 0 35392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__I
timestamp 1694700623
transform 1 0 21280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1694700623
transform -1 0 23072 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__I
timestamp 1694700623
transform -1 0 42000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__B
timestamp 1694700623
transform 1 0 32480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1694700623
transform -1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__I
timestamp 1694700623
transform 1 0 34384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1694700623
transform 1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B
timestamp 1694700623
transform -1 0 30240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1694700623
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1694700623
transform -1 0 43456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__B
timestamp 1694700623
transform 1 0 32256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1694700623
transform -1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1694700623
transform -1 0 39088 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1694700623
transform 1 0 46816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__C
timestamp 1694700623
transform 1 0 46368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__B
timestamp 1694700623
transform 1 0 45808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1694700623
transform 1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1694700623
transform 1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__B
timestamp 1694700623
transform 1 0 45472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1694700623
transform 1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B
timestamp 1694700623
transform 1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1694700623
transform 1 0 43904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1694700623
transform 1 0 30800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1694700623
transform 1 0 47824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__C
timestamp 1694700623
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__B
timestamp 1694700623
transform 1 0 46592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1694700623
transform 1 0 46256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__B
timestamp 1694700623
transform -1 0 47376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1694700623
transform 1 0 45248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__I
timestamp 1694700623
transform -1 0 22288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__B
timestamp 1694700623
transform 1 0 45136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1694700623
transform 1 0 45360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B
timestamp 1694700623
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1694700623
transform 1 0 49728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1694700623
transform 1 0 49728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1694700623
transform 1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1694700623
transform 1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__B
timestamp 1694700623
transform 1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A1
timestamp 1694700623
transform 1 0 23184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__I
timestamp 1694700623
transform 1 0 49952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__I
timestamp 1694700623
transform -1 0 25536 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__B
timestamp 1694700623
transform -1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__B
timestamp 1694700623
transform 1 0 20944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B
timestamp 1694700623
transform 1 0 18256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__I
timestamp 1694700623
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1694700623
transform 1 0 18368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__B
timestamp 1694700623
transform 1 0 20720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B
timestamp 1694700623
transform 1 0 4480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1694700623
transform 1 0 3248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1694700623
transform 1 0 3024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1694700623
transform 1 0 2912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__B
timestamp 1694700623
transform 1 0 4592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__B
timestamp 1694700623
transform 1 0 4480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__B
timestamp 1694700623
transform 1 0 5040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I
timestamp 1694700623
transform 1 0 21392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1694700623
transform 1 0 8176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__B
timestamp 1694700623
transform 1 0 7504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1694700623
transform 1 0 20720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__I
timestamp 1694700623
transform 1 0 41776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__B
timestamp 1694700623
transform 1 0 20832 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B
timestamp 1694700623
transform 1 0 6832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1694700623
transform 1 0 8400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1694700623
transform 1 0 12992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1694700623
transform -1 0 48608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1694700623
transform 1 0 12208 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1694700623
transform -1 0 13328 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1694700623
transform 1 0 15568 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__I
timestamp 1694700623
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B
timestamp 1694700623
transform -1 0 18592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1694700623
transform 1 0 53536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1694700623
transform 1 0 52976 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1694700623
transform 1 0 55104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1694700623
transform 1 0 53088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__I
timestamp 1694700623
transform -1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A1
timestamp 1694700623
transform -1 0 50736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__I
timestamp 1694700623
transform 1 0 48832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A1
timestamp 1694700623
transform 1 0 49616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A1
timestamp 1694700623
transform 1 0 50624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1694700623
transform -1 0 50736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1694700623
transform -1 0 49168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__I
timestamp 1694700623
transform 1 0 57568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1694700623
transform 1 0 58128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1694700623
transform 1 0 58128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1694700623
transform 1 0 44800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1694700623
transform 1 0 45248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1694700623
transform -1 0 48272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1694700623
transform 1 0 57792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__I
timestamp 1694700623
transform -1 0 41552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__I
timestamp 1694700623
transform 1 0 27552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__I
timestamp 1694700623
transform 1 0 37856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1694700623
transform -1 0 44016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A3
timestamp 1694700623
transform -1 0 45920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1694700623
transform 1 0 44352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1694700623
transform 1 0 42672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__I
timestamp 1694700623
transform 1 0 43568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1694700623
transform 1 0 44912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__B
timestamp 1694700623
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1694700623
transform 1 0 45472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1694700623
transform 1 0 47712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__B
timestamp 1694700623
transform -1 0 45360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1694700623
transform 1 0 44464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__B
timestamp 1694700623
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__I
timestamp 1694700623
transform -1 0 38528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1694700623
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__B
timestamp 1694700623
transform 1 0 30464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__B
timestamp 1694700623
transform 1 0 28448 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1694700623
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__B
timestamp 1694700623
transform 1 0 28560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1694700623
transform 1 0 31248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B
timestamp 1694700623
transform -1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1694700623
transform 1 0 30800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1694700623
transform 1 0 31472 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1694700623
transform 1 0 35504 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__C
timestamp 1694700623
transform 1 0 32928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__I
timestamp 1694700623
transform -1 0 50736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1694700623
transform 1 0 52640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1694700623
transform 1 0 50624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__B
timestamp 1694700623
transform 1 0 51968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__I
timestamp 1694700623
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__I
timestamp 1694700623
transform -1 0 51184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__I
timestamp 1694700623
transform -1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__I
timestamp 1694700623
transform 1 0 37520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B
timestamp 1694700623
transform -1 0 51296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__C
timestamp 1694700623
transform 1 0 52752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__B
timestamp 1694700623
transform 1 0 51184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__C
timestamp 1694700623
transform -1 0 52752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__B
timestamp 1694700623
transform 1 0 52080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__I
timestamp 1694700623
transform 1 0 43344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__I
timestamp 1694700623
transform 1 0 49504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A1
timestamp 1694700623
transform 1 0 43680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__I
timestamp 1694700623
transform 1 0 42784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1694700623
transform 1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A2
timestamp 1694700623
transform 1 0 43680 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1694700623
transform 1 0 43232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A1
timestamp 1694700623
transform 1 0 38416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__I
timestamp 1694700623
transform 1 0 51408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A1
timestamp 1694700623
transform 1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1694700623
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__B
timestamp 1694700623
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1694700623
transform -1 0 38080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A2
timestamp 1694700623
transform 1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1694700623
transform -1 0 37856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__A2
timestamp 1694700623
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__B
timestamp 1694700623
transform 1 0 28336 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A2
timestamp 1694700623
transform -1 0 27664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A2
timestamp 1694700623
transform 1 0 51408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1694700623
transform 1 0 50400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__B
timestamp 1694700623
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__I
timestamp 1694700623
transform 1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__I
timestamp 1694700623
transform 1 0 38976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__I
timestamp 1694700623
transform -1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1694700623
transform -1 0 33376 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A1
timestamp 1694700623
transform -1 0 33824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1694700623
transform -1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__C
timestamp 1694700623
transform -1 0 34048 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A1
timestamp 1694700623
transform 1 0 35728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1694700623
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A2
timestamp 1694700623
transform 1 0 35056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__B
timestamp 1694700623
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A1
timestamp 1694700623
transform 1 0 33152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1694700623
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1694700623
transform 1 0 36064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1694700623
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B
timestamp 1694700623
transform -1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1694700623
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1694700623
transform 1 0 28224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1694700623
transform -1 0 26768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__B
timestamp 1694700623
transform 1 0 27440 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__I
timestamp 1694700623
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2210__I
timestamp 1694700623
transform 1 0 24528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__I
timestamp 1694700623
transform 1 0 22176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A2
timestamp 1694700623
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1694700623
transform -1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1694700623
transform -1 0 20272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A1
timestamp 1694700623
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1694700623
transform -1 0 22176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__C
timestamp 1694700623
transform 1 0 22176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A1
timestamp 1694700623
transform 1 0 24304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1694700623
transform -1 0 24304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__A2
timestamp 1694700623
transform -1 0 23408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1694700623
transform 1 0 25200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A1
timestamp 1694700623
transform 1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__A2
timestamp 1694700623
transform 1 0 22400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A1
timestamp 1694700623
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1694700623
transform -1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__B
timestamp 1694700623
transform 1 0 20160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A2
timestamp 1694700623
transform 1 0 19376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__B
timestamp 1694700623
transform 1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A1
timestamp 1694700623
transform -1 0 34160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1694700623
transform -1 0 33712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1694700623
transform -1 0 37968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1694700623
transform 1 0 40992 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__B
timestamp 1694700623
transform 1 0 45920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1694700623
transform 1 0 41664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1694700623
transform 1 0 42224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__A2
timestamp 1694700623
transform 1 0 40992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__B
timestamp 1694700623
transform -1 0 39648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1694700623
transform 1 0 45696 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__B
timestamp 1694700623
transform 1 0 39984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1694700623
transform 1 0 43792 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__B
timestamp 1694700623
transform 1 0 44912 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1694700623
transform 1 0 55216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A1
timestamp 1694700623
transform 1 0 56000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__C
timestamp 1694700623
transform 1 0 57232 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__C
timestamp 1694700623
transform -1 0 53984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1694700623
transform 1 0 51520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1694700623
transform 1 0 51632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1694700623
transform 1 0 52080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1694700623
transform 1 0 47824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1694700623
transform 1 0 47488 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1694700623
transform 1 0 45808 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1694700623
transform 1 0 47936 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1694700623
transform 1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__C2
timestamp 1694700623
transform 1 0 45472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1694700623
transform 1 0 51072 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1694700623
transform -1 0 51296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__I
timestamp 1694700623
transform 1 0 32032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__I
timestamp 1694700623
transform 1 0 22288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__B
timestamp 1694700623
transform -1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1694700623
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__I
timestamp 1694700623
transform 1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1694700623
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1694700623
transform 1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1694700623
transform 1 0 39760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1694700623
transform 1 0 37744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__I
timestamp 1694700623
transform -1 0 33936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A2
timestamp 1694700623
transform -1 0 27776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A1
timestamp 1694700623
transform 1 0 27440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__I
timestamp 1694700623
transform 1 0 35952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1694700623
transform -1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__I
timestamp 1694700623
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1694700623
transform 1 0 30128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__I
timestamp 1694700623
transform -1 0 19824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1694700623
transform 1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A1
timestamp 1694700623
transform 1 0 31360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1694700623
transform 1 0 19264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1694700623
transform -1 0 18368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1694700623
transform 1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1694700623
transform -1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1694700623
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__B
timestamp 1694700623
transform 1 0 22848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1694700623
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1694700623
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1694700623
transform 1 0 32032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__C
timestamp 1694700623
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1694700623
transform 1 0 31808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1694700623
transform 1 0 29232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1694700623
transform -1 0 29456 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A1
timestamp 1694700623
transform 1 0 26880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1694700623
transform -1 0 25536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1694700623
transform -1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1694700623
transform 1 0 21168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1694700623
transform 1 0 20720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1694700623
transform 1 0 29344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1694700623
transform 1 0 15568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__I
timestamp 1694700623
transform -1 0 19600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1694700623
transform 1 0 15120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1694700623
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1694700623
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A1
timestamp 1694700623
transform 1 0 18032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__I
timestamp 1694700623
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1694700623
transform 1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__C
timestamp 1694700623
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2505__A1
timestamp 1694700623
transform -1 0 16016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A1
timestamp 1694700623
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__C
timestamp 1694700623
transform 1 0 18144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1694700623
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__C
timestamp 1694700623
transform -1 0 17920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B
timestamp 1694700623
transform -1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A1
timestamp 1694700623
transform -1 0 22624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__B
timestamp 1694700623
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__C
timestamp 1694700623
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1694700623
transform 1 0 42448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__B
timestamp 1694700623
transform -1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1694700623
transform -1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1694700623
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__A1
timestamp 1694700623
transform 1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__C
timestamp 1694700623
transform 1 0 37744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__CLK
timestamp 1694700623
transform 1 0 42000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__D
timestamp 1694700623
transform 1 0 41552 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2527__CLK
timestamp 1694700623
transform 1 0 30576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__CLK
timestamp 1694700623
transform 1 0 31808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__CLK
timestamp 1694700623
transform 1 0 31584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__CLK
timestamp 1694700623
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__CLK
timestamp 1694700623
transform 1 0 50288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__CLK
timestamp 1694700623
transform 1 0 44352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__CLK
timestamp 1694700623
transform -1 0 44016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__CLK
timestamp 1694700623
transform 1 0 41216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__CLK
timestamp 1694700623
transform 1 0 51184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__CLK
timestamp 1694700623
transform -1 0 50400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__CLK
timestamp 1694700623
transform 1 0 44912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__CLK
timestamp 1694700623
transform -1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__CLK
timestamp 1694700623
transform 1 0 43456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__CLK
timestamp 1694700623
transform 1 0 44240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__CLK
timestamp 1694700623
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__CLK
timestamp 1694700623
transform 1 0 22512 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__CLK
timestamp 1694700623
transform 1 0 19040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__CLK
timestamp 1694700623
transform -1 0 21616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__CLK
timestamp 1694700623
transform 1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__CLK
timestamp 1694700623
transform 1 0 25312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__CLK
timestamp 1694700623
transform 1 0 25872 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__CLK
timestamp 1694700623
transform 1 0 16128 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__CLK
timestamp 1694700623
transform 1 0 23408 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__CLK
timestamp 1694700623
transform -1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__CLK
timestamp 1694700623
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__CLK
timestamp 1694700623
transform 1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__CLK
timestamp 1694700623
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__CLK
timestamp 1694700623
transform 1 0 5376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__CLK
timestamp 1694700623
transform -1 0 5152 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__CLK
timestamp 1694700623
transform 1 0 4816 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__CLK
timestamp 1694700623
transform 1 0 5824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__CLK
timestamp 1694700623
transform 1 0 8736 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__CLK
timestamp 1694700623
transform 1 0 21952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__CLK
timestamp 1694700623
transform 1 0 21392 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__CLK
timestamp 1694700623
transform 1 0 7840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__CLK
timestamp 1694700623
transform 1 0 10192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__CLK
timestamp 1694700623
transform 1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__CLK
timestamp 1694700623
transform 1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__CLK
timestamp 1694700623
transform 1 0 10192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__CLK
timestamp 1694700623
transform -1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__CLK
timestamp 1694700623
transform 1 0 9744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__CLK
timestamp 1694700623
transform 1 0 11312 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1694700623
transform -1 0 12656 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1694700623
transform 1 0 16800 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1694700623
transform -1 0 20944 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__CLK
timestamp 1694700623
transform 1 0 56672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__CLK
timestamp 1694700623
transform 1 0 56224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__CLK
timestamp 1694700623
transform 1 0 54880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__CLK
timestamp 1694700623
transform 1 0 56672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__CLK
timestamp 1694700623
transform 1 0 53312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__CLK
timestamp 1694700623
transform 1 0 52416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__CLK
timestamp 1694700623
transform 1 0 53536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__CLK
timestamp 1694700623
transform 1 0 48720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__CLK
timestamp 1694700623
transform 1 0 50848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1694700623
transform 1 0 54656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1694700623
transform 1 0 53872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1694700623
transform 1 0 54656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1694700623
transform 1 0 55552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1694700623
transform 1 0 58128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1694700623
transform 1 0 58128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__CLK
timestamp 1694700623
transform 1 0 58128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__CLK
timestamp 1694700623
transform 1 0 58128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__CLK
timestamp 1694700623
transform 1 0 58128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__CLK
timestamp 1694700623
transform 1 0 54880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__CLK
timestamp 1694700623
transform 1 0 56672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__CLK
timestamp 1694700623
transform 1 0 56000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__CLK
timestamp 1694700623
transform 1 0 51408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1694700623
transform 1 0 50288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1694700623
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__CLK
timestamp 1694700623
transform 1 0 44352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__CLK
timestamp 1694700623
transform 1 0 45584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__CLK
timestamp 1694700623
transform 1 0 42112 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__CLK
timestamp 1694700623
transform -1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__CLK
timestamp 1694700623
transform 1 0 49952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__CLK
timestamp 1694700623
transform 1 0 49728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__CLK
timestamp 1694700623
transform 1 0 44688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__CLK
timestamp 1694700623
transform 1 0 36624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__CLK
timestamp 1694700623
transform 1 0 34384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__CLK
timestamp 1694700623
transform 1 0 25088 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__CLK
timestamp 1694700623
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__CLK
timestamp 1694700623
transform 1 0 34944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1694700623
transform 1 0 23184 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__CLK
timestamp 1694700623
transform 1 0 27664 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__CLK
timestamp 1694700623
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__CLK
timestamp 1694700623
transform -1 0 25536 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1694700623
transform 1 0 56000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1694700623
transform 1 0 57456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1694700623
transform 1 0 54880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1694700623
transform 1 0 57680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1694700623
transform 1 0 56672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1694700623
transform 1 0 50064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1694700623
transform 1 0 42784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__CLK
timestamp 1694700623
transform 1 0 41440 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__CLK
timestamp 1694700623
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__CLK
timestamp 1694700623
transform 1 0 40992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__CLK
timestamp 1694700623
transform 1 0 28560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1694700623
transform 1 0 55664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__CLK
timestamp 1694700623
transform 1 0 56000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1694700623
transform 1 0 53872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1694700623
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1694700623
transform 1 0 40320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__CLK
timestamp 1694700623
transform 1 0 37632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__CLK
timestamp 1694700623
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__CLK
timestamp 1694700623
transform 1 0 32032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__CLK
timestamp 1694700623
transform 1 0 38304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__CLK
timestamp 1694700623
transform 1 0 38304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1694700623
transform 1 0 9632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1694700623
transform 1 0 29232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1694700623
transform 1 0 28560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__CLK
timestamp 1694700623
transform 1 0 21392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__CLK
timestamp 1694700623
transform -1 0 21728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1694700623
transform 1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1694700623
transform 1 0 17472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1694700623
transform 1 0 17696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__CLK
timestamp 1694700623
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__CLK
timestamp 1694700623
transform 1 0 25312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__CLK
timestamp 1694700623
transform 1 0 23184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1694700623
transform 1 0 14784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__CLK
timestamp 1694700623
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__CLK
timestamp 1694700623
transform 1 0 43792 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__CLK
timestamp 1694700623
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__CLK
timestamp 1694700623
transform 1 0 42112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__CLK
timestamp 1694700623
transform 1 0 42784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1694700623
transform 1 0 40992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1694700623
transform 1 0 48160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1694700623
transform 1 0 41776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1694700623
transform 1 0 45360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1694700623
transform 1 0 44912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1694700623
transform 1 0 54880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1694700623
transform 1 0 54880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1694700623
transform 1 0 54880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__CLK
timestamp 1694700623
transform 1 0 53872 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__CLK
timestamp 1694700623
transform 1 0 54880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__CLK
timestamp 1694700623
transform 1 0 54880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1694700623
transform 1 0 58128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1694700623
transform 1 0 54992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1694700623
transform -1 0 41216 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__D
timestamp 1694700623
transform -1 0 40208 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__CLK
timestamp 1694700623
transform 1 0 54208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__CLK
timestamp 1694700623
transform 1 0 49840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__CLK
timestamp 1694700623
transform 1 0 43232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__CLK
timestamp 1694700623
transform -1 0 51856 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1694700623
transform 1 0 45808 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1694700623
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1694700623
transform 1 0 50400 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1694700623
transform 1 0 50400 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1694700623
transform 1 0 52080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1694700623
transform 1 0 52752 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1694700623
transform -1 0 55552 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1694700623
transform 1 0 54656 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1694700623
transform 1 0 54208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2677__CLK
timestamp 1694700623
transform -1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1694700623
transform -1 0 45584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__CLK
timestamp 1694700623
transform -1 0 41664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1694700623
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1694700623
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1694700623
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1694700623
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1694700623
transform 1 0 29904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1694700623
transform 1 0 30464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1694700623
transform 1 0 30912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1694700623
transform 1 0 28336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1694700623
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1694700623
transform 1 0 33936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1694700623
transform 1 0 19712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1694700623
transform -1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1694700623
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1694700623
transform -1 0 17920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1694700623
transform -1 0 19712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1694700623
transform 1 0 18032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1694700623
transform 1 0 30576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1694700623
transform 1 0 30240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1694700623
transform 1 0 27664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1694700623
transform 1 0 29680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1694700623
transform 1 0 27216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1694700623
transform -1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1694700623
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1694700623
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1694700623
transform 1 0 7168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1694700623
transform 1 0 8064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1694700623
transform 1 0 12768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1694700623
transform 1 0 13328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1694700623
transform 1 0 15008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1694700623
transform 1 0 15904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1694700623
transform 1 0 16352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1694700623
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1694700623
transform 1 0 23968 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1694700623
transform -1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1694700623
transform 1 0 27552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1694700623
transform 1 0 45248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1694700623
transform 1 0 38416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1694700623
transform 1 0 40320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1694700623
transform 1 0 41888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 21168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1694700623
transform -1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 15456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 28896 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 38752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 52864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 39984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 53872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 13328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 14448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1694700623
transform -1 0 25648 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 52752 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 40992 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1694700623
transform 1 0 52528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1694700623
transform -1 0 58352 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1694700623
transform -1 0 57680 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1694700623
transform -1 0 57456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1694700623
transform 1 0 58128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1694700623
transform -1 0 58352 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1694700623
transform -1 0 57680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1694700623
transform -1 0 57904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1694700623
transform -1 0 57680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1694700623
transform -1 0 58352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1694700623
transform -1 0 57456 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1694700623
transform 1 0 1792 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1694700623
transform 1 0 1792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1694700623
transform -1 0 30352 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1694700623
transform 1 0 39424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1694700623
transform 1 0 43008 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 30016 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 17584 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1694700623
transform 1 0 29680 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1694700623
transform 1 0 12544 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1694700623
transform 1 0 25088 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1694700623
transform 1 0 38976 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1694700623
transform 1 0 53088 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1694700623
transform 1 0 40208 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1694700623
transform 1 0 54096 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1694700623
transform -1 0 12544 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1694700623
transform 1 0 18032 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1694700623
transform 1 0 11536 0 -1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1694700623
transform 1 0 21952 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1694700623
transform 1 0 41216 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1694700623
transform 1 0 52976 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1694700623
transform 1 0 41104 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1694700623
transform 1 0 52752 0 1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1694700623
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1694700623
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1694700623
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1694700623
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 20608 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_182 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 21728 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1694700623
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1694700623
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1694700623
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1694700623
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1694700623
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1694700623
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_381
timestamp 1694700623
transform 1 0 44016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_397
timestamp 1694700623
transform 1 0 45808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1694700623
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1694700623
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1694700623
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1694700623
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1694700623
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1694700623
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1694700623
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1694700623
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1694700623
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1694700623
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1694700623
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1694700623
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1694700623
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1694700623
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1694700623
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_241
timestamp 1694700623
transform 1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_245
timestamp 1694700623
transform 1 0 28784 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1694700623
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1694700623
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_286
timestamp 1694700623
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_290
timestamp 1694700623
transform 1 0 33824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_292
timestamp 1694700623
transform 1 0 34048 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_322
timestamp 1694700623
transform 1 0 37408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_326
timestamp 1694700623
transform 1 0 37856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_331
timestamp 1694700623
transform 1 0 38416 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_347
timestamp 1694700623
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1694700623
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_410
timestamp 1694700623
transform 1 0 47264 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1694700623
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_426
timestamp 1694700623
transform 1 0 49056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_434
timestamp 1694700623
transform 1 0 49952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_467
timestamp 1694700623
transform 1 0 53648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_471
timestamp 1694700623
transform 1 0 54096 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_487
timestamp 1694700623
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1694700623
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_492
timestamp 1694700623
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_496
timestamp 1694700623
transform 1 0 56896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_498
timestamp 1694700623
transform 1 0 57120 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1694700623
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1694700623
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1694700623
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1694700623
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1694700623
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_139
timestamp 1694700623
transform 1 0 16912 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_155
timestamp 1694700623
transform 1 0 18704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_163
timestamp 1694700623
transform 1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_165
timestamp 1694700623
transform 1 0 19824 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1694700623
transform 1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1694700623
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1694700623
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_181
timestamp 1694700623
transform 1 0 21616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_189
timestamp 1694700623
transform 1 0 22512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_197
timestamp 1694700623
transform 1 0 23408 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_213
timestamp 1694700623
transform 1 0 25200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_217
timestamp 1694700623
transform 1 0 25648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_223
timestamp 1694700623
transform 1 0 26320 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_239
timestamp 1694700623
transform 1 0 28112 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1694700623
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_247
timestamp 1694700623
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_255
timestamp 1694700623
transform 1 0 29904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_259
timestamp 1694700623
transform 1 0 30352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_268
timestamp 1694700623
transform 1 0 31360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_272
timestamp 1694700623
transform 1 0 31808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_276
timestamp 1694700623
transform 1 0 32256 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_278
timestamp 1694700623
transform 1 0 32480 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_308
timestamp 1694700623
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_312
timestamp 1694700623
transform 1 0 36288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1694700623
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1694700623
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_354
timestamp 1694700623
transform 1 0 40992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_370
timestamp 1694700623
transform 1 0 42784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_378
timestamp 1694700623
transform 1 0 43680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_380
timestamp 1694700623
transform 1 0 43904 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_383
timestamp 1694700623
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1694700623
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_391
timestamp 1694700623
transform 1 0 45136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_393
timestamp 1694700623
transform 1 0 45360 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_404
timestamp 1694700623
transform 1 0 46592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_435
timestamp 1694700623
transform 1 0 50064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_439
timestamp 1694700623
transform 1 0 50512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_443
timestamp 1694700623
transform 1 0 50960 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1694700623
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1694700623
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1694700623
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1694700623
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1694700623
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1694700623
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1694700623
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1694700623
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1694700623
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1694700623
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1694700623
transform 1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1694700623
transform 1 0 18144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_152
timestamp 1694700623
transform 1 0 18368 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_163
timestamp 1694700623
transform 1 0 19600 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_187
timestamp 1694700623
transform 1 0 22288 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1694700623
transform 1 0 23184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_205
timestamp 1694700623
transform 1 0 24304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_209
timestamp 1694700623
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_212
timestamp 1694700623
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_228
timestamp 1694700623
transform 1 0 26880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_232
timestamp 1694700623
transform 1 0 27328 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_262
timestamp 1694700623
transform 1 0 30688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_272
timestamp 1694700623
transform 1 0 31808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_276
timestamp 1694700623
transform 1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_282
timestamp 1694700623
transform 1 0 32928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_286
timestamp 1694700623
transform 1 0 33376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_292
timestamp 1694700623
transform 1 0 34048 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_300
timestamp 1694700623
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_302
timestamp 1694700623
transform 1 0 35168 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_307
timestamp 1694700623
transform 1 0 35728 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_339
timestamp 1694700623
transform 1 0 39312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1694700623
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1694700623
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_352
timestamp 1694700623
transform 1 0 40768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_387
timestamp 1694700623
transform 1 0 44688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_397
timestamp 1694700623
transform 1 0 45808 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_414
timestamp 1694700623
transform 1 0 47712 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_418
timestamp 1694700623
transform 1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1694700623
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1694700623
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1694700623
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1694700623
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1694700623
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1694700623
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1694700623
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1694700623
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1694700623
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_123
timestamp 1694700623
transform 1 0 15120 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_165
timestamp 1694700623
transform 1 0 19824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_189
timestamp 1694700623
transform 1 0 22512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_193
timestamp 1694700623
transform 1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_195
timestamp 1694700623
transform 1 0 23184 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_216
timestamp 1694700623
transform 1 0 25536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_236
timestamp 1694700623
transform 1 0 27776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_240
timestamp 1694700623
transform 1 0 28224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_244
timestamp 1694700623
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1694700623
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_255
timestamp 1694700623
transform 1 0 29904 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_274
timestamp 1694700623
transform 1 0 32032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_278
timestamp 1694700623
transform 1 0 32480 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_312
timestamp 1694700623
transform 1 0 36288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_314
timestamp 1694700623
transform 1 0 36512 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1694700623
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_337
timestamp 1694700623
transform 1 0 39088 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_341
timestamp 1694700623
transform 1 0 39536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_363
timestamp 1694700623
transform 1 0 42000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_367
timestamp 1694700623
transform 1 0 42448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_369
timestamp 1694700623
transform 1 0 42672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_378
timestamp 1694700623
transform 1 0 43680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_382
timestamp 1694700623
transform 1 0 44128 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1694700623
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_387
timestamp 1694700623
transform 1 0 44688 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_395
timestamp 1694700623
transform 1 0 45584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_399
timestamp 1694700623
transform 1 0 46032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_401
timestamp 1694700623
transform 1 0 46256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_404
timestamp 1694700623
transform 1 0 46592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_408
timestamp 1694700623
transform 1 0 47040 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_416
timestamp 1694700623
transform 1 0 47936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_426
timestamp 1694700623
transform 1 0 49056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_448
timestamp 1694700623
transform 1 0 51520 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_452
timestamp 1694700623
transform 1 0 51968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_454
timestamp 1694700623
transform 1 0 52192 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_486
timestamp 1694700623
transform 1 0 55776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_490
timestamp 1694700623
transform 1 0 56224 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_506
timestamp 1694700623
transform 1 0 58016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_508
timestamp 1694700623
transform 1 0 58240 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1694700623
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1694700623
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1694700623
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1694700623
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1694700623
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_150
timestamp 1694700623
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_170
timestamp 1694700623
transform 1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_180
timestamp 1694700623
transform 1 0 21504 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_188
timestamp 1694700623
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1694700623
transform 1 0 25088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_216
timestamp 1694700623
transform 1 0 25536 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_233
timestamp 1694700623
transform 1 0 27440 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_263
timestamp 1694700623
transform 1 0 30800 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_267
timestamp 1694700623
transform 1 0 31248 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_270
timestamp 1694700623
transform 1 0 31584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_274
timestamp 1694700623
transform 1 0 32032 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_278
timestamp 1694700623
transform 1 0 32480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_282
timestamp 1694700623
transform 1 0 32928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_286
timestamp 1694700623
transform 1 0 33376 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_299
timestamp 1694700623
transform 1 0 34832 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_318
timestamp 1694700623
transform 1 0 36960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_338
timestamp 1694700623
transform 1 0 39200 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_360
timestamp 1694700623
transform 1 0 41664 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_384
timestamp 1694700623
transform 1 0 44352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_388
timestamp 1694700623
transform 1 0 44800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_396
timestamp 1694700623
transform 1 0 45696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_399
timestamp 1694700623
transform 1 0 46032 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_415
timestamp 1694700623
transform 1 0 47824 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_419
timestamp 1694700623
transform 1 0 48272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_422
timestamp 1694700623
transform 1 0 48608 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_450
timestamp 1694700623
transform 1 0 51744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_454
timestamp 1694700623
transform 1 0 52192 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_459
timestamp 1694700623
transform 1 0 52752 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_475
timestamp 1694700623
transform 1 0 54544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_483
timestamp 1694700623
transform 1 0 55440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_487
timestamp 1694700623
transform 1 0 55888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_489
timestamp 1694700623
transform 1 0 56112 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1694700623
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1694700623
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1694700623
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1694700623
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1694700623
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1694700623
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1694700623
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1694700623
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_177
timestamp 1694700623
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_209
timestamp 1694700623
transform 1 0 24752 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_233
timestamp 1694700623
transform 1 0 27440 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1694700623
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1694700623
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1694700623
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_259
timestamp 1694700623
transform 1 0 30352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_276
timestamp 1694700623
transform 1 0 32256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_280
timestamp 1694700623
transform 1 0 32704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_284
timestamp 1694700623
transform 1 0 33152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_286
timestamp 1694700623
transform 1 0 33376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_293
timestamp 1694700623
transform 1 0 34160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_297
timestamp 1694700623
transform 1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1694700623
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_333
timestamp 1694700623
transform 1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_335
timestamp 1694700623
transform 1 0 38864 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_344
timestamp 1694700623
transform 1 0 39872 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_376
timestamp 1694700623
transform 1 0 43456 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_384
timestamp 1694700623
transform 1 0 44352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_387
timestamp 1694700623
transform 1 0 44688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_407
timestamp 1694700623
transform 1 0 46928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_409
timestamp 1694700623
transform 1 0 47152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1694700623
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1694700623
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1694700623
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1694700623
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1694700623
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1694700623
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_72
timestamp 1694700623
transform 1 0 9408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_104
timestamp 1694700623
transform 1 0 12992 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_108
timestamp 1694700623
transform 1 0 13440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_110
timestamp 1694700623
transform 1 0 13664 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1694700623
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_146
timestamp 1694700623
transform 1 0 17696 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_162
timestamp 1694700623
transform 1 0 19488 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_178
timestamp 1694700623
transform 1 0 21280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_182
timestamp 1694700623
transform 1 0 21728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_190
timestamp 1694700623
transform 1 0 22624 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1694700623
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_212
timestamp 1694700623
transform 1 0 25088 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_244
timestamp 1694700623
transform 1 0 28672 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_260
timestamp 1694700623
transform 1 0 30464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1694700623
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1694700623
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1694700623
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_291
timestamp 1694700623
transform 1 0 33936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_307
timestamp 1694700623
transform 1 0 35728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_315
timestamp 1694700623
transform 1 0 36624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_317
timestamp 1694700623
transform 1 0 36848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_326
timestamp 1694700623
transform 1 0 37856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_334
timestamp 1694700623
transform 1 0 38752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_336
timestamp 1694700623
transform 1 0 38976 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1694700623
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_352
timestamp 1694700623
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_360
timestamp 1694700623
transform 1 0 41664 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_381
timestamp 1694700623
transform 1 0 44016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_383
timestamp 1694700623
transform 1 0 44240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_415
timestamp 1694700623
transform 1 0 47824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1694700623
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_422
timestamp 1694700623
transform 1 0 48608 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_430
timestamp 1694700623
transform 1 0 49504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_440
timestamp 1694700623
transform 1 0 50624 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_448
timestamp 1694700623
transform 1 0 51520 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_452
timestamp 1694700623
transform 1 0 51968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_483
timestamp 1694700623
transform 1 0 55440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_487
timestamp 1694700623
transform 1 0 55888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_489
timestamp 1694700623
transform 1 0 56112 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1694700623
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1694700623
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1694700623
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1694700623
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1694700623
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1694700623
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_107
timestamp 1694700623
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_123
timestamp 1694700623
transform 1 0 15120 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_127
timestamp 1694700623
transform 1 0 15568 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_132
timestamp 1694700623
transform 1 0 16128 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_140
timestamp 1694700623
transform 1 0 17024 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_164
timestamp 1694700623
transform 1 0 19712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_168
timestamp 1694700623
transform 1 0 20160 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1694700623
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1694700623
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_177
timestamp 1694700623
transform 1 0 21168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_184
timestamp 1694700623
transform 1 0 21952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_188
timestamp 1694700623
transform 1 0 22400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_192
timestamp 1694700623
transform 1 0 22848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_194
timestamp 1694700623
transform 1 0 23072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1694700623
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_251
timestamp 1694700623
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_253
timestamp 1694700623
transform 1 0 29680 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_274
timestamp 1694700623
transform 1 0 32032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_278
timestamp 1694700623
transform 1 0 32480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_298
timestamp 1694700623
transform 1 0 34720 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_302
timestamp 1694700623
transform 1 0 35168 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1694700623
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_321
timestamp 1694700623
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_360
timestamp 1694700623
transform 1 0 41664 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_384
timestamp 1694700623
transform 1 0 44352 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_387
timestamp 1694700623
transform 1 0 44688 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_419
timestamp 1694700623
transform 1 0 48272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_435
timestamp 1694700623
transform 1 0 50064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_437
timestamp 1694700623
transform 1 0 50288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_445
timestamp 1694700623
transform 1 0 51184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_449
timestamp 1694700623
transform 1 0 51632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_465
timestamp 1694700623
transform 1 0 53424 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_497
timestamp 1694700623
transform 1 0 57008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1694700623
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1694700623
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1694700623
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_72
timestamp 1694700623
transform 1 0 9408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_104
timestamp 1694700623
transform 1 0 12992 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_120
timestamp 1694700623
transform 1 0 14784 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_132
timestamp 1694700623
transform 1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1694700623
transform 1 0 17248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_166
timestamp 1694700623
transform 1 0 19936 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_174
timestamp 1694700623
transform 1 0 20832 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_178
timestamp 1694700623
transform 1 0 21280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1694700623
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_212
timestamp 1694700623
transform 1 0 25088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_216
timestamp 1694700623
transform 1 0 25536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_224
timestamp 1694700623
transform 1 0 26432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_261
timestamp 1694700623
transform 1 0 30576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_263
timestamp 1694700623
transform 1 0 30800 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_269
timestamp 1694700623
transform 1 0 31472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_273
timestamp 1694700623
transform 1 0 31920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1694700623
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1694700623
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1694700623
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1694700623
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_352
timestamp 1694700623
transform 1 0 40768 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_356
timestamp 1694700623
transform 1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_358
timestamp 1694700623
transform 1 0 41440 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_367
timestamp 1694700623
transform 1 0 42448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_369
timestamp 1694700623
transform 1 0 42672 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_401
timestamp 1694700623
transform 1 0 46256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_411
timestamp 1694700623
transform 1 0 47376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1694700623
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_422
timestamp 1694700623
transform 1 0 48608 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_438
timestamp 1694700623
transform 1 0 50400 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_442
timestamp 1694700623
transform 1 0 50848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_444
timestamp 1694700623
transform 1 0 51072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_450
timestamp 1694700623
transform 1 0 51744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_454
timestamp 1694700623
transform 1 0 52192 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1694700623
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_492
timestamp 1694700623
transform 1 0 56448 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_500
timestamp 1694700623
transform 1 0 57344 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_504
timestamp 1694700623
transform 1 0 57792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_506
timestamp 1694700623
transform 1 0 58016 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1694700623
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1694700623
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1694700623
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1694700623
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1694700623
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_144
timestamp 1694700623
transform 1 0 17472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_148
timestamp 1694700623
transform 1 0 17920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_152
timestamp 1694700623
transform 1 0 18368 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_165
timestamp 1694700623
transform 1 0 19824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1694700623
transform 1 0 20272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_173
timestamp 1694700623
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_183
timestamp 1694700623
transform 1 0 21840 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_199
timestamp 1694700623
transform 1 0 23632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1694700623
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1694700623
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1694700623
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_251
timestamp 1694700623
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_255
timestamp 1694700623
transform 1 0 29904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_259
timestamp 1694700623
transform 1 0 30352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_263
timestamp 1694700623
transform 1 0 30800 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_267
timestamp 1694700623
transform 1 0 31248 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_280
timestamp 1694700623
transform 1 0 32704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_284
timestamp 1694700623
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_288
timestamp 1694700623
transform 1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_292
timestamp 1694700623
transform 1 0 34048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_300
timestamp 1694700623
transform 1 0 34944 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_303
timestamp 1694700623
transform 1 0 35280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1694700623
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1694700623
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1694700623
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_328
timestamp 1694700623
transform 1 0 38080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_338
timestamp 1694700623
transform 1 0 39200 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_370
timestamp 1694700623
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_374
timestamp 1694700623
transform 1 0 43232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1694700623
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1694700623
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_387
timestamp 1694700623
transform 1 0 44688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_403
timestamp 1694700623
transform 1 0 46480 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_433
timestamp 1694700623
transform 1 0 49840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_437
timestamp 1694700623
transform 1 0 50288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_441
timestamp 1694700623
transform 1 0 50736 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_486
timestamp 1694700623
transform 1 0 55776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_490
timestamp 1694700623
transform 1 0 56224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_502
timestamp 1694700623
transform 1 0 57568 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1694700623
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1694700623
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1694700623
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1694700623
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1694700623
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1694700623
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_171
timestamp 1694700623
transform 1 0 20496 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_175
timestamp 1694700623
transform 1 0 20944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_179
timestamp 1694700623
transform 1 0 21392 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_197
timestamp 1694700623
transform 1 0 23408 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_201
timestamp 1694700623
transform 1 0 23856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_205
timestamp 1694700623
transform 1 0 24304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1694700623
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1694700623
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1694700623
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_224
timestamp 1694700623
transform 1 0 26432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1694700623
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_242
timestamp 1694700623
transform 1 0 28448 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_250
timestamp 1694700623
transform 1 0 29344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_252
timestamp 1694700623
transform 1 0 29568 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1694700623
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_290
timestamp 1694700623
transform 1 0 33824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_292
timestamp 1694700623
transform 1 0 34048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_330
timestamp 1694700623
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_332
timestamp 1694700623
transform 1 0 38528 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1694700623
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_358
timestamp 1694700623
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_362
timestamp 1694700623
transform 1 0 41888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_366
timestamp 1694700623
transform 1 0 42336 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_370
timestamp 1694700623
transform 1 0 42784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_378
timestamp 1694700623
transform 1 0 43680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_382
timestamp 1694700623
transform 1 0 44128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_384
timestamp 1694700623
transform 1 0 44352 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_389
timestamp 1694700623
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_405
timestamp 1694700623
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_417
timestamp 1694700623
transform 1 0 48048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1694700623
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_422
timestamp 1694700623
transform 1 0 48608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_430
timestamp 1694700623
transform 1 0 49504 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_456
timestamp 1694700623
transform 1 0 52416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_460
timestamp 1694700623
transform 1 0 52864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_488
timestamp 1694700623
transform 1 0 56000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1694700623
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1694700623
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1694700623
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1694700623
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1694700623
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1694700623
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1694700623
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_139
timestamp 1694700623
transform 1 0 16912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_143
timestamp 1694700623
transform 1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1694700623
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_183
timestamp 1694700623
transform 1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_211
timestamp 1694700623
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215
timestamp 1694700623
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_231
timestamp 1694700623
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_235
timestamp 1694700623
transform 1 0 27664 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1694700623
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1694700623
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_249
timestamp 1694700623
transform 1 0 29232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_293
timestamp 1694700623
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_311
timestamp 1694700623
transform 1 0 36176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1694700623
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_321
timestamp 1694700623
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_329
timestamp 1694700623
transform 1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_333
timestamp 1694700623
transform 1 0 38640 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_368
timestamp 1694700623
transform 1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_372
timestamp 1694700623
transform 1 0 43008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_374
timestamp 1694700623
transform 1 0 43232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1694700623
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_399
timestamp 1694700623
transform 1 0 46032 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_407
timestamp 1694700623
transform 1 0 46928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_420
timestamp 1694700623
transform 1 0 48384 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_436
timestamp 1694700623
transform 1 0 50176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_440
timestamp 1694700623
transform 1 0 50624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_442
timestamp 1694700623
transform 1 0 50848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_445
timestamp 1694700623
transform 1 0 51184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_449
timestamp 1694700623
transform 1 0 51632 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_453
timestamp 1694700623
transform 1 0 52080 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_457
timestamp 1694700623
transform 1 0 52528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_459
timestamp 1694700623
transform 1 0 52752 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_462
timestamp 1694700623
transform 1 0 53088 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_494
timestamp 1694700623
transform 1 0 56672 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_502
timestamp 1694700623
transform 1 0 57568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_506
timestamp 1694700623
transform 1 0 58016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_508
timestamp 1694700623
transform 1 0 58240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1694700623
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1694700623
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1694700623
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1694700623
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1694700623
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1694700623
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1694700623
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_146
timestamp 1694700623
transform 1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_150
timestamp 1694700623
transform 1 0 18144 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1694700623
transform 1 0 21952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_203
timestamp 1694700623
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1694700623
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1694700623
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_212
timestamp 1694700623
transform 1 0 25088 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_228
timestamp 1694700623
transform 1 0 26880 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_258
timestamp 1694700623
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_262
timestamp 1694700623
transform 1 0 30688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_270
timestamp 1694700623
transform 1 0 31584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_288
timestamp 1694700623
transform 1 0 33600 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_305
timestamp 1694700623
transform 1 0 35504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_309
timestamp 1694700623
transform 1 0 35952 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_317
timestamp 1694700623
transform 1 0 36848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_321
timestamp 1694700623
transform 1 0 37296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_325
timestamp 1694700623
transform 1 0 37744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_329
timestamp 1694700623
transform 1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_333
timestamp 1694700623
transform 1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_343
timestamp 1694700623
transform 1 0 39760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1694700623
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1694700623
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_352
timestamp 1694700623
transform 1 0 40768 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_356
timestamp 1694700623
transform 1 0 41216 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_372
timestamp 1694700623
transform 1 0 43008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_376
timestamp 1694700623
transform 1 0 43456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_385
timestamp 1694700623
transform 1 0 44464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_393
timestamp 1694700623
transform 1 0 45360 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_417
timestamp 1694700623
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1694700623
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_422
timestamp 1694700623
transform 1 0 48608 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_430
timestamp 1694700623
transform 1 0 49504 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_434
timestamp 1694700623
transform 1 0 49952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_444
timestamp 1694700623
transform 1 0 51072 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_452
timestamp 1694700623
transform 1 0 51968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_456
timestamp 1694700623
transform 1 0 52416 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_492
timestamp 1694700623
transform 1 0 56448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_496
timestamp 1694700623
transform 1 0 56896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_504
timestamp 1694700623
transform 1 0 57792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1694700623
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1694700623
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1694700623
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1694700623
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1694700623
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1694700623
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1694700623
transform 1 0 16912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_147
timestamp 1694700623
transform 1 0 17808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_149
timestamp 1694700623
transform 1 0 18032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_158
timestamp 1694700623
transform 1 0 19040 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1694700623
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1694700623
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1694700623
transform 1 0 21616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_183
timestamp 1694700623
transform 1 0 21840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_186
timestamp 1694700623
transform 1 0 22176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_192
timestamp 1694700623
transform 1 0 22848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_194
timestamp 1694700623
transform 1 0 23072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_232
timestamp 1694700623
transform 1 0 27328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_236
timestamp 1694700623
transform 1 0 27776 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1694700623
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_247
timestamp 1694700623
transform 1 0 29008 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_279
timestamp 1694700623
transform 1 0 32592 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_287
timestamp 1694700623
transform 1 0 33488 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_290
timestamp 1694700623
transform 1 0 33824 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_306
timestamp 1694700623
transform 1 0 35616 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1694700623
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1694700623
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_346
timestamp 1694700623
transform 1 0 40096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_350
timestamp 1694700623
transform 1 0 40544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_352
timestamp 1694700623
transform 1 0 40768 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_375
timestamp 1694700623
transform 1 0 43344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_377
timestamp 1694700623
transform 1 0 43568 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_380
timestamp 1694700623
transform 1 0 43904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1694700623
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_392
timestamp 1694700623
transform 1 0 45248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_400
timestamp 1694700623
transform 1 0 46144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_402
timestamp 1694700623
transform 1 0 46368 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_419
timestamp 1694700623
transform 1 0 48272 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_469
timestamp 1694700623
transform 1 0 53872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_471
timestamp 1694700623
transform 1 0 54096 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_501
timestamp 1694700623
transform 1 0 57456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1694700623
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1694700623
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1694700623
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1694700623
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1694700623
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_142
timestamp 1694700623
transform 1 0 17248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_174
timestamp 1694700623
transform 1 0 20832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_190
timestamp 1694700623
transform 1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_192
timestamp 1694700623
transform 1 0 22848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1694700623
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1694700623
transform 1 0 25088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1694700623
transform 1 0 25984 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_253
timestamp 1694700623
transform 1 0 29680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_257
timestamp 1694700623
transform 1 0 30128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_265
timestamp 1694700623
transform 1 0 31024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_267
timestamp 1694700623
transform 1 0 31248 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1694700623
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_282
timestamp 1694700623
transform 1 0 32928 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1694700623
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_397
timestamp 1694700623
transform 1 0 45808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_401
timestamp 1694700623
transform 1 0 46256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_415
timestamp 1694700623
transform 1 0 47824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1694700623
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_422
timestamp 1694700623
transform 1 0 48608 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_431
timestamp 1694700623
transform 1 0 49616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_433
timestamp 1694700623
transform 1 0 49840 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_442
timestamp 1694700623
transform 1 0 50848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_459
timestamp 1694700623
transform 1 0 52752 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_467
timestamp 1694700623
transform 1 0 53648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_469
timestamp 1694700623
transform 1 0 53872 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_474
timestamp 1694700623
transform 1 0 54432 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1694700623
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1694700623
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1694700623
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1694700623
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1694700623
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1694700623
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1694700623
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_123
timestamp 1694700623
transform 1 0 15120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_127
timestamp 1694700623
transform 1 0 15568 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_157
timestamp 1694700623
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_159
timestamp 1694700623
transform 1 0 19152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_162
timestamp 1694700623
transform 1 0 19488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_166
timestamp 1694700623
transform 1 0 19936 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1694700623
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1694700623
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_185
timestamp 1694700623
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1694700623
transform 1 0 22288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_198
timestamp 1694700623
transform 1 0 23520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_202
timestamp 1694700623
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_204
timestamp 1694700623
transform 1 0 24192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_211
timestamp 1694700623
transform 1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_215
timestamp 1694700623
transform 1 0 25424 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_231
timestamp 1694700623
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1694700623
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_247
timestamp 1694700623
transform 1 0 29008 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_256
timestamp 1694700623
transform 1 0 30016 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_272
timestamp 1694700623
transform 1 0 31808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_282
timestamp 1694700623
transform 1 0 32928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_286
timestamp 1694700623
transform 1 0 33376 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_296
timestamp 1694700623
transform 1 0 34496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_300
timestamp 1694700623
transform 1 0 34944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_308
timestamp 1694700623
transform 1 0 35840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1694700623
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1694700623
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1694700623
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_325
timestamp 1694700623
transform 1 0 37744 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_328
timestamp 1694700623
transform 1 0 38080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_332
timestamp 1694700623
transform 1 0 38528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_348
timestamp 1694700623
transform 1 0 40320 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_356
timestamp 1694700623
transform 1 0 41216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_360
timestamp 1694700623
transform 1 0 41664 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_376
timestamp 1694700623
transform 1 0 43456 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_384
timestamp 1694700623
transform 1 0 44352 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_387
timestamp 1694700623
transform 1 0 44688 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_391
timestamp 1694700623
transform 1 0 45136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_398
timestamp 1694700623
transform 1 0 45920 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_451
timestamp 1694700623
transform 1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_457
timestamp 1694700623
transform 1 0 52528 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_473
timestamp 1694700623
transform 1 0 54320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_477
timestamp 1694700623
transform 1 0 54768 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1694700623
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1694700623
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1694700623
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1694700623
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_108
timestamp 1694700623
transform 1 0 13440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1694700623
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1694700623
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1694700623
transform 1 0 17696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_160
timestamp 1694700623
transform 1 0 19264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1694700623
transform 1 0 22960 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1694700623
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1694700623
transform 1 0 25088 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_228
timestamp 1694700623
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_232
timestamp 1694700623
transform 1 0 27328 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1694700623
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_286
timestamp 1694700623
transform 1 0 33376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_290
timestamp 1694700623
transform 1 0 33824 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_322
timestamp 1694700623
transform 1 0 37408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_338
timestamp 1694700623
transform 1 0 39200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1694700623
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1694700623
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_356
timestamp 1694700623
transform 1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_360
timestamp 1694700623
transform 1 0 41664 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_392
timestamp 1694700623
transform 1 0 45248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_408
timestamp 1694700623
transform 1 0 47040 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1694700623
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_422
timestamp 1694700623
transform 1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_430
timestamp 1694700623
transform 1 0 49504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_438
timestamp 1694700623
transform 1 0 50400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_442
timestamp 1694700623
transform 1 0 50848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_444
timestamp 1694700623
transform 1 0 51072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_455
timestamp 1694700623
transform 1 0 52304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_459
timestamp 1694700623
transform 1 0 52752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_472
timestamp 1694700623
transform 1 0 54208 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_488
timestamp 1694700623
transform 1 0 56000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_492
timestamp 1694700623
transform 1 0 56448 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_500
timestamp 1694700623
transform 1 0 57344 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_503
timestamp 1694700623
transform 1 0 57680 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1694700623
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1694700623
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1694700623
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1694700623
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1694700623
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_139
timestamp 1694700623
transform 1 0 16912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1694700623
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1694700623
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1694700623
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_185
timestamp 1694700623
transform 1 0 22064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_189
timestamp 1694700623
transform 1 0 22512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_196
timestamp 1694700623
transform 1 0 23296 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_228
timestamp 1694700623
transform 1 0 26880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1694700623
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_240
timestamp 1694700623
transform 1 0 28224 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1694700623
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_247
timestamp 1694700623
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_255
timestamp 1694700623
transform 1 0 29904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_259
timestamp 1694700623
transform 1 0 30352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_276
timestamp 1694700623
transform 1 0 32256 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_292
timestamp 1694700623
transform 1 0 34048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_296
timestamp 1694700623
transform 1 0 34496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_298
timestamp 1694700623
transform 1 0 34720 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_307
timestamp 1694700623
transform 1 0 35728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1694700623
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1694700623
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1694700623
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_323
timestamp 1694700623
transform 1 0 37520 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_353
timestamp 1694700623
transform 1 0 40880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_355
timestamp 1694700623
transform 1 0 41104 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1694700623
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_391
timestamp 1694700623
transform 1 0 45136 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_399
timestamp 1694700623
transform 1 0 46032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_403
timestamp 1694700623
transform 1 0 46480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_414
timestamp 1694700623
transform 1 0 47712 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_430
timestamp 1694700623
transform 1 0 49504 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_434
timestamp 1694700623
transform 1 0 49952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_436
timestamp 1694700623
transform 1 0 50176 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_453
timestamp 1694700623
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_469
timestamp 1694700623
transform 1 0 53872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_471
timestamp 1694700623
transform 1 0 54096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_501
timestamp 1694700623
transform 1 0 57456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1694700623
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1694700623
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1694700623
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1694700623
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1694700623
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1694700623
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_155
timestamp 1694700623
transform 1 0 18704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_159
timestamp 1694700623
transform 1 0 19152 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_175
timestamp 1694700623
transform 1 0 20944 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_179
timestamp 1694700623
transform 1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_189
timestamp 1694700623
transform 1 0 22512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_191
timestamp 1694700623
transform 1 0 22736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1694700623
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_249
timestamp 1694700623
transform 1 0 29232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_265
timestamp 1694700623
transform 1 0 31024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_267
timestamp 1694700623
transform 1 0 31248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_270
timestamp 1694700623
transform 1 0 31584 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1694700623
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1694700623
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_300
timestamp 1694700623
transform 1 0 34944 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_330
timestamp 1694700623
transform 1 0 38304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_334
timestamp 1694700623
transform 1 0 38752 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_338
timestamp 1694700623
transform 1 0 39200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_348
timestamp 1694700623
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1694700623
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1694700623
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_371
timestamp 1694700623
transform 1 0 42896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_375
timestamp 1694700623
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_387
timestamp 1694700623
transform 1 0 44688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1694700623
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_422
timestamp 1694700623
transform 1 0 48608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_430
timestamp 1694700623
transform 1 0 49504 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_434
timestamp 1694700623
transform 1 0 49952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_436
timestamp 1694700623
transform 1 0 50176 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_450
timestamp 1694700623
transform 1 0 51744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_452
timestamp 1694700623
transform 1 0 51968 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_477
timestamp 1694700623
transform 1 0 54768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1694700623
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1694700623
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1694700623
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1694700623
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1694700623
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1694700623
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1694700623
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1694700623
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1694700623
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1694700623
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_144
timestamp 1694700623
transform 1 0 17472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_148
timestamp 1694700623
transform 1 0 17920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_158
timestamp 1694700623
transform 1 0 19040 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1694700623
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1694700623
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_193
timestamp 1694700623
transform 1 0 22960 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_197
timestamp 1694700623
transform 1 0 23408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_207
timestamp 1694700623
transform 1 0 24528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_215
timestamp 1694700623
transform 1 0 25424 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_219
timestamp 1694700623
transform 1 0 25872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_221
timestamp 1694700623
transform 1 0 26096 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_232
timestamp 1694700623
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_240
timestamp 1694700623
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1694700623
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_247
timestamp 1694700623
transform 1 0 29008 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_251
timestamp 1694700623
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_253
timestamp 1694700623
transform 1 0 29680 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_262
timestamp 1694700623
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_266
timestamp 1694700623
transform 1 0 31136 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_282
timestamp 1694700623
transform 1 0 32928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_286
timestamp 1694700623
transform 1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_302
timestamp 1694700623
transform 1 0 35168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_306
timestamp 1694700623
transform 1 0 35616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_310
timestamp 1694700623
transform 1 0 36064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1694700623
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_341
timestamp 1694700623
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_345
timestamp 1694700623
transform 1 0 39984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_353
timestamp 1694700623
transform 1 0 40880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_357
timestamp 1694700623
transform 1 0 41328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_367
timestamp 1694700623
transform 1 0 42448 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1694700623
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_387
timestamp 1694700623
transform 1 0 44688 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_391
timestamp 1694700623
transform 1 0 45136 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_402
timestamp 1694700623
transform 1 0 46368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_406
timestamp 1694700623
transform 1 0 46816 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_436
timestamp 1694700623
transform 1 0 50176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1694700623
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_457
timestamp 1694700623
transform 1 0 52528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_461
timestamp 1694700623
transform 1 0 52976 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_493
timestamp 1694700623
transform 1 0 56560 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1694700623
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1694700623
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1694700623
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1694700623
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1694700623
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1694700623
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1694700623
transform 1 0 17920 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_159
timestamp 1694700623
transform 1 0 19152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_189
timestamp 1694700623
transform 1 0 22512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1694700623
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1694700623
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1694700623
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_220
timestamp 1694700623
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_222
timestamp 1694700623
transform 1 0 26208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1694700623
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1694700623
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_322
timestamp 1694700623
transform 1 0 37408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_324
timestamp 1694700623
transform 1 0 37632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_327
timestamp 1694700623
transform 1 0 37968 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_343
timestamp 1694700623
transform 1 0 39760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_347
timestamp 1694700623
transform 1 0 40208 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_389
timestamp 1694700623
transform 1 0 44912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_397
timestamp 1694700623
transform 1 0 45808 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1694700623
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_422
timestamp 1694700623
transform 1 0 48608 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_430
timestamp 1694700623
transform 1 0 49504 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_434
timestamp 1694700623
transform 1 0 49952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_438
timestamp 1694700623
transform 1 0 50400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_442
timestamp 1694700623
transform 1 0 50848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_446
timestamp 1694700623
transform 1 0 51296 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_478
timestamp 1694700623
transform 1 0 54880 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1694700623
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_492
timestamp 1694700623
transform 1 0 56448 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_500
timestamp 1694700623
transform 1 0 57344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_504
timestamp 1694700623
transform 1 0 57792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_506
timestamp 1694700623
transform 1 0 58016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1694700623
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1694700623
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1694700623
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1694700623
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1694700623
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1694700623
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_158
timestamp 1694700623
transform 1 0 19040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_162
timestamp 1694700623
transform 1 0 19488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_166
timestamp 1694700623
transform 1 0 19936 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1694700623
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1694700623
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_190
timestamp 1694700623
transform 1 0 22624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_194
timestamp 1694700623
transform 1 0 23072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_202
timestamp 1694700623
transform 1 0 23968 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_206
timestamp 1694700623
transform 1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_208
timestamp 1694700623
transform 1 0 24640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_211
timestamp 1694700623
transform 1 0 24976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_227
timestamp 1694700623
transform 1 0 26768 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_235
timestamp 1694700623
transform 1 0 27664 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1694700623
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1694700623
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_255
timestamp 1694700623
transform 1 0 29904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_259
timestamp 1694700623
transform 1 0 30352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_289
timestamp 1694700623
transform 1 0 33712 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_293
timestamp 1694700623
transform 1 0 34160 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1694700623
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1694700623
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1694700623
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_349
timestamp 1694700623
transform 1 0 40432 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_357
timestamp 1694700623
transform 1 0 41328 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_360
timestamp 1694700623
transform 1 0 41664 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_376
timestamp 1694700623
transform 1 0 43456 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1694700623
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_387
timestamp 1694700623
transform 1 0 44688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_403
timestamp 1694700623
transform 1 0 46480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_407
timestamp 1694700623
transform 1 0 46928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_411
timestamp 1694700623
transform 1 0 47376 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_443
timestamp 1694700623
transform 1 0 50960 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1694700623
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_457
timestamp 1694700623
transform 1 0 52528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_473
timestamp 1694700623
transform 1 0 54320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_477
timestamp 1694700623
transform 1 0 54768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_479
timestamp 1694700623
transform 1 0 54992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1694700623
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1694700623
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1694700623
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1694700623
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1694700623
transform 1 0 17248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_168
timestamp 1694700623
transform 1 0 20160 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_176
timestamp 1694700623
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1694700623
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_249
timestamp 1694700623
transform 1 0 29232 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_265
timestamp 1694700623
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1694700623
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1694700623
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1694700623
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_282
timestamp 1694700623
transform 1 0 32928 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_286
timestamp 1694700623
transform 1 0 33376 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_321
timestamp 1694700623
transform 1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_323
timestamp 1694700623
transform 1 0 37520 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_326
timestamp 1694700623
transform 1 0 37856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_340
timestamp 1694700623
transform 1 0 39424 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1694700623
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_354
timestamp 1694700623
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_363
timestamp 1694700623
transform 1 0 42000 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_379
timestamp 1694700623
transform 1 0 43792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_387
timestamp 1694700623
transform 1 0 44688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_391
timestamp 1694700623
transform 1 0 45136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_395
timestamp 1694700623
transform 1 0 45584 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_399
timestamp 1694700623
transform 1 0 46032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_401
timestamp 1694700623
transform 1 0 46256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_404
timestamp 1694700623
transform 1 0 46592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_413
timestamp 1694700623
transform 1 0 47600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1694700623
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1694700623
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_422
timestamp 1694700623
transform 1 0 48608 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_434
timestamp 1694700623
transform 1 0 49952 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_450
timestamp 1694700623
transform 1 0 51744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_452
timestamp 1694700623
transform 1 0 51968 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_482
timestamp 1694700623
transform 1 0 55328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1694700623
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_500
timestamp 1694700623
transform 1 0 57344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1694700623
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1694700623
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1694700623
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1694700623
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1694700623
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1694700623
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1694700623
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_177
timestamp 1694700623
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_193
timestamp 1694700623
transform 1 0 22960 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_197
timestamp 1694700623
transform 1 0 23408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_199
timestamp 1694700623
transform 1 0 23632 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_247
timestamp 1694700623
transform 1 0 29008 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_279
timestamp 1694700623
transform 1 0 32592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_283
timestamp 1694700623
transform 1 0 33040 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_317
timestamp 1694700623
transform 1 0 36848 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_353
timestamp 1694700623
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1694700623
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1694700623
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_391
timestamp 1694700623
transform 1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_403
timestamp 1694700623
transform 1 0 46480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_443
timestamp 1694700623
transform 1 0 50960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_447
timestamp 1694700623
transform 1 0 51408 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_457
timestamp 1694700623
transform 1 0 52528 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_473
timestamp 1694700623
transform 1 0 54320 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_482
timestamp 1694700623
transform 1 0 55328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_490
timestamp 1694700623
transform 1 0 56224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_507
timestamp 1694700623
transform 1 0 58128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1694700623
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1694700623
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1694700623
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_104
timestamp 1694700623
transform 1 0 12992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_108
timestamp 1694700623
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_110
timestamp 1694700623
transform 1 0 13664 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1694700623
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_146
timestamp 1694700623
transform 1 0 17696 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_162
timestamp 1694700623
transform 1 0 19488 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_165
timestamp 1694700623
transform 1 0 19824 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_181
timestamp 1694700623
transform 1 0 21616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_185
timestamp 1694700623
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_195
timestamp 1694700623
transform 1 0 23184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1694700623
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1694700623
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_221
timestamp 1694700623
transform 1 0 26096 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_229
timestamp 1694700623
transform 1 0 26992 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_233
timestamp 1694700623
transform 1 0 27440 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1694700623
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1694700623
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1694700623
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1694700623
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_290
timestamp 1694700623
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_294
timestamp 1694700623
transform 1 0 34272 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_326
timestamp 1694700623
transform 1 0 37856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_336
timestamp 1694700623
transform 1 0 38976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_340
timestamp 1694700623
transform 1 0 39424 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1694700623
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_352
timestamp 1694700623
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_356
timestamp 1694700623
transform 1 0 41216 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_370
timestamp 1694700623
transform 1 0 42784 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_384
timestamp 1694700623
transform 1 0 44352 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_422
timestamp 1694700623
transform 1 0 48608 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_438
timestamp 1694700623
transform 1 0 50400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_468
timestamp 1694700623
transform 1 0 53760 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_474
timestamp 1694700623
transform 1 0 54432 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_478
timestamp 1694700623
transform 1 0 54880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1694700623
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_497
timestamp 1694700623
transform 1 0 57008 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_505
timestamp 1694700623
transform 1 0 57904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1694700623
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1694700623
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1694700623
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1694700623
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1694700623
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_139
timestamp 1694700623
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_141
timestamp 1694700623
transform 1 0 17136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_144
timestamp 1694700623
transform 1 0 17472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_148
timestamp 1694700623
transform 1 0 17920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_152
timestamp 1694700623
transform 1 0 18368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_154
timestamp 1694700623
transform 1 0 18592 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_171
timestamp 1694700623
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1694700623
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1694700623
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_230
timestamp 1694700623
transform 1 0 27104 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1694700623
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1694700623
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_251
timestamp 1694700623
transform 1 0 29456 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_267
timestamp 1694700623
transform 1 0 31248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_272
timestamp 1694700623
transform 1 0 31808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_276
timestamp 1694700623
transform 1 0 32256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_284
timestamp 1694700623
transform 1 0 33152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_291
timestamp 1694700623
transform 1 0 33936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_299
timestamp 1694700623
transform 1 0 34832 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_303
timestamp 1694700623
transform 1 0 35280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1694700623
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1694700623
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1694700623
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1694700623
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_333
timestamp 1694700623
transform 1 0 38640 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_365
timestamp 1694700623
transform 1 0 42224 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1694700623
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1694700623
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_407
timestamp 1694700623
transform 1 0 46928 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_439
timestamp 1694700623
transform 1 0 50512 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_470
timestamp 1694700623
transform 1 0 53984 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_478
timestamp 1694700623
transform 1 0 54880 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_508
timestamp 1694700623
transform 1 0 58240 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1694700623
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_66
timestamp 1694700623
transform 1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1694700623
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_105
timestamp 1694700623
transform 1 0 13104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_109
timestamp 1694700623
transform 1 0 13552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_121
timestamp 1694700623
transform 1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_125
timestamp 1694700623
transform 1 0 15344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_129
timestamp 1694700623
transform 1 0 15792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_152
timestamp 1694700623
transform 1 0 18368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1694700623
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1694700623
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_162
timestamp 1694700623
transform 1 0 19488 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_200
timestamp 1694700623
transform 1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1694700623
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1694700623
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_217
timestamp 1694700623
transform 1 0 25648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_225
timestamp 1694700623
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_237
timestamp 1694700623
transform 1 0 27888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1694700623
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_253
timestamp 1694700623
transform 1 0 29680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_257
timestamp 1694700623
transform 1 0 30128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_265
timestamp 1694700623
transform 1 0 31024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_275
timestamp 1694700623
transform 1 0 32144 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1694700623
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_296
timestamp 1694700623
transform 1 0 34496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_300
timestamp 1694700623
transform 1 0 34944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_331
timestamp 1694700623
transform 1 0 38416 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_340
timestamp 1694700623
transform 1 0 39424 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1694700623
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_358
timestamp 1694700623
transform 1 0 41440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_360
timestamp 1694700623
transform 1 0 41664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_379
timestamp 1694700623
transform 1 0 43792 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_383
timestamp 1694700623
transform 1 0 44240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_386
timestamp 1694700623
transform 1 0 44576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_390
timestamp 1694700623
transform 1 0 45024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_394
timestamp 1694700623
transform 1 0 45472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_398
timestamp 1694700623
transform 1 0 45920 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_414
timestamp 1694700623
transform 1 0 47712 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_418
timestamp 1694700623
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_422
timestamp 1694700623
transform 1 0 48608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_426
timestamp 1694700623
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_467
timestamp 1694700623
transform 1 0 53648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_471
timestamp 1694700623
transform 1 0 54096 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_487
timestamp 1694700623
transform 1 0 55888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1694700623
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_506
timestamp 1694700623
transform 1 0 58016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1694700623
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1694700623
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1694700623
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_37
timestamp 1694700623
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_53
timestamp 1694700623
transform 1 0 7280 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_57
timestamp 1694700623
transform 1 0 7728 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_59
timestamp 1694700623
transform 1 0 7952 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_68
timestamp 1694700623
transform 1 0 8960 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_100
timestamp 1694700623
transform 1 0 12544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1694700623
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_107
timestamp 1694700623
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_121
timestamp 1694700623
transform 1 0 14896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1694700623
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_128
timestamp 1694700623
transform 1 0 15680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_168
timestamp 1694700623
transform 1 0 20160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1694700623
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1694700623
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1694700623
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_186
timestamp 1694700623
transform 1 0 22176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_190
timestamp 1694700623
transform 1 0 22624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_194
timestamp 1694700623
transform 1 0 23072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_197
timestamp 1694700623
transform 1 0 23408 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_210
timestamp 1694700623
transform 1 0 24864 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_214
timestamp 1694700623
transform 1 0 25312 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_238
timestamp 1694700623
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_242
timestamp 1694700623
transform 1 0 28448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_256
timestamp 1694700623
transform 1 0 30016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_260
timestamp 1694700623
transform 1 0 30464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_262
timestamp 1694700623
transform 1 0 30688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_269
timestamp 1694700623
transform 1 0 31472 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_287
timestamp 1694700623
transform 1 0 33488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_295
timestamp 1694700623
transform 1 0 34384 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_302
timestamp 1694700623
transform 1 0 35168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_309
timestamp 1694700623
transform 1 0 35952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1694700623
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_333
timestamp 1694700623
transform 1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_354
timestamp 1694700623
transform 1 0 40992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_356
timestamp 1694700623
transform 1 0 41216 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_365
timestamp 1694700623
transform 1 0 42224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_369
timestamp 1694700623
transform 1 0 42672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1694700623
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_375
timestamp 1694700623
transform 1 0 43344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1694700623
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_435
timestamp 1694700623
transform 1 0 50064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_439
timestamp 1694700623
transform 1 0 50512 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_470
timestamp 1694700623
transform 1 0 53984 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_486
timestamp 1694700623
transform 1 0 55776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_490
timestamp 1694700623
transform 1 0 56224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_496
timestamp 1694700623
transform 1 0 56896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_500
timestamp 1694700623
transform 1 0 57344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1694700623
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_34
timestamp 1694700623
transform 1 0 5152 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_38
timestamp 1694700623
transform 1 0 5600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1694700623
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1694700623
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1694700623
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_88
timestamp 1694700623
transform 1 0 11200 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_132
timestamp 1694700623
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_161
timestamp 1694700623
transform 1 0 19376 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_177
timestamp 1694700623
transform 1 0 21168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_185
timestamp 1694700623
transform 1 0 22064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1694700623
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1694700623
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_217
timestamp 1694700623
transform 1 0 25648 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_238
timestamp 1694700623
transform 1 0 28000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_254
timestamp 1694700623
transform 1 0 29792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_261
timestamp 1694700623
transform 1 0 30576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1694700623
transform 1 0 31024 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1694700623
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1694700623
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1694700623
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_282
timestamp 1694700623
transform 1 0 32928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1694700623
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_288
timestamp 1694700623
transform 1 0 33600 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_293
timestamp 1694700623
transform 1 0 34160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_297
timestamp 1694700623
transform 1 0 34608 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_313
timestamp 1694700623
transform 1 0 36400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_317
timestamp 1694700623
transform 1 0 36848 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_321
timestamp 1694700623
transform 1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_325
timestamp 1694700623
transform 1 0 37744 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_333
timestamp 1694700623
transform 1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_335
timestamp 1694700623
transform 1 0 38864 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1694700623
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_360
timestamp 1694700623
transform 1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_364
timestamp 1694700623
transform 1 0 42112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_395
timestamp 1694700623
transform 1 0 45584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_403
timestamp 1694700623
transform 1 0 46480 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_407
timestamp 1694700623
transform 1 0 46928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_415
timestamp 1694700623
transform 1 0 47824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1694700623
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_422
timestamp 1694700623
transform 1 0 48608 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_454
timestamp 1694700623
transform 1 0 52192 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_460
timestamp 1694700623
transform 1 0 52864 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_476
timestamp 1694700623
transform 1 0 54656 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_484
timestamp 1694700623
transform 1 0 55552 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1694700623
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_500
timestamp 1694700623
transform 1 0 57344 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_504
timestamp 1694700623
transform 1 0 57792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_506
timestamp 1694700623
transform 1 0 58016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1694700623
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1694700623
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1694700623
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_53
timestamp 1694700623
transform 1 0 7280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_61
timestamp 1694700623
transform 1 0 8176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_65
timestamp 1694700623
transform 1 0 8624 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_72
timestamp 1694700623
transform 1 0 9408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_76
timestamp 1694700623
transform 1 0 9856 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_92
timestamp 1694700623
transform 1 0 11648 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_96
timestamp 1694700623
transform 1 0 12096 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_123
timestamp 1694700623
transform 1 0 15120 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_139
timestamp 1694700623
transform 1 0 16912 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_147
timestamp 1694700623
transform 1 0 17808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_149
timestamp 1694700623
transform 1 0 18032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_152
timestamp 1694700623
transform 1 0 18368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_156
timestamp 1694700623
transform 1 0 18816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_160
timestamp 1694700623
transform 1 0 19264 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_163
timestamp 1694700623
transform 1 0 19600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1694700623
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1694700623
transform 1 0 21168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_193
timestamp 1694700623
transform 1 0 22960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_201
timestamp 1694700623
transform 1 0 23856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_210
timestamp 1694700623
transform 1 0 24864 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_229
timestamp 1694700623
transform 1 0 26992 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_237
timestamp 1694700623
transform 1 0 27888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_241
timestamp 1694700623
transform 1 0 28336 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1694700623
transform 1 0 29008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_249
timestamp 1694700623
transform 1 0 29232 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_252
timestamp 1694700623
transform 1 0 29568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_256
timestamp 1694700623
transform 1 0 30016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_260
timestamp 1694700623
transform 1 0 30464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_292
timestamp 1694700623
transform 1 0 34048 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_308
timestamp 1694700623
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1694700623
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1694700623
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1694700623
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_331
timestamp 1694700623
transform 1 0 38416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_335
timestamp 1694700623
transform 1 0 38864 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_343
timestamp 1694700623
transform 1 0 39760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_373
timestamp 1694700623
transform 1 0 43120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_377
timestamp 1694700623
transform 1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_395
timestamp 1694700623
transform 1 0 45584 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_427
timestamp 1694700623
transform 1 0 49168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_443
timestamp 1694700623
transform 1 0 50960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1694700623
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_470
timestamp 1694700623
transform 1 0 53984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_478
timestamp 1694700623
transform 1 0 54880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1694700623
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1694700623
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_26
timestamp 1694700623
transform 1 0 4256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_28
timestamp 1694700623
transform 1 0 4480 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_58
timestamp 1694700623
transform 1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_62
timestamp 1694700623
transform 1 0 8288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_110
timestamp 1694700623
transform 1 0 13664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_124
timestamp 1694700623
transform 1 0 15232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_132
timestamp 1694700623
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1694700623
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_152
timestamp 1694700623
transform 1 0 18368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_154
timestamp 1694700623
transform 1 0 18592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_190
timestamp 1694700623
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_194
timestamp 1694700623
transform 1 0 23072 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_244
timestamp 1694700623
transform 1 0 28672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_248
timestamp 1694700623
transform 1 0 29120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_256
timestamp 1694700623
transform 1 0 30016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_260
timestamp 1694700623
transform 1 0 30464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_272
timestamp 1694700623
transform 1 0 31808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_276
timestamp 1694700623
transform 1 0 32256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1694700623
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_290
timestamp 1694700623
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_294
timestamp 1694700623
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_303
timestamp 1694700623
transform 1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_305
timestamp 1694700623
transform 1 0 35504 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_312
timestamp 1694700623
transform 1 0 36288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_320
timestamp 1694700623
transform 1 0 37184 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_324
timestamp 1694700623
transform 1 0 37632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_342
timestamp 1694700623
transform 1 0 39648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_352
timestamp 1694700623
transform 1 0 40768 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_382
timestamp 1694700623
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_386
timestamp 1694700623
transform 1 0 44576 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_418
timestamp 1694700623
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_422
timestamp 1694700623
transform 1 0 48608 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_438
timestamp 1694700623
transform 1 0 50400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_442
timestamp 1694700623
transform 1 0 50848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_444
timestamp 1694700623
transform 1 0 51072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_474
timestamp 1694700623
transform 1 0 54432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_478
timestamp 1694700623
transform 1 0 54880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_485
timestamp 1694700623
transform 1 0 55664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_489
timestamp 1694700623
transform 1 0 56112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1694700623
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1694700623
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1694700623
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_37
timestamp 1694700623
transform 1 0 5488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_45
timestamp 1694700623
transform 1 0 6384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_49
timestamp 1694700623
transform 1 0 6832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_51
timestamp 1694700623
transform 1 0 7056 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_88
timestamp 1694700623
transform 1 0 11200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1694700623
transform 1 0 12768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1694700623
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1694700623
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_121
timestamp 1694700623
transform 1 0 14896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_125
timestamp 1694700623
transform 1 0 15344 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_165
timestamp 1694700623
transform 1 0 19824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1694700623
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_177
timestamp 1694700623
transform 1 0 21168 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_209
timestamp 1694700623
transform 1 0 24752 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_225
timestamp 1694700623
transform 1 0 26544 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_233
timestamp 1694700623
transform 1 0 27440 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1694700623
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1694700623
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_251
timestamp 1694700623
transform 1 0 29456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_255
timestamp 1694700623
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_257
timestamp 1694700623
transform 1 0 30128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_310
timestamp 1694700623
transform 1 0 36064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_312
timestamp 1694700623
transform 1 0 36288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_317
timestamp 1694700623
transform 1 0 36848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1694700623
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_360
timestamp 1694700623
transform 1 0 41664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_364
timestamp 1694700623
transform 1 0 42112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_368
timestamp 1694700623
transform 1 0 42560 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_379
timestamp 1694700623
transform 1 0 43792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1694700623
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_387
timestamp 1694700623
transform 1 0 44688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_391
timestamp 1694700623
transform 1 0 45136 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_423
timestamp 1694700623
transform 1 0 48720 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_427
timestamp 1694700623
transform 1 0 49168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_437
timestamp 1694700623
transform 1 0 50288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_441
timestamp 1694700623
transform 1 0 50736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_449
timestamp 1694700623
transform 1 0 51632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_453
timestamp 1694700623
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_468
timestamp 1694700623
transform 1 0 53760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_470
timestamp 1694700623
transform 1 0 53984 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_497
timestamp 1694700623
transform 1 0 57008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1694700623
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1694700623
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_18
timestamp 1694700623
transform 1 0 3360 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_22
timestamp 1694700623
transform 1 0 3808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_24
timestamp 1694700623
transform 1 0 4032 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_54
timestamp 1694700623
transform 1 0 7392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1694700623
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_127
timestamp 1694700623
transform 1 0 15568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_129
timestamp 1694700623
transform 1 0 15792 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_147
timestamp 1694700623
transform 1 0 17808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_151
timestamp 1694700623
transform 1 0 18256 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_167
timestamp 1694700623
transform 1 0 20048 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_171
timestamp 1694700623
transform 1 0 20496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_190
timestamp 1694700623
transform 1 0 22624 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_197
timestamp 1694700623
transform 1 0 23408 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_218
timestamp 1694700623
transform 1 0 25760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_226
timestamp 1694700623
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_240
timestamp 1694700623
transform 1 0 28224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_247
timestamp 1694700623
transform 1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_251
timestamp 1694700623
transform 1 0 29456 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_255
timestamp 1694700623
transform 1 0 29904 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_259
timestamp 1694700623
transform 1 0 30352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_270
timestamp 1694700623
transform 1 0 31584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_274
timestamp 1694700623
transform 1 0 32032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1694700623
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_282
timestamp 1694700623
transform 1 0 32928 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_298
timestamp 1694700623
transform 1 0 34720 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_302
timestamp 1694700623
transform 1 0 35168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_312
timestamp 1694700623
transform 1 0 36288 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_314
timestamp 1694700623
transform 1 0 36512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_323
timestamp 1694700623
transform 1 0 37520 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_339
timestamp 1694700623
transform 1 0 39312 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_343
timestamp 1694700623
transform 1 0 39760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1694700623
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_352
timestamp 1694700623
transform 1 0 40768 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_368
timestamp 1694700623
transform 1 0 42560 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_383
timestamp 1694700623
transform 1 0 44240 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_415
timestamp 1694700623
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1694700623
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_422
timestamp 1694700623
transform 1 0 48608 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_438
timestamp 1694700623
transform 1 0 50400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_450
timestamp 1694700623
transform 1 0 51744 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_458
timestamp 1694700623
transform 1 0 52640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_460
timestamp 1694700623
transform 1 0 52864 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_467
timestamp 1694700623
transform 1 0 53648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_471
timestamp 1694700623
transform 1 0 54096 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_487
timestamp 1694700623
transform 1 0 55888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_489
timestamp 1694700623
transform 1 0 56112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_492
timestamp 1694700623
transform 1 0 56448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_499
timestamp 1694700623
transform 1 0 57232 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_505
timestamp 1694700623
transform 1 0 57904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1694700623
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1694700623
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1694700623
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_121
timestamp 1694700623
transform 1 0 14896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_125
timestamp 1694700623
transform 1 0 15344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_129
timestamp 1694700623
transform 1 0 15792 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_145
timestamp 1694700623
transform 1 0 17584 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_153
timestamp 1694700623
transform 1 0 18480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_165
timestamp 1694700623
transform 1 0 19824 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_173
timestamp 1694700623
transform 1 0 20720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1694700623
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_189
timestamp 1694700623
transform 1 0 22512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_193
timestamp 1694700623
transform 1 0 22960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_201
timestamp 1694700623
transform 1 0 23856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_213
timestamp 1694700623
transform 1 0 25200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_215
timestamp 1694700623
transform 1 0 25424 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_262
timestamp 1694700623
transform 1 0 30688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_271
timestamp 1694700623
transform 1 0 31696 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_287
timestamp 1694700623
transform 1 0 33488 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_299
timestamp 1694700623
transform 1 0 34832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_309
timestamp 1694700623
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1694700623
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_346
timestamp 1694700623
transform 1 0 40096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_350
timestamp 1694700623
transform 1 0 40544 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1694700623
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1694700623
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_387
timestamp 1694700623
transform 1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_395
timestamp 1694700623
transform 1 0 45584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_399
timestamp 1694700623
transform 1 0 46032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_440
timestamp 1694700623
transform 1 0 50624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_444
timestamp 1694700623
transform 1 0 51072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_452
timestamp 1694700623
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1694700623
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_463
timestamp 1694700623
transform 1 0 53200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_471
timestamp 1694700623
transform 1 0 54096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_473
timestamp 1694700623
transform 1 0 54320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1694700623
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_34
timestamp 1694700623
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_50
timestamp 1694700623
transform 1 0 6944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_54
timestamp 1694700623
transform 1 0 7392 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1694700623
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_92
timestamp 1694700623
transform 1 0 11648 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_119
timestamp 1694700623
transform 1 0 14672 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_135
timestamp 1694700623
transform 1 0 16464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1694700623
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_142
timestamp 1694700623
transform 1 0 17248 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_174
timestamp 1694700623
transform 1 0 20832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_176
timestamp 1694700623
transform 1 0 21056 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_199
timestamp 1694700623
transform 1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1694700623
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1694700623
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_216
timestamp 1694700623
transform 1 0 25536 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_232
timestamp 1694700623
transform 1 0 27328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_234
timestamp 1694700623
transform 1 0 27552 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1694700623
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_282
timestamp 1694700623
transform 1 0 32928 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_298
timestamp 1694700623
transform 1 0 34720 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_301
timestamp 1694700623
transform 1 0 35056 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_310
timestamp 1694700623
transform 1 0 36064 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_342
timestamp 1694700623
transform 1 0 39648 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_352
timestamp 1694700623
transform 1 0 40768 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_360
timestamp 1694700623
transform 1 0 41664 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_393
timestamp 1694700623
transform 1 0 45360 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_397
timestamp 1694700623
transform 1 0 45808 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_413
timestamp 1694700623
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_417
timestamp 1694700623
transform 1 0 48048 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1694700623
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_422
timestamp 1694700623
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_424
timestamp 1694700623
transform 1 0 48832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_427
timestamp 1694700623
transform 1 0 49168 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_431
timestamp 1694700623
transform 1 0 49616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_438
timestamp 1694700623
transform 1 0 50400 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_470
timestamp 1694700623
transform 1 0 53984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1694700623
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1694700623
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_500
timestamp 1694700623
transform 1 0 57344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_502
timestamp 1694700623
transform 1 0 57568 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1694700623
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1694700623
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1694700623
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_53
timestamp 1694700623
transform 1 0 7280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_57
timestamp 1694700623
transform 1 0 7728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_73
timestamp 1694700623
transform 1 0 9520 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_92
timestamp 1694700623
transform 1 0 11648 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_102
timestamp 1694700623
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1694700623
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_120
timestamp 1694700623
transform 1 0 14784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_161
timestamp 1694700623
transform 1 0 19376 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_169
timestamp 1694700623
transform 1 0 20272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1694700623
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1694700623
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_193
timestamp 1694700623
transform 1 0 22960 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_197
timestamp 1694700623
transform 1 0 23408 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_199
timestamp 1694700623
transform 1 0 23632 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_229
timestamp 1694700623
transform 1 0 26992 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_233
timestamp 1694700623
transform 1 0 27440 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1694700623
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_247
timestamp 1694700623
transform 1 0 29008 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_263
timestamp 1694700623
transform 1 0 30800 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_296
timestamp 1694700623
transform 1 0 34496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_300
timestamp 1694700623
transform 1 0 34944 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_309
timestamp 1694700623
transform 1 0 35952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1694700623
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_329
timestamp 1694700623
transform 1 0 38192 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_362
timestamp 1694700623
transform 1 0 41888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_366
timestamp 1694700623
transform 1 0 42336 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_374
timestamp 1694700623
transform 1 0 43232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_376
timestamp 1694700623
transform 1 0 43456 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1694700623
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_391
timestamp 1694700623
transform 1 0 45136 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_421
timestamp 1694700623
transform 1 0 48496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_425
timestamp 1694700623
transform 1 0 48944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_443
timestamp 1694700623
transform 1 0 50960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1694700623
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_457
timestamp 1694700623
transform 1 0 52528 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_473
timestamp 1694700623
transform 1 0 54320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_477
timestamp 1694700623
transform 1 0 54768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_479
timestamp 1694700623
transform 1 0 54992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1694700623
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_34
timestamp 1694700623
transform 1 0 5152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_50
timestamp 1694700623
transform 1 0 6944 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_58
timestamp 1694700623
transform 1 0 7840 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_62
timestamp 1694700623
transform 1 0 8288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_91
timestamp 1694700623
transform 1 0 11536 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_106
timestamp 1694700623
transform 1 0 13216 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1694700623
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_142
timestamp 1694700623
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_150
timestamp 1694700623
transform 1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_152
timestamp 1694700623
transform 1 0 18368 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_159
timestamp 1694700623
transform 1 0 19152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_163
timestamp 1694700623
transform 1 0 19600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_167
timestamp 1694700623
transform 1 0 20048 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_170
timestamp 1694700623
transform 1 0 20384 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_208
timestamp 1694700623
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_212
timestamp 1694700623
transform 1 0 25088 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_228
timestamp 1694700623
transform 1 0 26880 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_236
timestamp 1694700623
transform 1 0 27776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_240
timestamp 1694700623
transform 1 0 28224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_242
timestamp 1694700623
transform 1 0 28448 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_245
timestamp 1694700623
transform 1 0 28784 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_261
timestamp 1694700623
transform 1 0 30576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_263
timestamp 1694700623
transform 1 0 30800 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1694700623
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_284
timestamp 1694700623
transform 1 0 33152 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1694700623
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_352
timestamp 1694700623
transform 1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1694700623
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_372
timestamp 1694700623
transform 1 0 43008 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_387
timestamp 1694700623
transform 1 0 44688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_391
timestamp 1694700623
transform 1 0 45136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_399
timestamp 1694700623
transform 1 0 46032 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_413
timestamp 1694700623
transform 1 0 47600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1694700623
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1694700623
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1694700623
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_432
timestamp 1694700623
transform 1 0 49728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_444
timestamp 1694700623
transform 1 0 51072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_446
timestamp 1694700623
transform 1 0 51296 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_449
timestamp 1694700623
transform 1 0 51632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_455
timestamp 1694700623
transform 1 0 52304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_465
timestamp 1694700623
transform 1 0 53424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_472
timestamp 1694700623
transform 1 0 54208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_482
timestamp 1694700623
transform 1 0 55328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_492
timestamp 1694700623
transform 1 0 56448 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_500
timestamp 1694700623
transform 1 0 57344 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_504
timestamp 1694700623
transform 1 0 57792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_506
timestamp 1694700623
transform 1 0 58016 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1694700623
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1694700623
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_37
timestamp 1694700623
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_69
timestamp 1694700623
transform 1 0 9072 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_85
timestamp 1694700623
transform 1 0 10864 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_89
timestamp 1694700623
transform 1 0 11312 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_115
timestamp 1694700623
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_119
timestamp 1694700623
transform 1 0 14672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_151
timestamp 1694700623
transform 1 0 18256 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_168
timestamp 1694700623
transform 1 0 20160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1694700623
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1694700623
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1694700623
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_210
timestamp 1694700623
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_220
timestamp 1694700623
transform 1 0 25984 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_228
timestamp 1694700623
transform 1 0 26880 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_232
timestamp 1694700623
transform 1 0 27328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1694700623
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_247
timestamp 1694700623
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_253
timestamp 1694700623
transform 1 0 29680 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_261
timestamp 1694700623
transform 1 0 30576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_309
timestamp 1694700623
transform 1 0 35952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1694700623
transform 1 0 36400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_325
timestamp 1694700623
transform 1 0 37744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_367
timestamp 1694700623
transform 1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_375
timestamp 1694700623
transform 1 0 43344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1694700623
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_387
timestamp 1694700623
transform 1 0 44688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_403
timestamp 1694700623
transform 1 0 46480 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_411
timestamp 1694700623
transform 1 0 47376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_415
timestamp 1694700623
transform 1 0 47824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_417
timestamp 1694700623
transform 1 0 48048 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_486
timestamp 1694700623
transform 1 0 55776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_490
timestamp 1694700623
transform 1 0 56224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_494
timestamp 1694700623
transform 1 0 56672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_505
timestamp 1694700623
transform 1 0 57904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1694700623
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_34
timestamp 1694700623
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_50
timestamp 1694700623
transform 1 0 6944 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_58
timestamp 1694700623
transform 1 0 7840 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_127
timestamp 1694700623
transform 1 0 15568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_135
timestamp 1694700623
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1694700623
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1694700623
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_144
timestamp 1694700623
transform 1 0 17472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_161
timestamp 1694700623
transform 1 0 19376 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_193
timestamp 1694700623
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_195
timestamp 1694700623
transform 1 0 23184 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_204
timestamp 1694700623
transform 1 0 24192 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_208
timestamp 1694700623
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1694700623
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_251
timestamp 1694700623
transform 1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_253
timestamp 1694700623
transform 1 0 29680 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_278
timestamp 1694700623
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_344
timestamp 1694700623
transform 1 0 39872 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_352
timestamp 1694700623
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_368
timestamp 1694700623
transform 1 0 42560 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_376
timestamp 1694700623
transform 1 0 43456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_387
timestamp 1694700623
transform 1 0 44688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_391
timestamp 1694700623
transform 1 0 45136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_393
timestamp 1694700623
transform 1 0 45360 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_412
timestamp 1694700623
transform 1 0 47488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1694700623
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_422
timestamp 1694700623
transform 1 0 48608 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_454
timestamp 1694700623
transform 1 0 52192 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_470
timestamp 1694700623
transform 1 0 53984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_474
timestamp 1694700623
transform 1 0 54432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_481
timestamp 1694700623
transform 1 0 55216 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_489
timestamp 1694700623
transform 1 0 56112 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_492
timestamp 1694700623
transform 1 0 56448 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_501
timestamp 1694700623
transform 1 0 57456 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1694700623
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_6
timestamp 1694700623
transform 1 0 2016 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_22
timestamp 1694700623
transform 1 0 3808 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_30
timestamp 1694700623
transform 1 0 4704 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1694700623
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1694700623
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_53
timestamp 1694700623
transform 1 0 7280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_97
timestamp 1694700623
transform 1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1694700623
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_117
timestamp 1694700623
transform 1 0 14448 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_125
timestamp 1694700623
transform 1 0 15344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_145
timestamp 1694700623
transform 1 0 17584 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_150
timestamp 1694700623
transform 1 0 18144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_168
timestamp 1694700623
transform 1 0 20160 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_172
timestamp 1694700623
transform 1 0 20608 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_206
timestamp 1694700623
transform 1 0 24416 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_222
timestamp 1694700623
transform 1 0 26208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_230
timestamp 1694700623
transform 1 0 27104 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_234
timestamp 1694700623
transform 1 0 27552 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1694700623
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1694700623
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1694700623
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_317
timestamp 1694700623
transform 1 0 36848 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_332
timestamp 1694700623
transform 1 0 38528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_336
timestamp 1694700623
transform 1 0 38976 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_368
timestamp 1694700623
transform 1 0 42560 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1694700623
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_392
timestamp 1694700623
transform 1 0 45248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_396
timestamp 1694700623
transform 1 0 45696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_427
timestamp 1694700623
transform 1 0 49168 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_432
timestamp 1694700623
transform 1 0 49728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_436
timestamp 1694700623
transform 1 0 50176 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1694700623
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1694700623
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_457
timestamp 1694700623
transform 1 0 52528 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_467
timestamp 1694700623
transform 1 0 53648 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_483
timestamp 1694700623
transform 1 0 55440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_491
timestamp 1694700623
transform 1 0 56336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_493
timestamp 1694700623
transform 1 0 56560 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_499
timestamp 1694700623
transform 1 0 57232 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_507
timestamp 1694700623
transform 1 0 58128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_10
timestamp 1694700623
transform 1 0 2464 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_42
timestamp 1694700623
transform 1 0 6048 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_58
timestamp 1694700623
transform 1 0 7840 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1694700623
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1694700623
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_88
timestamp 1694700623
transform 1 0 11200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_97
timestamp 1694700623
transform 1 0 12208 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_113
timestamp 1694700623
transform 1 0 14000 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_121
timestamp 1694700623
transform 1 0 14896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_123
timestamp 1694700623
transform 1 0 15120 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_134
timestamp 1694700623
transform 1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1694700623
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_176
timestamp 1694700623
transform 1 0 21056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_180
timestamp 1694700623
transform 1 0 21504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_188
timestamp 1694700623
transform 1 0 22400 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_198
timestamp 1694700623
transform 1 0 23520 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1694700623
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_220
timestamp 1694700623
transform 1 0 25984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1694700623
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_234
timestamp 1694700623
transform 1 0 27552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_238
timestamp 1694700623
transform 1 0 28000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_240
timestamp 1694700623
transform 1 0 28224 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_243
timestamp 1694700623
transform 1 0 28560 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_272
timestamp 1694700623
transform 1 0 31808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_274
timestamp 1694700623
transform 1 0 32032 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1694700623
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_284
timestamp 1694700623
transform 1 0 33152 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_311
timestamp 1694700623
transform 1 0 36176 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_315
timestamp 1694700623
transform 1 0 36624 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_341
timestamp 1694700623
transform 1 0 39536 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1694700623
transform 1 0 40432 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1694700623
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1694700623
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1694700623
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_397
timestamp 1694700623
transform 1 0 45808 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_413
timestamp 1694700623
transform 1 0 47600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1694700623
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1694700623
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_422
timestamp 1694700623
transform 1 0 48608 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_430
timestamp 1694700623
transform 1 0 49504 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_434
timestamp 1694700623
transform 1 0 49952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_442
timestamp 1694700623
transform 1 0 50848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_446
timestamp 1694700623
transform 1 0 51296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_448
timestamp 1694700623
transform 1 0 51520 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_455
timestamp 1694700623
transform 1 0 52304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_467
timestamp 1694700623
transform 1 0 53648 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_475
timestamp 1694700623
transform 1 0 54544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_477
timestamp 1694700623
transform 1 0 54768 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1694700623
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_507
timestamp 1694700623
transform 1 0 58128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_31
timestamp 1694700623
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1694700623
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_53
timestamp 1694700623
transform 1 0 7280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_61
timestamp 1694700623
transform 1 0 8176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_78
timestamp 1694700623
transform 1 0 10080 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_82
timestamp 1694700623
transform 1 0 10528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1694700623
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_123
timestamp 1694700623
transform 1 0 15120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_183
timestamp 1694700623
transform 1 0 21840 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_187
timestamp 1694700623
transform 1 0 22288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_196
timestamp 1694700623
transform 1 0 23296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_210
timestamp 1694700623
transform 1 0 24864 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_218
timestamp 1694700623
transform 1 0 25760 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_222
timestamp 1694700623
transform 1 0 26208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_224
timestamp 1694700623
transform 1 0 26432 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1694700623
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_247
timestamp 1694700623
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_255
timestamp 1694700623
transform 1 0 29904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_259
timestamp 1694700623
transform 1 0 30352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_294
timestamp 1694700623
transform 1 0 34272 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_296
timestamp 1694700623
transform 1 0 34496 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_312
timestamp 1694700623
transform 1 0 36288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1694700623
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_334
timestamp 1694700623
transform 1 0 38752 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_350
timestamp 1694700623
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_358
timestamp 1694700623
transform 1 0 41440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_362
timestamp 1694700623
transform 1 0 41888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_370
timestamp 1694700623
transform 1 0 42784 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_374
timestamp 1694700623
transform 1 0 43232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_376
timestamp 1694700623
transform 1 0 43456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1694700623
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_387
timestamp 1694700623
transform 1 0 44688 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_419
timestamp 1694700623
transform 1 0 48272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_423
timestamp 1694700623
transform 1 0 48720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_425
timestamp 1694700623
transform 1 0 48944 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_457
timestamp 1694700623
transform 1 0 52528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_461
timestamp 1694700623
transform 1 0 52976 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_491
timestamp 1694700623
transform 1 0 56336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_501
timestamp 1694700623
transform 1 0 57456 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1694700623
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_10
timestamp 1694700623
transform 1 0 2464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_56
timestamp 1694700623
transform 1 0 7616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_91
timestamp 1694700623
transform 1 0 11536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_106
timestamp 1694700623
transform 1 0 13216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_114
timestamp 1694700623
transform 1 0 14112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_118
timestamp 1694700623
transform 1 0 14560 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_155
timestamp 1694700623
transform 1 0 18704 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_179
timestamp 1694700623
transform 1 0 21392 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_183
timestamp 1694700623
transform 1 0 21840 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_218
timestamp 1694700623
transform 1 0 25760 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_256
timestamp 1694700623
transform 1 0 30016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_260
timestamp 1694700623
transform 1 0 30464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_269
timestamp 1694700623
transform 1 0 31472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_277
timestamp 1694700623
transform 1 0 32368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1694700623
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_330
timestamp 1694700623
transform 1 0 38304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_345
timestamp 1694700623
transform 1 0 39984 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1694700623
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_381
timestamp 1694700623
transform 1 0 44016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_385
timestamp 1694700623
transform 1 0 44464 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_401
timestamp 1694700623
transform 1 0 46256 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_408
timestamp 1694700623
transform 1 0 47040 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1694700623
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1694700623
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1694700623
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_492
timestamp 1694700623
transform 1 0 56448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_496
timestamp 1694700623
transform 1 0 56896 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_504
timestamp 1694700623
transform 1 0 57792 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1694700623
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2
timestamp 1694700623
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_18
timestamp 1694700623
transform 1 0 3360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_20
timestamp 1694700623
transform 1 0 3584 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_26
timestamp 1694700623
transform 1 0 4256 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_30
timestamp 1694700623
transform 1 0 4704 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1694700623
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1694700623
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_55
timestamp 1694700623
transform 1 0 7504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_63
timestamp 1694700623
transform 1 0 8400 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_79
timestamp 1694700623
transform 1 0 10192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1694700623
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_107
timestamp 1694700623
transform 1 0 13328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_142
timestamp 1694700623
transform 1 0 17248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_146
timestamp 1694700623
transform 1 0 17696 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_183
timestamp 1694700623
transform 1 0 21840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_187
timestamp 1694700623
transform 1 0 22288 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_195
timestamp 1694700623
transform 1 0 23184 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_199
timestamp 1694700623
transform 1 0 23632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_209
timestamp 1694700623
transform 1 0 24752 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_217
timestamp 1694700623
transform 1 0 25648 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_252
timestamp 1694700623
transform 1 0 29568 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_308
timestamp 1694700623
transform 1 0 35840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1694700623
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1694700623
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_330
timestamp 1694700623
transform 1 0 38304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_355
timestamp 1694700623
transform 1 0 41104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_357
timestamp 1694700623
transform 1 0 41328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_366
timestamp 1694700623
transform 1 0 42336 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1694700623
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1694700623
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_387
timestamp 1694700623
transform 1 0 44688 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_430
timestamp 1694700623
transform 1 0 49504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_434
timestamp 1694700623
transform 1 0 49952 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_450
timestamp 1694700623
transform 1 0 51744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1694700623
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1694700623
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_465
timestamp 1694700623
transform 1 0 53424 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_468
timestamp 1694700623
transform 1 0 53760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_476
timestamp 1694700623
transform 1 0 54656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1694700623
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_34
timestamp 1694700623
transform 1 0 5152 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_38
timestamp 1694700623
transform 1 0 5600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_40
timestamp 1694700623
transform 1 0 5824 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_62
timestamp 1694700623
transform 1 0 8288 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_72
timestamp 1694700623
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_80
timestamp 1694700623
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_84
timestamp 1694700623
transform 1 0 10752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_107
timestamp 1694700623
transform 1 0 13328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_115
timestamp 1694700623
transform 1 0 14224 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_119
timestamp 1694700623
transform 1 0 14672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1694700623
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1694700623
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1694700623
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_148
timestamp 1694700623
transform 1 0 17920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_176
timestamp 1694700623
transform 1 0 21056 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_192
timestamp 1694700623
transform 1 0 22848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_194
timestamp 1694700623
transform 1 0 23072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1694700623
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_240
timestamp 1694700623
transform 1 0 28224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_248
timestamp 1694700623
transform 1 0 29120 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_252
timestamp 1694700623
transform 1 0 29568 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1694700623
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1694700623
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_303
timestamp 1694700623
transform 1 0 35280 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_331
timestamp 1694700623
transform 1 0 38416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_352
timestamp 1694700623
transform 1 0 40768 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_384
timestamp 1694700623
transform 1 0 44352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_386
timestamp 1694700623
transform 1 0 44576 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_389
timestamp 1694700623
transform 1 0 44912 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_405
timestamp 1694700623
transform 1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_413
timestamp 1694700623
transform 1 0 47600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_417
timestamp 1694700623
transform 1 0 48048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1694700623
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_422
timestamp 1694700623
transform 1 0 48608 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_431
timestamp 1694700623
transform 1 0 49616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_464
timestamp 1694700623
transform 1 0 53312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_474
timestamp 1694700623
transform 1 0 54432 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_492
timestamp 1694700623
transform 1 0 56448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_496
timestamp 1694700623
transform 1 0 56896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_500
timestamp 1694700623
transform 1 0 57344 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_31
timestamp 1694700623
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_37
timestamp 1694700623
transform 1 0 5488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_45
timestamp 1694700623
transform 1 0 6384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_51
timestamp 1694700623
transform 1 0 7056 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_83
timestamp 1694700623
transform 1 0 10640 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_87
timestamp 1694700623
transform 1 0 11088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1694700623
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1694700623
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1694700623
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_165
timestamp 1694700623
transform 1 0 19824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_177
timestamp 1694700623
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_181
timestamp 1694700623
transform 1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_183
timestamp 1694700623
transform 1 0 21840 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_240
timestamp 1694700623
transform 1 0 28224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1694700623
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_247
timestamp 1694700623
transform 1 0 29008 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_263
timestamp 1694700623
transform 1 0 30800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_285
timestamp 1694700623
transform 1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_293
timestamp 1694700623
transform 1 0 34160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_295
timestamp 1694700623
transform 1 0 34384 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_304
timestamp 1694700623
transform 1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1694700623
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1694700623
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_317
timestamp 1694700623
transform 1 0 36848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_321
timestamp 1694700623
transform 1 0 37296 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_328
timestamp 1694700623
transform 1 0 38080 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_344
timestamp 1694700623
transform 1 0 39872 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_352
timestamp 1694700623
transform 1 0 40768 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_356
timestamp 1694700623
transform 1 0 41216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_358
timestamp 1694700623
transform 1 0 41440 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_367
timestamp 1694700623
transform 1 0 42448 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_371
timestamp 1694700623
transform 1 0 42896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1694700623
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_400
timestamp 1694700623
transform 1 0 46144 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_408
timestamp 1694700623
transform 1 0 47040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_414
timestamp 1694700623
transform 1 0 47712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_422
timestamp 1694700623
transform 1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_430
timestamp 1694700623
transform 1 0 49504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_434
timestamp 1694700623
transform 1 0 49952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_438
timestamp 1694700623
transform 1 0 50400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_448
timestamp 1694700623
transform 1 0 51520 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1694700623
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1694700623
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1694700623
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_506
timestamp 1694700623
transform 1 0 58016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_508
timestamp 1694700623
transform 1 0 58240 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_2
timestamp 1694700623
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_6
timestamp 1694700623
transform 1 0 2016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_37
timestamp 1694700623
transform 1 0 5488 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_53
timestamp 1694700623
transform 1 0 7280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_55
timestamp 1694700623
transform 1 0 7504 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_62
timestamp 1694700623
transform 1 0 8288 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_72
timestamp 1694700623
transform 1 0 9408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_104
timestamp 1694700623
transform 1 0 12992 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_112
timestamp 1694700623
transform 1 0 13888 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_115
timestamp 1694700623
transform 1 0 14224 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_119
timestamp 1694700623
transform 1 0 14672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_173
timestamp 1694700623
transform 1 0 20720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_177
timestamp 1694700623
transform 1 0 21168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_181
timestamp 1694700623
transform 1 0 21616 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_203
timestamp 1694700623
transform 1 0 24080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1694700623
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1694700623
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1694700623
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1694700623
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1694700623
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1694700623
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1694700623
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_290
timestamp 1694700623
transform 1 0 33824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_336
timestamp 1694700623
transform 1 0 38976 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_344
timestamp 1694700623
transform 1 0 39872 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_360
timestamp 1694700623
transform 1 0 41664 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_368
timestamp 1694700623
transform 1 0 42560 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_372
timestamp 1694700623
transform 1 0 43008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1694700623
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_422
timestamp 1694700623
transform 1 0 48608 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_438
timestamp 1694700623
transform 1 0 50400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_454
timestamp 1694700623
transform 1 0 52192 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_470
timestamp 1694700623
transform 1 0 53984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_478
timestamp 1694700623
transform 1 0 54880 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_482
timestamp 1694700623
transform 1 0 55328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_484
timestamp 1694700623
transform 1 0 55552 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_505
timestamp 1694700623
transform 1 0 57904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1694700623
transform 1 0 1568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_10
timestamp 1694700623
transform 1 0 2464 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_17
timestamp 1694700623
transform 1 0 3248 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_19
timestamp 1694700623
transform 1 0 3472 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_42
timestamp 1694700623
transform 1 0 6048 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_81
timestamp 1694700623
transform 1 0 10416 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_89
timestamp 1694700623
transform 1 0 11312 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_93
timestamp 1694700623
transform 1 0 11760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_95
timestamp 1694700623
transform 1 0 11984 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1694700623
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_114
timestamp 1694700623
transform 1 0 14112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_116
timestamp 1694700623
transform 1 0 14336 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1694700623
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_185
timestamp 1694700623
transform 1 0 22064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_189
timestamp 1694700623
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_191
timestamp 1694700623
transform 1 0 22736 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_202
timestamp 1694700623
transform 1 0 23968 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_220
timestamp 1694700623
transform 1 0 25984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_239
timestamp 1694700623
transform 1 0 28112 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_243
timestamp 1694700623
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_252
timestamp 1694700623
transform 1 0 29568 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_268
timestamp 1694700623
transform 1 0 31360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1694700623
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1694700623
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1694700623
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_333
timestamp 1694700623
transform 1 0 38640 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_341
timestamp 1694700623
transform 1 0 39536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_374
timestamp 1694700623
transform 1 0 43232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_378
timestamp 1694700623
transform 1 0 43680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1694700623
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1694700623
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_396
timestamp 1694700623
transform 1 0 45696 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_412
timestamp 1694700623
transform 1 0 47488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_428
timestamp 1694700623
transform 1 0 49280 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_442
timestamp 1694700623
transform 1 0 50848 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_446
timestamp 1694700623
transform 1 0 51296 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_467
timestamp 1694700623
transform 1 0 53648 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_475
timestamp 1694700623
transform 1 0 54544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_2
timestamp 1694700623
transform 1 0 1568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_10
timestamp 1694700623
transform 1 0 2464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_14
timestamp 1694700623
transform 1 0 2912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_16
timestamp 1694700623
transform 1 0 3136 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_19
timestamp 1694700623
transform 1 0 3472 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_27
timestamp 1694700623
transform 1 0 4368 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_31
timestamp 1694700623
transform 1 0 4816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_33
timestamp 1694700623
transform 1 0 5040 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_63
timestamp 1694700623
transform 1 0 8400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_77
timestamp 1694700623
transform 1 0 9968 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_81
timestamp 1694700623
transform 1 0 10416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_83
timestamp 1694700623
transform 1 0 10640 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_121
timestamp 1694700623
transform 1 0 14896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_123
timestamp 1694700623
transform 1 0 15120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_142
timestamp 1694700623
transform 1 0 17248 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_186
timestamp 1694700623
transform 1 0 22176 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_194
timestamp 1694700623
transform 1 0 23072 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_261
timestamp 1694700623
transform 1 0 30576 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_277
timestamp 1694700623
transform 1 0 32368 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1694700623
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_284
timestamp 1694700623
transform 1 0 33152 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_310
timestamp 1694700623
transform 1 0 36064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_343
timestamp 1694700623
transform 1 0 39760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_347
timestamp 1694700623
transform 1 0 40208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1694700623
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_362
timestamp 1694700623
transform 1 0 41888 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_370
timestamp 1694700623
transform 1 0 42784 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_374
timestamp 1694700623
transform 1 0 43232 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_381
timestamp 1694700623
transform 1 0 44016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_387
timestamp 1694700623
transform 1 0 44688 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1694700623
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_422
timestamp 1694700623
transform 1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_424
timestamp 1694700623
transform 1 0 48832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_454
timestamp 1694700623
transform 1 0 52192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_458
timestamp 1694700623
transform 1 0 52640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_489
timestamp 1694700623
transform 1 0 56112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_492
timestamp 1694700623
transform 1 0 56448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_504
timestamp 1694700623
transform 1 0 57792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_506
timestamp 1694700623
transform 1 0 58016 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1694700623
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_10
timestamp 1694700623
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_12
timestamp 1694700623
transform 1 0 2688 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_25
timestamp 1694700623
transform 1 0 4144 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1694700623
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1694700623
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_53
timestamp 1694700623
transform 1 0 7280 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_61
timestamp 1694700623
transform 1 0 8176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_71
timestamp 1694700623
transform 1 0 9296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_87
timestamp 1694700623
transform 1 0 11088 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_120
timestamp 1694700623
transform 1 0 14784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_177
timestamp 1694700623
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_181
timestamp 1694700623
transform 1 0 21616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_187
timestamp 1694700623
transform 1 0 22288 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_203
timestamp 1694700623
transform 1 0 24080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_207
timestamp 1694700623
transform 1 0 24528 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_225
timestamp 1694700623
transform 1 0 26544 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_237
timestamp 1694700623
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_239
timestamp 1694700623
transform 1 0 28112 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_269
timestamp 1694700623
transform 1 0 31472 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_277
timestamp 1694700623
transform 1 0 32368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_281
timestamp 1694700623
transform 1 0 32816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_285
timestamp 1694700623
transform 1 0 33264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_289
timestamp 1694700623
transform 1 0 33712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_293
timestamp 1694700623
transform 1 0 34160 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_309
timestamp 1694700623
transform 1 0 35952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_335
timestamp 1694700623
transform 1 0 38864 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_348
timestamp 1694700623
transform 1 0 40320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_352
timestamp 1694700623
transform 1 0 40768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_387
timestamp 1694700623
transform 1 0 44688 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_398
timestamp 1694700623
transform 1 0 45920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_408
timestamp 1694700623
transform 1 0 47040 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_424
timestamp 1694700623
transform 1 0 48832 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_428
timestamp 1694700623
transform 1 0 49280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_430
timestamp 1694700623
transform 1 0 49504 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_438
timestamp 1694700623
transform 1 0 50400 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_446
timestamp 1694700623
transform 1 0 51296 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1694700623
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_457
timestamp 1694700623
transform 1 0 52528 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_461
timestamp 1694700623
transform 1 0 52976 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_35
timestamp 1694700623
transform 1 0 5264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_39
timestamp 1694700623
transform 1 0 5712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_55
timestamp 1694700623
transform 1 0 7504 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_63
timestamp 1694700623
transform 1 0 8400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1694700623
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1694700623
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_72
timestamp 1694700623
transform 1 0 9408 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_104
timestamp 1694700623
transform 1 0 12992 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_120
timestamp 1694700623
transform 1 0 14784 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_124
timestamp 1694700623
transform 1 0 15232 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_130
timestamp 1694700623
transform 1 0 15904 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1694700623
transform 1 0 16688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1694700623
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_142
timestamp 1694700623
transform 1 0 17248 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_193
timestamp 1694700623
transform 1 0 22960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_197
timestamp 1694700623
transform 1 0 23408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_205
timestamp 1694700623
transform 1 0 24304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1694700623
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_212
timestamp 1694700623
transform 1 0 25088 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_244
timestamp 1694700623
transform 1 0 28672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_260
timestamp 1694700623
transform 1 0 30464 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_268
timestamp 1694700623
transform 1 0 31360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_270
timestamp 1694700623
transform 1 0 31584 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1694700623
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_282
timestamp 1694700623
transform 1 0 32928 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1694700623
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_382
timestamp 1694700623
transform 1 0 44128 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_386
timestamp 1694700623
transform 1 0 44576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_388
timestamp 1694700623
transform 1 0 44800 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_422
timestamp 1694700623
transform 1 0 48608 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_454
timestamp 1694700623
transform 1 0 52192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_458
timestamp 1694700623
transform 1 0 52640 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_487
timestamp 1694700623
transform 1 0 55888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1694700623
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_492
timestamp 1694700623
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_502
timestamp 1694700623
transform 1 0 57568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_506
timestamp 1694700623
transform 1 0 58016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1694700623
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_2
timestamp 1694700623
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_6
timestamp 1694700623
transform 1 0 2016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_8
timestamp 1694700623
transform 1 0 2240 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_15
timestamp 1694700623
transform 1 0 3024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_45
timestamp 1694700623
transform 1 0 6384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_49
timestamp 1694700623
transform 1 0 6832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_71
timestamp 1694700623
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_75
timestamp 1694700623
transform 1 0 9744 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_91
timestamp 1694700623
transform 1 0 11536 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_99
timestamp 1694700623
transform 1 0 12432 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_103
timestamp 1694700623
transform 1 0 12880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_113
timestamp 1694700623
transform 1 0 14000 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_121
timestamp 1694700623
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_197
timestamp 1694700623
transform 1 0 23408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_201
timestamp 1694700623
transform 1 0 23856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_211
timestamp 1694700623
transform 1 0 24976 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_221
timestamp 1694700623
transform 1 0 26096 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_237
timestamp 1694700623
transform 1 0 27888 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_247
timestamp 1694700623
transform 1 0 29008 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_263
timestamp 1694700623
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_285
timestamp 1694700623
transform 1 0 33264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_287
timestamp 1694700623
transform 1 0 33488 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_304
timestamp 1694700623
transform 1 0 35392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_308
timestamp 1694700623
transform 1 0 35840 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1694700623
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1694700623
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1694700623
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_327
timestamp 1694700623
transform 1 0 37968 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_343
timestamp 1694700623
transform 1 0 39760 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_347
timestamp 1694700623
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_349
timestamp 1694700623
transform 1 0 40432 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1694700623
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_410
timestamp 1694700623
transform 1 0 47264 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_457
timestamp 1694700623
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_465
timestamp 1694700623
transform 1 0 53424 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_469
timestamp 1694700623
transform 1 0 53872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_485
timestamp 1694700623
transform 1 0 55664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_487
timestamp 1694700623
transform 1 0 55888 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_498
timestamp 1694700623
transform 1 0 57120 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_504
timestamp 1694700623
transform 1 0 57792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_506
timestamp 1694700623
transform 1 0 58016 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_2
timestamp 1694700623
transform 1 0 1568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_10
timestamp 1694700623
transform 1 0 2464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_14
timestamp 1694700623
transform 1 0 2912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_17
timestamp 1694700623
transform 1 0 3248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_25
timestamp 1694700623
transform 1 0 4144 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_29
timestamp 1694700623
transform 1 0 4592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_35
timestamp 1694700623
transform 1 0 5264 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_39
timestamp 1694700623
transform 1 0 5712 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1694700623
transform 1 0 9072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_80
timestamp 1694700623
transform 1 0 10304 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_112
timestamp 1694700623
transform 1 0 13888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_114
timestamp 1694700623
transform 1 0 14112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_131
timestamp 1694700623
transform 1 0 16016 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1694700623
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_142
timestamp 1694700623
transform 1 0 17248 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_174
timestamp 1694700623
transform 1 0 20832 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_177
timestamp 1694700623
transform 1 0 21168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_179
timestamp 1694700623
transform 1 0 21392 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_201
timestamp 1694700623
transform 1 0 23856 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_224
timestamp 1694700623
transform 1 0 26432 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_246
timestamp 1694700623
transform 1 0 28896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_250
timestamp 1694700623
transform 1 0 29344 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_266
timestamp 1694700623
transform 1 0 31136 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1694700623
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_313
timestamp 1694700623
transform 1 0 36400 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_317
timestamp 1694700623
transform 1 0 36848 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_325
timestamp 1694700623
transform 1 0 37744 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_329
timestamp 1694700623
transform 1 0 38192 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_332
timestamp 1694700623
transform 1 0 38528 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_348
timestamp 1694700623
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_352
timestamp 1694700623
transform 1 0 40768 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_368
timestamp 1694700623
transform 1 0 42560 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_376
timestamp 1694700623
transform 1 0 43456 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_378
timestamp 1694700623
transform 1 0 43680 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_381
timestamp 1694700623
transform 1 0 44016 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_413
timestamp 1694700623
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_417
timestamp 1694700623
transform 1 0 48048 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_428
timestamp 1694700623
transform 1 0 49280 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_432
timestamp 1694700623
transform 1 0 49728 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_462
timestamp 1694700623
transform 1 0 53088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_466
timestamp 1694700623
transform 1 0 53536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_474
timestamp 1694700623
transform 1 0 54432 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_478
timestamp 1694700623
transform 1 0 54880 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_500
timestamp 1694700623
transform 1 0 57344 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_2
timestamp 1694700623
transform 1 0 1568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_10
timestamp 1694700623
transform 1 0 2464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_16
timestamp 1694700623
transform 1 0 3136 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_32
timestamp 1694700623
transform 1 0 4928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1694700623
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_37
timestamp 1694700623
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_53
timestamp 1694700623
transform 1 0 7280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_57
timestamp 1694700623
transform 1 0 7728 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_66
timestamp 1694700623
transform 1 0 8736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1694700623
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_111
timestamp 1694700623
transform 1 0 13776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_130
timestamp 1694700623
transform 1 0 15904 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_138
timestamp 1694700623
transform 1 0 16800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_155
timestamp 1694700623
transform 1 0 18704 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_163
timestamp 1694700623
transform 1 0 19600 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1694700623
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_181
timestamp 1694700623
transform 1 0 21616 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_189
timestamp 1694700623
transform 1 0 22512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_195
timestamp 1694700623
transform 1 0 23184 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_227
timestamp 1694700623
transform 1 0 26768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_241
timestamp 1694700623
transform 1 0 28336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_262
timestamp 1694700623
transform 1 0 30688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_293
timestamp 1694700623
transform 1 0 34160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_297
timestamp 1694700623
transform 1 0 34608 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1694700623
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_317
timestamp 1694700623
transform 1 0 36848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_321
timestamp 1694700623
transform 1 0 37296 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_330
timestamp 1694700623
transform 1 0 38304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_332
timestamp 1694700623
transform 1 0 38528 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_362
timestamp 1694700623
transform 1 0 41888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_366
timestamp 1694700623
transform 1 0 42336 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_382
timestamp 1694700623
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1694700623
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_387
timestamp 1694700623
transform 1 0 44688 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_396
timestamp 1694700623
transform 1 0 45696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_400
timestamp 1694700623
transform 1 0 46144 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_422
timestamp 1694700623
transform 1 0 48608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_432
timestamp 1694700623
transform 1 0 49728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_436
timestamp 1694700623
transform 1 0 50176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_438
timestamp 1694700623
transform 1 0 50400 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_447
timestamp 1694700623
transform 1 0 51408 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_457
timestamp 1694700623
transform 1 0 52528 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_473
timestamp 1694700623
transform 1 0 54320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_477
timestamp 1694700623
transform 1 0 54768 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2
timestamp 1694700623
transform 1 0 1568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_6
timestamp 1694700623
transform 1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_14
timestamp 1694700623
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_16
timestamp 1694700623
transform 1 0 3136 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_40
timestamp 1694700623
transform 1 0 5824 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_56
timestamp 1694700623
transform 1 0 7616 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_64
timestamp 1694700623
transform 1 0 8512 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1694700623
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_105
timestamp 1694700623
transform 1 0 13104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_127
timestamp 1694700623
transform 1 0 15568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_135
timestamp 1694700623
transform 1 0 16464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1694700623
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_142
timestamp 1694700623
transform 1 0 17248 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_167
timestamp 1694700623
transform 1 0 20048 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_183
timestamp 1694700623
transform 1 0 21840 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_191
timestamp 1694700623
transform 1 0 22736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_195
timestamp 1694700623
transform 1 0 23184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_212
timestamp 1694700623
transform 1 0 25088 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_216
timestamp 1694700623
transform 1 0 25536 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_236
timestamp 1694700623
transform 1 0 27776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_240
timestamp 1694700623
transform 1 0 28224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_276
timestamp 1694700623
transform 1 0 32256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_282
timestamp 1694700623
transform 1 0 32928 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_290
timestamp 1694700623
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_294
timestamp 1694700623
transform 1 0 34272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_296
timestamp 1694700623
transform 1 0 34496 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_305
timestamp 1694700623
transform 1 0 35504 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1694700623
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_358
timestamp 1694700623
transform 1 0 41440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_362
timestamp 1694700623
transform 1 0 41888 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_378
timestamp 1694700623
transform 1 0 43680 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_382
timestamp 1694700623
transform 1 0 44128 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_403
timestamp 1694700623
transform 1 0 46480 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_411
timestamp 1694700623
transform 1 0 47376 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_446
timestamp 1694700623
transform 1 0 51296 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_454
timestamp 1694700623
transform 1 0 52192 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_458
timestamp 1694700623
transform 1 0 52640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_460
timestamp 1694700623
transform 1 0 52864 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_469
timestamp 1694700623
transform 1 0 53872 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_483
timestamp 1694700623
transform 1 0 55440 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_487
timestamp 1694700623
transform 1 0 55888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_489
timestamp 1694700623
transform 1 0 56112 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1694700623
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1694700623
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1694700623
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_43
timestamp 1694700623
transform 1 0 6160 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_75
timestamp 1694700623
transform 1 0 9744 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1694700623
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_107
timestamp 1694700623
transform 1 0 13328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_109
timestamp 1694700623
transform 1 0 13552 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_116
timestamp 1694700623
transform 1 0 14336 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_132
timestamp 1694700623
transform 1 0 16128 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_140
timestamp 1694700623
transform 1 0 17024 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_153
timestamp 1694700623
transform 1 0 18480 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_169
timestamp 1694700623
transform 1 0 20272 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_173
timestamp 1694700623
transform 1 0 20720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_177
timestamp 1694700623
transform 1 0 21168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_185
timestamp 1694700623
transform 1 0 22064 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_212
timestamp 1694700623
transform 1 0 25088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1694700623
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1694700623
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_255
timestamp 1694700623
transform 1 0 29904 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_287
timestamp 1694700623
transform 1 0 33488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_291
timestamp 1694700623
transform 1 0 33936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_293
timestamp 1694700623
transform 1 0 34160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_307
timestamp 1694700623
transform 1 0 35728 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_343
timestamp 1694700623
transform 1 0 39760 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_351
timestamp 1694700623
transform 1 0 40656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_376
timestamp 1694700623
transform 1 0 43456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_380
timestamp 1694700623
transform 1 0 43904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_382
timestamp 1694700623
transform 1 0 44128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_416
timestamp 1694700623
transform 1 0 47936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_422
timestamp 1694700623
transform 1 0 48608 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_430
timestamp 1694700623
transform 1 0 49504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_434
timestamp 1694700623
transform 1 0 49952 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_450
timestamp 1694700623
transform 1 0 51744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1694700623
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_488
timestamp 1694700623
transform 1 0 56000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_492
timestamp 1694700623
transform 1 0 56448 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_508
timestamp 1694700623
transform 1 0 58240 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_2
timestamp 1694700623
transform 1 0 1568 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_18
timestamp 1694700623
transform 1 0 3360 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_22
timestamp 1694700623
transform 1 0 3808 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_24
timestamp 1694700623
transform 1 0 4032 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_45
timestamp 1694700623
transform 1 0 6384 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_53
timestamp 1694700623
transform 1 0 7280 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_57
timestamp 1694700623
transform 1 0 7728 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_72
timestamp 1694700623
transform 1 0 9408 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_76
timestamp 1694700623
transform 1 0 9856 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_101
timestamp 1694700623
transform 1 0 12656 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_103
timestamp 1694700623
transform 1 0 12880 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_106
timestamp 1694700623
transform 1 0 13216 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_133
timestamp 1694700623
transform 1 0 16240 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_137
timestamp 1694700623
transform 1 0 16688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1694700623
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_142
timestamp 1694700623
transform 1 0 17248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_172
timestamp 1694700623
transform 1 0 20608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_174
timestamp 1694700623
transform 1 0 20832 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_177
timestamp 1694700623
transform 1 0 21168 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_212
timestamp 1694700623
transform 1 0 25088 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_228
timestamp 1694700623
transform 1 0 26880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_238
timestamp 1694700623
transform 1 0 28000 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_270
timestamp 1694700623
transform 1 0 31584 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_274
timestamp 1694700623
transform 1 0 32032 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_276
timestamp 1694700623
transform 1 0 32256 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1694700623
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_282
timestamp 1694700623
transform 1 0 32928 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_298
timestamp 1694700623
transform 1 0 34720 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_306
timestamp 1694700623
transform 1 0 35616 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_308
timestamp 1694700623
transform 1 0 35840 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_324
timestamp 1694700623
transform 1 0 37632 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_340
timestamp 1694700623
transform 1 0 39424 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_348
timestamp 1694700623
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_352
timestamp 1694700623
transform 1 0 40768 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_356
timestamp 1694700623
transform 1 0 41216 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_362
timestamp 1694700623
transform 1 0 41888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_364
timestamp 1694700623
transform 1 0 42112 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_370
timestamp 1694700623
transform 1 0 42784 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_372
timestamp 1694700623
transform 1 0 43008 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_381
timestamp 1694700623
transform 1 0 44016 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_413
timestamp 1694700623
transform 1 0 47600 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_417
timestamp 1694700623
transform 1 0 48048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1694700623
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_422
timestamp 1694700623
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_438
timestamp 1694700623
transform 1 0 50400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_440
timestamp 1694700623
transform 1 0 50624 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_470
timestamp 1694700623
transform 1 0 53984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_474
timestamp 1694700623
transform 1 0 54432 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_480
timestamp 1694700623
transform 1 0 55104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1694700623
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1694700623
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1694700623
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1694700623
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_37
timestamp 1694700623
transform 1 0 5488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_39
timestamp 1694700623
transform 1 0 5712 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_77
timestamp 1694700623
transform 1 0 9968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_81
timestamp 1694700623
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_85
timestamp 1694700623
transform 1 0 10864 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_92
timestamp 1694700623
transform 1 0 11648 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_100
timestamp 1694700623
transform 1 0 12544 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_104
timestamp 1694700623
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_107
timestamp 1694700623
transform 1 0 13328 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_164
timestamp 1694700623
transform 1 0 19712 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1694700623
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_185
timestamp 1694700623
transform 1 0 22064 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_220
timestamp 1694700623
transform 1 0 25984 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_236
timestamp 1694700623
transform 1 0 27776 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1694700623
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_247
timestamp 1694700623
transform 1 0 29008 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_263
timestamp 1694700623
transform 1 0 30800 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_265
timestamp 1694700623
transform 1 0 31024 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_287
timestamp 1694700623
transform 1 0 33488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_291
timestamp 1694700623
transform 1 0 33936 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_307
timestamp 1694700623
transform 1 0 35728 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_317
timestamp 1694700623
transform 1 0 36848 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_349
timestamp 1694700623
transform 1 0 40432 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_357
timestamp 1694700623
transform 1 0 41328 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_359
timestamp 1694700623
transform 1 0 41552 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_369
timestamp 1694700623
transform 1 0 42672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_375
timestamp 1694700623
transform 1 0 43344 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_383
timestamp 1694700623
transform 1 0 44240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_387
timestamp 1694700623
transform 1 0 44688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_403
timestamp 1694700623
transform 1 0 46480 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_433
timestamp 1694700623
transform 1 0 49840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_435
timestamp 1694700623
transform 1 0 50064 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_446
timestamp 1694700623
transform 1 0 51296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_450
timestamp 1694700623
transform 1 0 51744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_452
timestamp 1694700623
transform 1 0 51968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_465
timestamp 1694700623
transform 1 0 53424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_467
timestamp 1694700623
transform 1 0 53648 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_2
timestamp 1694700623
transform 1 0 1568 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_10
timestamp 1694700623
transform 1 0 2464 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_34
timestamp 1694700623
transform 1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_38
timestamp 1694700623
transform 1 0 5600 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_54
timestamp 1694700623
transform 1 0 7392 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_82
timestamp 1694700623
transform 1 0 10528 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_108
timestamp 1694700623
transform 1 0 13440 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_122
timestamp 1694700623
transform 1 0 15008 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_138
timestamp 1694700623
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_142
timestamp 1694700623
transform 1 0 17248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_183
timestamp 1694700623
transform 1 0 21840 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_191
timestamp 1694700623
transform 1 0 22736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_195
timestamp 1694700623
transform 1 0 23184 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_202
timestamp 1694700623
transform 1 0 23968 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_212
timestamp 1694700623
transform 1 0 25088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_228
timestamp 1694700623
transform 1 0 26880 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_236
timestamp 1694700623
transform 1 0 27776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_258
timestamp 1694700623
transform 1 0 30240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_262
timestamp 1694700623
transform 1 0 30688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_294
timestamp 1694700623
transform 1 0 34272 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_306
timestamp 1694700623
transform 1 0 35616 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_314
timestamp 1694700623
transform 1 0 36512 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_341
timestamp 1694700623
transform 1 0 39536 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1694700623
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_366
timestamp 1694700623
transform 1 0 42336 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_398
timestamp 1694700623
transform 1 0 45920 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_406
timestamp 1694700623
transform 1 0 46816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_408
timestamp 1694700623
transform 1 0 47040 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_413
timestamp 1694700623
transform 1 0 47600 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1694700623
transform 1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1694700623
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_422
timestamp 1694700623
transform 1 0 48608 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_430
timestamp 1694700623
transform 1 0 49504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_432
timestamp 1694700623
transform 1 0 49728 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_435
timestamp 1694700623
transform 1 0 50064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_437
timestamp 1694700623
transform 1 0 50288 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_445
timestamp 1694700623
transform 1 0 51184 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_459
timestamp 1694700623
transform 1 0 52752 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_475
timestamp 1694700623
transform 1 0 54544 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_483
timestamp 1694700623
transform 1 0 55440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_487
timestamp 1694700623
transform 1 0 55888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_489
timestamp 1694700623
transform 1 0 56112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1694700623
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1694700623
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_42
timestamp 1694700623
transform 1 0 6048 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_58
timestamp 1694700623
transform 1 0 7840 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_62
timestamp 1694700623
transform 1 0 8288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_64
timestamp 1694700623
transform 1 0 8512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_80
timestamp 1694700623
transform 1 0 10304 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_94
timestamp 1694700623
transform 1 0 11872 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_102
timestamp 1694700623
transform 1 0 12768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_104
timestamp 1694700623
transform 1 0 12992 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_107
timestamp 1694700623
transform 1 0 13328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_109
timestamp 1694700623
transform 1 0 13552 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_118
timestamp 1694700623
transform 1 0 14560 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_150
timestamp 1694700623
transform 1 0 18144 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_158
timestamp 1694700623
transform 1 0 19040 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_166
timestamp 1694700623
transform 1 0 19936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1694700623
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_177
timestamp 1694700623
transform 1 0 21168 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_209
timestamp 1694700623
transform 1 0 24752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_211
timestamp 1694700623
transform 1 0 24976 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_243
timestamp 1694700623
transform 1 0 28560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_267
timestamp 1694700623
transform 1 0 31248 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_271
timestamp 1694700623
transform 1 0 31696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_273
timestamp 1694700623
transform 1 0 31920 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_289
timestamp 1694700623
transform 1 0 33712 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_293
timestamp 1694700623
transform 1 0 34160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_295
timestamp 1694700623
transform 1 0 34384 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1694700623
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_317
timestamp 1694700623
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_325
timestamp 1694700623
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_329
timestamp 1694700623
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_368
timestamp 1694700623
transform 1 0 42560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_372
timestamp 1694700623
transform 1 0 43008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_380
timestamp 1694700623
transform 1 0 43904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1694700623
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_395
timestamp 1694700623
transform 1 0 45584 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_399
timestamp 1694700623
transform 1 0 46032 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_403
timestamp 1694700623
transform 1 0 46480 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_413
timestamp 1694700623
transform 1 0 47600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_417
timestamp 1694700623
transform 1 0 48048 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_449
timestamp 1694700623
transform 1 0 51632 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_453
timestamp 1694700623
transform 1 0 52080 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_457
timestamp 1694700623
transform 1 0 52528 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_473
timestamp 1694700623
transform 1 0 54320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_477
timestamp 1694700623
transform 1 0 54768 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_2
timestamp 1694700623
transform 1 0 1568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_10
timestamp 1694700623
transform 1 0 2464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_14
timestamp 1694700623
transform 1 0 2912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_44
timestamp 1694700623
transform 1 0 6272 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_60
timestamp 1694700623
transform 1 0 8064 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1694700623
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_72
timestamp 1694700623
transform 1 0 9408 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_88
timestamp 1694700623
transform 1 0 11200 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_96
timestamp 1694700623
transform 1 0 12096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_100
timestamp 1694700623
transform 1 0 12544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_109
timestamp 1694700623
transform 1 0 13552 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_117
timestamp 1694700623
transform 1 0 14448 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_126
timestamp 1694700623
transform 1 0 15456 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_134
timestamp 1694700623
transform 1 0 16352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_138
timestamp 1694700623
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1694700623
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1694700623
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_212
timestamp 1694700623
transform 1 0 25088 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_228
timestamp 1694700623
transform 1 0 26880 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_236
timestamp 1694700623
transform 1 0 27776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_259
timestamp 1694700623
transform 1 0 30352 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_275
timestamp 1694700623
transform 1 0 32144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1694700623
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_282
timestamp 1694700623
transform 1 0 32928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_298
timestamp 1694700623
transform 1 0 34720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_306
timestamp 1694700623
transform 1 0 35616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_335
timestamp 1694700623
transform 1 0 38864 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_343
timestamp 1694700623
transform 1 0 39760 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_347
timestamp 1694700623
transform 1 0 40208 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1694700623
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_363
timestamp 1694700623
transform 1 0 42000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_367
timestamp 1694700623
transform 1 0 42448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_371
timestamp 1694700623
transform 1 0 42896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_373
timestamp 1694700623
transform 1 0 43120 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_405
timestamp 1694700623
transform 1 0 46704 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_426
timestamp 1694700623
transform 1 0 49056 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_442
timestamp 1694700623
transform 1 0 50848 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_446
timestamp 1694700623
transform 1 0 51296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_448
timestamp 1694700623
transform 1 0 51520 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_465
timestamp 1694700623
transform 1 0 53424 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_473
timestamp 1694700623
transform 1 0 54320 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_477
timestamp 1694700623
transform 1 0 54768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_489
timestamp 1694700623
transform 1 0 56112 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_500
timestamp 1694700623
transform 1 0 57344 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1694700623
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_2
timestamp 1694700623
transform 1 0 1568 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_18
timestamp 1694700623
transform 1 0 3360 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_26
timestamp 1694700623
transform 1 0 4256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_28
timestamp 1694700623
transform 1 0 4480 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_31
timestamp 1694700623
transform 1 0 4816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_37
timestamp 1694700623
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_45
timestamp 1694700623
transform 1 0 6384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_49
timestamp 1694700623
transform 1 0 6832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_51
timestamp 1694700623
transform 1 0 7056 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_69
timestamp 1694700623
transform 1 0 9072 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_73
timestamp 1694700623
transform 1 0 9520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_75
timestamp 1694700623
transform 1 0 9744 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_82
timestamp 1694700623
transform 1 0 10528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_86
timestamp 1694700623
transform 1 0 10976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_88
timestamp 1694700623
transform 1 0 11200 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_95
timestamp 1694700623
transform 1 0 11984 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1694700623
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_137
timestamp 1694700623
transform 1 0 16688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_145
timestamp 1694700623
transform 1 0 17584 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_149
timestamp 1694700623
transform 1 0 18032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_151
timestamp 1694700623
transform 1 0 18256 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_164
timestamp 1694700623
transform 1 0 19712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_166
timestamp 1694700623
transform 1 0 19936 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_177
timestamp 1694700623
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_181
timestamp 1694700623
transform 1 0 21616 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_185
timestamp 1694700623
transform 1 0 22064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_210
timestamp 1694700623
transform 1 0 24864 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1694700623
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1694700623
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_247
timestamp 1694700623
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_255
timestamp 1694700623
transform 1 0 29904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_259
timestamp 1694700623
transform 1 0 30352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_292
timestamp 1694700623
transform 1 0 34048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_300
timestamp 1694700623
transform 1 0 34944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_302
timestamp 1694700623
transform 1 0 35168 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1694700623
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_317
timestamp 1694700623
transform 1 0 36848 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_333
timestamp 1694700623
transform 1 0 38640 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_342
timestamp 1694700623
transform 1 0 39648 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_358
timestamp 1694700623
transform 1 0 41440 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_366
timestamp 1694700623
transform 1 0 42336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_370
timestamp 1694700623
transform 1 0 42784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_380
timestamp 1694700623
transform 1 0 43904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1694700623
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_387
timestamp 1694700623
transform 1 0 44688 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_447
timestamp 1694700623
transform 1 0 51408 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1694700623
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_457
timestamp 1694700623
transform 1 0 52528 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_465
timestamp 1694700623
transform 1 0 53424 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_469
timestamp 1694700623
transform 1 0 53872 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_476
timestamp 1694700623
transform 1 0 54656 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_484
timestamp 1694700623
transform 1 0 55552 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_493
timestamp 1694700623
transform 1 0 56560 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_2
timestamp 1694700623
transform 1 0 1568 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_18
timestamp 1694700623
transform 1 0 3360 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_26
timestamp 1694700623
transform 1 0 4256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_30
timestamp 1694700623
transform 1 0 4704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_32
timestamp 1694700623
transform 1 0 4928 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_72
timestamp 1694700623
transform 1 0 9408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_76
timestamp 1694700623
transform 1 0 9856 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_107
timestamp 1694700623
transform 1 0 13328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_111
timestamp 1694700623
transform 1 0 13776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_115
timestamp 1694700623
transform 1 0 14224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_117
timestamp 1694700623
transform 1 0 14448 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_123
timestamp 1694700623
transform 1 0 15120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1694700623
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_206
timestamp 1694700623
transform 1 0 24416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1694700623
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_216
timestamp 1694700623
transform 1 0 25536 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_248
timestamp 1694700623
transform 1 0 29120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_264
timestamp 1694700623
transform 1 0 30912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_282
timestamp 1694700623
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_284
timestamp 1694700623
transform 1 0 33152 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_297
timestamp 1694700623
transform 1 0 34608 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_318
timestamp 1694700623
transform 1 0 36960 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1694700623
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_356
timestamp 1694700623
transform 1 0 41216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_364
timestamp 1694700623
transform 1 0 42112 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_395
timestamp 1694700623
transform 1 0 45584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_399
timestamp 1694700623
transform 1 0 46032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_410
timestamp 1694700623
transform 1 0 47264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_414
timestamp 1694700623
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1694700623
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_422
timestamp 1694700623
transform 1 0 48608 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_438
timestamp 1694700623
transform 1 0 50400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_477
timestamp 1694700623
transform 1 0 54768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_481
timestamp 1694700623
transform 1 0 55216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1694700623
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_492
timestamp 1694700623
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_496
timestamp 1694700623
transform 1 0 56896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_498
timestamp 1694700623
transform 1 0 57120 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_2
timestamp 1694700623
transform 1 0 1568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_10
timestamp 1694700623
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_12
timestamp 1694700623
transform 1 0 2688 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_30
timestamp 1694700623
transform 1 0 4704 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1694700623
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_37
timestamp 1694700623
transform 1 0 5488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_45
timestamp 1694700623
transform 1 0 6384 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_49
timestamp 1694700623
transform 1 0 6832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_71
timestamp 1694700623
transform 1 0 9296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_85
timestamp 1694700623
transform 1 0 10864 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1694700623
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_107
timestamp 1694700623
transform 1 0 13328 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_139
timestamp 1694700623
transform 1 0 16912 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_143
timestamp 1694700623
transform 1 0 17360 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1694700623
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_177
timestamp 1694700623
transform 1 0 21168 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_185
timestamp 1694700623
transform 1 0 22064 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_211
timestamp 1694700623
transform 1 0 24976 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1694700623
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_261
timestamp 1694700623
transform 1 0 30576 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_277
timestamp 1694700623
transform 1 0 32368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_281
timestamp 1694700623
transform 1 0 32816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_285
timestamp 1694700623
transform 1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_287
timestamp 1694700623
transform 1 0 33488 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_329
timestamp 1694700623
transform 1 0 38192 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_337
timestamp 1694700623
transform 1 0 39088 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_339
timestamp 1694700623
transform 1 0 39312 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_350
timestamp 1694700623
transform 1 0 40544 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_362
timestamp 1694700623
transform 1 0 41888 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_378
timestamp 1694700623
transform 1 0 43680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_382
timestamp 1694700623
transform 1 0 44128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1694700623
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_387
timestamp 1694700623
transform 1 0 44688 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_419
timestamp 1694700623
transform 1 0 48272 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_435
timestamp 1694700623
transform 1 0 50064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_443
timestamp 1694700623
transform 1 0 50960 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1694700623
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_463
timestamp 1694700623
transform 1 0 53200 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_467
timestamp 1694700623
transform 1 0 53648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_39
timestamp 1694700623
transform 1 0 5712 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_55
timestamp 1694700623
transform 1 0 7504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_63
timestamp 1694700623
transform 1 0 8400 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_67
timestamp 1694700623
transform 1 0 8848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_69
timestamp 1694700623
transform 1 0 9072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_72
timestamp 1694700623
transform 1 0 9408 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_80
timestamp 1694700623
transform 1 0 10304 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_84
timestamp 1694700623
transform 1 0 10752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_91
timestamp 1694700623
transform 1 0 11536 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_107
timestamp 1694700623
transform 1 0 13328 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_111
timestamp 1694700623
transform 1 0 13776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_133
timestamp 1694700623
transform 1 0 16240 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_137
timestamp 1694700623
transform 1 0 16688 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1694700623
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_142
timestamp 1694700623
transform 1 0 17248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_150
timestamp 1694700623
transform 1 0 18144 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_153
timestamp 1694700623
transform 1 0 18480 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_185
timestamp 1694700623
transform 1 0 22064 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_201
timestamp 1694700623
transform 1 0 23856 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1694700623
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_212
timestamp 1694700623
transform 1 0 25088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_220
timestamp 1694700623
transform 1 0 25984 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_224
timestamp 1694700623
transform 1 0 26432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_253
timestamp 1694700623
transform 1 0 29680 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_257
timestamp 1694700623
transform 1 0 30128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_271
timestamp 1694700623
transform 1 0 31696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_275
timestamp 1694700623
transform 1 0 32144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1694700623
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1694700623
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_286
timestamp 1694700623
transform 1 0 33376 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_318
timestamp 1694700623
transform 1 0 36960 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_334
timestamp 1694700623
transform 1 0 38752 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_338
timestamp 1694700623
transform 1 0 39200 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_347
timestamp 1694700623
transform 1 0 40208 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1694700623
transform 1 0 40432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1694700623
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_369
timestamp 1694700623
transform 1 0 42672 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_385
timestamp 1694700623
transform 1 0 44464 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_393
timestamp 1694700623
transform 1 0 45360 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1694700623
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1694700623
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_422
timestamp 1694700623
transform 1 0 48608 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_438
timestamp 1694700623
transform 1 0 50400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_440
timestamp 1694700623
transform 1 0 50624 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_453
timestamp 1694700623
transform 1 0 52080 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_469
timestamp 1694700623
transform 1 0 53872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_473
timestamp 1694700623
transform 1 0 54320 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_482
timestamp 1694700623
transform 1 0 55328 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_500
timestamp 1694700623
transform 1 0 57344 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1694700623
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_2
timestamp 1694700623
transform 1 0 1568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_10
timestamp 1694700623
transform 1 0 2464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_33
timestamp 1694700623
transform 1 0 5040 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1694700623
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_69
timestamp 1694700623
transform 1 0 9072 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_90
timestamp 1694700623
transform 1 0 11424 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_92
timestamp 1694700623
transform 1 0 11648 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_95
timestamp 1694700623
transform 1 0 11984 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_99
timestamp 1694700623
transform 1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_103
timestamp 1694700623
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_107
timestamp 1694700623
transform 1 0 13328 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_111
timestamp 1694700623
transform 1 0 13776 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_115
timestamp 1694700623
transform 1 0 14224 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_120
timestamp 1694700623
transform 1 0 14784 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_154
timestamp 1694700623
transform 1 0 18592 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_170
timestamp 1694700623
transform 1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1694700623
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_177
timestamp 1694700623
transform 1 0 21168 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_193
timestamp 1694700623
transform 1 0 22960 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_203
timestamp 1694700623
transform 1 0 24080 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_219
timestamp 1694700623
transform 1 0 25872 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_227
timestamp 1694700623
transform 1 0 26768 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_231
timestamp 1694700623
transform 1 0 27216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_233
timestamp 1694700623
transform 1 0 27440 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_242
timestamp 1694700623
transform 1 0 28448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1694700623
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_247
timestamp 1694700623
transform 1 0 29008 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_272
timestamp 1694700623
transform 1 0 31808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_292
timestamp 1694700623
transform 1 0 34048 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_294
timestamp 1694700623
transform 1 0 34272 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_305
timestamp 1694700623
transform 1 0 35504 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_313
timestamp 1694700623
transform 1 0 36400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_317
timestamp 1694700623
transform 1 0 36848 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_321
timestamp 1694700623
transform 1 0 37296 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_375
timestamp 1694700623
transform 1 0 43344 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_416
timestamp 1694700623
transform 1 0 47936 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_424
timestamp 1694700623
transform 1 0 48832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_432
timestamp 1694700623
transform 1 0 49728 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_439
timestamp 1694700623
transform 1 0 50512 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_466
timestamp 1694700623
transform 1 0 53536 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_474
timestamp 1694700623
transform 1 0 54432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_505
timestamp 1694700623
transform 1 0 57904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1694700623
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1694700623
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_26
timestamp 1694700623
transform 1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_30
timestamp 1694700623
transform 1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_32
timestamp 1694700623
transform 1 0 4928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_35
timestamp 1694700623
transform 1 0 5264 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_51
timestamp 1694700623
transform 1 0 7056 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_59
timestamp 1694700623
transform 1 0 7952 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_68
timestamp 1694700623
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_72
timestamp 1694700623
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_74
timestamp 1694700623
transform 1 0 9632 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_77
timestamp 1694700623
transform 1 0 9968 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_86
timestamp 1694700623
transform 1 0 10976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_93
timestamp 1694700623
transform 1 0 11760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_116
timestamp 1694700623
transform 1 0 14336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_133
timestamp 1694700623
transform 1 0 16240 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_137
timestamp 1694700623
transform 1 0 16688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_139
timestamp 1694700623
transform 1 0 16912 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_142
timestamp 1694700623
transform 1 0 17248 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_152
timestamp 1694700623
transform 1 0 18368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_177
timestamp 1694700623
transform 1 0 21168 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_185
timestamp 1694700623
transform 1 0 22064 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_209
timestamp 1694700623
transform 1 0 24752 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_212
timestamp 1694700623
transform 1 0 25088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_216
timestamp 1694700623
transform 1 0 25536 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_232
timestamp 1694700623
transform 1 0 27328 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_240
timestamp 1694700623
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_244
timestamp 1694700623
transform 1 0 28672 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_260
timestamp 1694700623
transform 1 0 30464 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_264
timestamp 1694700623
transform 1 0 30912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_266
timestamp 1694700623
transform 1 0 31136 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_269
timestamp 1694700623
transform 1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_282
timestamp 1694700623
transform 1 0 32928 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_344
timestamp 1694700623
transform 1 0 39872 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_348
timestamp 1694700623
transform 1 0 40320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_352
timestamp 1694700623
transform 1 0 40768 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_384
timestamp 1694700623
transform 1 0 44352 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_392
timestamp 1694700623
transform 1 0 45248 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_397
timestamp 1694700623
transform 1 0 45808 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_419
timestamp 1694700623
transform 1 0 48272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_426
timestamp 1694700623
transform 1 0 49056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_430
timestamp 1694700623
transform 1 0 49504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_432
timestamp 1694700623
transform 1 0 49728 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_439
timestamp 1694700623
transform 1 0 50512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_470
timestamp 1694700623
transform 1 0 53984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_474
timestamp 1694700623
transform 1 0 54432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_488
timestamp 1694700623
transform 1 0 56000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_492
timestamp 1694700623
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1694700623
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_2
timestamp 1694700623
transform 1 0 1568 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_18
timestamp 1694700623
transform 1 0 3360 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_22
timestamp 1694700623
transform 1 0 3808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_24
timestamp 1694700623
transform 1 0 4032 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_33
timestamp 1694700623
transform 1 0 5040 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_45
timestamp 1694700623
transform 1 0 6384 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_87
timestamp 1694700623
transform 1 0 11088 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_91
timestamp 1694700623
transform 1 0 11536 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_93
timestamp 1694700623
transform 1 0 11760 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_102
timestamp 1694700623
transform 1 0 12768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1694700623
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_125
timestamp 1694700623
transform 1 0 15344 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_129
timestamp 1694700623
transform 1 0 15792 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_131
timestamp 1694700623
transform 1 0 16016 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_171
timestamp 1694700623
transform 1 0 20496 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_233
timestamp 1694700623
transform 1 0 27440 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_237
timestamp 1694700623
transform 1 0 27888 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_247
timestamp 1694700623
transform 1 0 29008 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_249
timestamp 1694700623
transform 1 0 29232 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_265
timestamp 1694700623
transform 1 0 31024 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_298
timestamp 1694700623
transform 1 0 34720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_302
timestamp 1694700623
transform 1 0 35168 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_306
timestamp 1694700623
transform 1 0 35616 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_329
timestamp 1694700623
transform 1 0 38192 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_361
timestamp 1694700623
transform 1 0 41776 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_379
timestamp 1694700623
transform 1 0 43792 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_383
timestamp 1694700623
transform 1 0 44240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_387
timestamp 1694700623
transform 1 0 44688 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_403
timestamp 1694700623
transform 1 0 46480 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_436
timestamp 1694700623
transform 1 0 50176 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_440
timestamp 1694700623
transform 1 0 50624 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_448
timestamp 1694700623
transform 1 0 51520 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_452
timestamp 1694700623
transform 1 0 51968 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_454
timestamp 1694700623
transform 1 0 52192 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_457
timestamp 1694700623
transform 1 0 52528 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_473
timestamp 1694700623
transform 1 0 54320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_477
timestamp 1694700623
transform 1 0 54768 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_479
timestamp 1694700623
transform 1 0 54992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_486
timestamp 1694700623
transform 1 0 55776 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_502
timestamp 1694700623
transform 1 0 57568 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_506
timestamp 1694700623
transform 1 0 58016 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_508
timestamp 1694700623
transform 1 0 58240 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_51
timestamp 1694700623
transform 1 0 7056 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_55
timestamp 1694700623
transform 1 0 7504 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_57
timestamp 1694700623
transform 1 0 7728 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1694700623
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_85
timestamp 1694700623
transform 1 0 10864 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_101
timestamp 1694700623
transform 1 0 12656 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_105
timestamp 1694700623
transform 1 0 13104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_114
timestamp 1694700623
transform 1 0 14112 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_130
timestamp 1694700623
transform 1 0 15904 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_138
timestamp 1694700623
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_142
timestamp 1694700623
transform 1 0 17248 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_158
timestamp 1694700623
transform 1 0 19040 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_160
timestamp 1694700623
transform 1 0 19264 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_174
timestamp 1694700623
transform 1 0 20832 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_182
timestamp 1694700623
transform 1 0 21728 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_186
timestamp 1694700623
transform 1 0 22176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_188
timestamp 1694700623
transform 1 0 22400 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_212
timestamp 1694700623
transform 1 0 25088 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_242
timestamp 1694700623
transform 1 0 28448 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_246
timestamp 1694700623
transform 1 0 28896 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_248
timestamp 1694700623
transform 1 0 29120 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_272
timestamp 1694700623
transform 1 0 31808 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_279
timestamp 1694700623
transform 1 0 32592 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_282
timestamp 1694700623
transform 1 0 32928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_286
timestamp 1694700623
transform 1 0 33376 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_302
timestamp 1694700623
transform 1 0 35168 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_306
timestamp 1694700623
transform 1 0 35616 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_308
timestamp 1694700623
transform 1 0 35840 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_338
timestamp 1694700623
transform 1 0 39200 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1694700623
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_352
timestamp 1694700623
transform 1 0 40768 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_360
timestamp 1694700623
transform 1 0 41664 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_393
timestamp 1694700623
transform 1 0 45360 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_409
timestamp 1694700623
transform 1 0 47152 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_417
timestamp 1694700623
transform 1 0 48048 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_419
timestamp 1694700623
transform 1 0 48272 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_422
timestamp 1694700623
transform 1 0 48608 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_438
timestamp 1694700623
transform 1 0 50400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_442
timestamp 1694700623
transform 1 0 50848 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_454
timestamp 1694700623
transform 1 0 52192 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_456
timestamp 1694700623
transform 1 0 52416 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_459
timestamp 1694700623
transform 1 0 52752 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_475
timestamp 1694700623
transform 1 0 54544 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_483
timestamp 1694700623
transform 1 0 55440 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_487
timestamp 1694700623
transform 1 0 55888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_489
timestamp 1694700623
transform 1 0 56112 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_492
timestamp 1694700623
transform 1 0 56448 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_508
timestamp 1694700623
transform 1 0 58240 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_10
timestamp 1694700623
transform 1 0 2464 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_18
timestamp 1694700623
transform 1 0 3360 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_20
timestamp 1694700623
transform 1 0 3584 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_29
timestamp 1694700623
transform 1 0 4592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_33
timestamp 1694700623
transform 1 0 5040 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_42
timestamp 1694700623
transform 1 0 6048 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_74
timestamp 1694700623
transform 1 0 9632 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_76
timestamp 1694700623
transform 1 0 9856 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_100
timestamp 1694700623
transform 1 0 12544 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1694700623
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_113
timestamp 1694700623
transform 1 0 14000 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_119
timestamp 1694700623
transform 1 0 14672 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_123
timestamp 1694700623
transform 1 0 15120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_127
timestamp 1694700623
transform 1 0 15568 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_139
timestamp 1694700623
transform 1 0 16912 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1694700623
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_177
timestamp 1694700623
transform 1 0 21168 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_209
timestamp 1694700623
transform 1 0 24752 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_217
timestamp 1694700623
transform 1 0 25648 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_221
timestamp 1694700623
transform 1 0 26096 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_223
timestamp 1694700623
transform 1 0 26320 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1694700623
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_247
timestamp 1694700623
transform 1 0 29008 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_251
timestamp 1694700623
transform 1 0 29456 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_264
timestamp 1694700623
transform 1 0 30912 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_296
timestamp 1694700623
transform 1 0 34496 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_304
timestamp 1694700623
transform 1 0 35392 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1694700623
transform 1 0 36512 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1694700623
transform 1 0 36848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1694700623
transform 1 0 37744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_329
timestamp 1694700623
transform 1 0 38192 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_359
timestamp 1694700623
transform 1 0 41552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_363
timestamp 1694700623
transform 1 0 42000 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_376
timestamp 1694700623
transform 1 0 43456 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_384
timestamp 1694700623
transform 1 0 44352 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_416
timestamp 1694700623
transform 1 0 47936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_420
timestamp 1694700623
transform 1 0 48384 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_436
timestamp 1694700623
transform 1 0 50176 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_444
timestamp 1694700623
transform 1 0 51072 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_448
timestamp 1694700623
transform 1 0 51520 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_450
timestamp 1694700623
transform 1 0 51744 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_457
timestamp 1694700623
transform 1 0 52528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_485
timestamp 1694700623
transform 1 0 55664 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_501
timestamp 1694700623
transform 1 0 57456 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_505
timestamp 1694700623
transform 1 0 57904 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_2
timestamp 1694700623
transform 1 0 1568 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_6
timestamp 1694700623
transform 1 0 2016 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_38
timestamp 1694700623
transform 1 0 5600 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_46
timestamp 1694700623
transform 1 0 6496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_50
timestamp 1694700623
transform 1 0 6944 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_52
timestamp 1694700623
transform 1 0 7168 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_59
timestamp 1694700623
transform 1 0 7952 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_63
timestamp 1694700623
transform 1 0 8400 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_67
timestamp 1694700623
transform 1 0 8848 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1694700623
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_72
timestamp 1694700623
transform 1 0 9408 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_88
timestamp 1694700623
transform 1 0 11200 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_125
timestamp 1694700623
transform 1 0 15344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_139
timestamp 1694700623
transform 1 0 16912 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_151
timestamp 1694700623
transform 1 0 18256 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_183
timestamp 1694700623
transform 1 0 21840 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_199
timestamp 1694700623
transform 1 0 23632 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_207
timestamp 1694700623
transform 1 0 24528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1694700623
transform 1 0 24752 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_212
timestamp 1694700623
transform 1 0 25088 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_234
timestamp 1694700623
transform 1 0 27552 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_238
timestamp 1694700623
transform 1 0 28000 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_254
timestamp 1694700623
transform 1 0 29792 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_262
timestamp 1694700623
transform 1 0 30688 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_266
timestamp 1694700623
transform 1 0 31136 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_274
timestamp 1694700623
transform 1 0 32032 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_278
timestamp 1694700623
transform 1 0 32480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_282
timestamp 1694700623
transform 1 0 32928 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_298
timestamp 1694700623
transform 1 0 34720 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_302
timestamp 1694700623
transform 1 0 35168 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_323
timestamp 1694700623
transform 1 0 37520 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_331
timestamp 1694700623
transform 1 0 38416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_335
timestamp 1694700623
transform 1 0 38864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_337
timestamp 1694700623
transform 1 0 39088 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_360
timestamp 1694700623
transform 1 0 41664 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_375
timestamp 1694700623
transform 1 0 43344 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_383
timestamp 1694700623
transform 1 0 44240 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_387
timestamp 1694700623
transform 1 0 44688 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_394
timestamp 1694700623
transform 1 0 45472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_398
timestamp 1694700623
transform 1 0 45920 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_414
timestamp 1694700623
transform 1 0 47712 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_436
timestamp 1694700623
transform 1 0 50176 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_440
timestamp 1694700623
transform 1 0 50624 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_444
timestamp 1694700623
transform 1 0 51072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_474
timestamp 1694700623
transform 1 0 54432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_478
timestamp 1694700623
transform 1 0 54880 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_486
timestamp 1694700623
transform 1 0 55776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_498
timestamp 1694700623
transform 1 0 57120 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_500
timestamp 1694700623
transform 1 0 57344 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1694700623
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1694700623
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_37
timestamp 1694700623
transform 1 0 5488 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_39
timestamp 1694700623
transform 1 0 5712 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_42
timestamp 1694700623
transform 1 0 6048 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_59
timestamp 1694700623
transform 1 0 7952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_90
timestamp 1694700623
transform 1 0 11424 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_130
timestamp 1694700623
transform 1 0 15904 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_149
timestamp 1694700623
transform 1 0 18032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_177
timestamp 1694700623
transform 1 0 21168 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_181
timestamp 1694700623
transform 1 0 21616 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_183
timestamp 1694700623
transform 1 0 21840 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_186
timestamp 1694700623
transform 1 0 22176 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_188
timestamp 1694700623
transform 1 0 22400 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_231
timestamp 1694700623
transform 1 0 27216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_243
timestamp 1694700623
transform 1 0 28560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_252
timestamp 1694700623
transform 1 0 29568 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_256
timestamp 1694700623
transform 1 0 30016 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_286
timestamp 1694700623
transform 1 0 33376 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_290
timestamp 1694700623
transform 1 0 33824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_300
timestamp 1694700623
transform 1 0 34944 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_308
timestamp 1694700623
transform 1 0 35840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_312
timestamp 1694700623
transform 1 0 36288 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_314
timestamp 1694700623
transform 1 0 36512 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_317
timestamp 1694700623
transform 1 0 36848 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_335
timestamp 1694700623
transform 1 0 38864 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_343
timestamp 1694700623
transform 1 0 39760 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_387
timestamp 1694700623
transform 1 0 44688 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_403
timestamp 1694700623
transform 1 0 46480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_405
timestamp 1694700623
transform 1 0 46704 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_457
timestamp 1694700623
transform 1 0 52528 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_473
timestamp 1694700623
transform 1 0 54320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_477
timestamp 1694700623
transform 1 0 54768 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_2
timestamp 1694700623
transform 1 0 1568 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_10
timestamp 1694700623
transform 1 0 2464 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_63
timestamp 1694700623
transform 1 0 8400 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_67
timestamp 1694700623
transform 1 0 8848 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_69
timestamp 1694700623
transform 1 0 9072 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_72
timestamp 1694700623
transform 1 0 9408 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_80
timestamp 1694700623
transform 1 0 10304 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_82
timestamp 1694700623
transform 1 0 10528 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_109
timestamp 1694700623
transform 1 0 13552 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_113
timestamp 1694700623
transform 1 0 14000 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_117
timestamp 1694700623
transform 1 0 14448 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_133
timestamp 1694700623
transform 1 0 16240 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_137
timestamp 1694700623
transform 1 0 16688 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_139
timestamp 1694700623
transform 1 0 16912 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_152
timestamp 1694700623
transform 1 0 18368 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_154
timestamp 1694700623
transform 1 0 18592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_223
timestamp 1694700623
transform 1 0 26320 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_227
timestamp 1694700623
transform 1 0 26768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_258
timestamp 1694700623
transform 1 0 30240 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_262
timestamp 1694700623
transform 1 0 30688 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_278
timestamp 1694700623
transform 1 0 32480 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_318
timestamp 1694700623
transform 1 0 36960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_348
timestamp 1694700623
transform 1 0 40320 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_352
timestamp 1694700623
transform 1 0 40768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_360
timestamp 1694700623
transform 1 0 41664 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_364
timestamp 1694700623
transform 1 0 42112 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_372
timestamp 1694700623
transform 1 0 43008 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_404
timestamp 1694700623
transform 1 0 46592 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_422
timestamp 1694700623
transform 1 0 48608 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_437
timestamp 1694700623
transform 1 0 50288 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_441
timestamp 1694700623
transform 1 0 50736 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_448
timestamp 1694700623
transform 1 0 51520 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_456
timestamp 1694700623
transform 1 0 52416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_466
timestamp 1694700623
transform 1 0 53536 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_508
timestamp 1694700623
transform 1 0 58240 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1694700623
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1694700623
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_37
timestamp 1694700623
transform 1 0 5488 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_52
timestamp 1694700623
transform 1 0 7168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_54
timestamp 1694700623
transform 1 0 7392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_57
timestamp 1694700623
transform 1 0 7728 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_89
timestamp 1694700623
transform 1 0 11312 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_99
timestamp 1694700623
transform 1 0 12432 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_103
timestamp 1694700623
transform 1 0 12880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_107
timestamp 1694700623
transform 1 0 13328 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_139
timestamp 1694700623
transform 1 0 16912 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_155
timestamp 1694700623
transform 1 0 18704 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_163
timestamp 1694700623
transform 1 0 19600 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_171
timestamp 1694700623
transform 1 0 20496 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_177
timestamp 1694700623
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_179
timestamp 1694700623
transform 1 0 21392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_213
timestamp 1694700623
transform 1 0 25200 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_217
timestamp 1694700623
transform 1 0 25648 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_221
timestamp 1694700623
transform 1 0 26096 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_237
timestamp 1694700623
transform 1 0 27888 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_247
timestamp 1694700623
transform 1 0 29008 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_263
timestamp 1694700623
transform 1 0 30800 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_271
timestamp 1694700623
transform 1 0 31696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_275
timestamp 1694700623
transform 1 0 32144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_282
timestamp 1694700623
transform 1 0 32928 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_290
timestamp 1694700623
transform 1 0 33824 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_294
timestamp 1694700623
transform 1 0 34272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_307
timestamp 1694700623
transform 1 0 35728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_325
timestamp 1694700623
transform 1 0 37744 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_327
timestamp 1694700623
transform 1 0 37968 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_334
timestamp 1694700623
transform 1 0 38752 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_366
timestamp 1694700623
transform 1 0 42336 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_380
timestamp 1694700623
transform 1 0 43904 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_384
timestamp 1694700623
transform 1 0 44352 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_387
timestamp 1694700623
transform 1 0 44688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_391
timestamp 1694700623
transform 1 0 45136 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_423
timestamp 1694700623
transform 1 0 48720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_429
timestamp 1694700623
transform 1 0 49392 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_445
timestamp 1694700623
transform 1 0 51184 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_453
timestamp 1694700623
transform 1 0 52080 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_507
timestamp 1694700623
transform 1 0 58128 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_2
timestamp 1694700623
transform 1 0 1568 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_34
timestamp 1694700623
transform 1 0 5152 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_42
timestamp 1694700623
transform 1 0 6048 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_46
timestamp 1694700623
transform 1 0 6496 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_55
timestamp 1694700623
transform 1 0 7504 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_67
timestamp 1694700623
transform 1 0 8848 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_69
timestamp 1694700623
transform 1 0 9072 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_87
timestamp 1694700623
transform 1 0 11088 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_95
timestamp 1694700623
transform 1 0 11984 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_99
timestamp 1694700623
transform 1 0 12432 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_101
timestamp 1694700623
transform 1 0 12656 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_115
timestamp 1694700623
transform 1 0 14224 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_125
timestamp 1694700623
transform 1 0 15344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_129
timestamp 1694700623
transform 1 0 15792 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_138
timestamp 1694700623
transform 1 0 16800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_142
timestamp 1694700623
transform 1 0 17248 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_150
timestamp 1694700623
transform 1 0 18144 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_154
timestamp 1694700623
transform 1 0 18592 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_172
timestamp 1694700623
transform 1 0 20608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_176
timestamp 1694700623
transform 1 0 21056 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_208
timestamp 1694700623
transform 1 0 24640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_212
timestamp 1694700623
transform 1 0 25088 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_228
timestamp 1694700623
transform 1 0 26880 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_232
timestamp 1694700623
transform 1 0 27328 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_234
timestamp 1694700623
transform 1 0 27552 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_237
timestamp 1694700623
transform 1 0 27888 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_253
timestamp 1694700623
transform 1 0 29680 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_261
timestamp 1694700623
transform 1 0 30576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_265
timestamp 1694700623
transform 1 0 31024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_269
timestamp 1694700623
transform 1 0 31472 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_277
timestamp 1694700623
transform 1 0 32368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_279
timestamp 1694700623
transform 1 0 32592 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_282
timestamp 1694700623
transform 1 0 32928 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_314
timestamp 1694700623
transform 1 0 36512 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_328
timestamp 1694700623
transform 1 0 38080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_342
timestamp 1694700623
transform 1 0 39648 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_384
timestamp 1694700623
transform 1 0 44352 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_412
timestamp 1694700623
transform 1 0 47488 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_451
timestamp 1694700623
transform 1 0 51856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_463
timestamp 1694700623
transform 1 0 53200 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_497
timestamp 1694700623
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_501
timestamp 1694700623
transform 1 0 57456 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_2
timestamp 1694700623
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1694700623
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_37
timestamp 1694700623
transform 1 0 5488 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_53
timestamp 1694700623
transform 1 0 7280 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_67
timestamp 1694700623
transform 1 0 8848 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_107
timestamp 1694700623
transform 1 0 13328 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_115
timestamp 1694700623
transform 1 0 14224 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_150
timestamp 1694700623
transform 1 0 18144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_154
timestamp 1694700623
transform 1 0 18592 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_168
timestamp 1694700623
transform 1 0 20160 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_172
timestamp 1694700623
transform 1 0 20608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_174
timestamp 1694700623
transform 1 0 20832 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_203
timestamp 1694700623
transform 1 0 24080 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_219
timestamp 1694700623
transform 1 0 25872 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_241
timestamp 1694700623
transform 1 0 28336 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_247
timestamp 1694700623
transform 1 0 29008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_249
timestamp 1694700623
transform 1 0 29232 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_262
timestamp 1694700623
transform 1 0 30688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_264
timestamp 1694700623
transform 1 0 30912 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_270
timestamp 1694700623
transform 1 0 31584 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_272
timestamp 1694700623
transform 1 0 31808 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_280
timestamp 1694700623
transform 1 0 32704 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_284
timestamp 1694700623
transform 1 0 33152 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_300
timestamp 1694700623
transform 1 0 34944 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_308
timestamp 1694700623
transform 1 0 35840 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_312
timestamp 1694700623
transform 1 0 36288 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_314
timestamp 1694700623
transform 1 0 36512 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_317
timestamp 1694700623
transform 1 0 36848 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_333
timestamp 1694700623
transform 1 0 38640 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_341
timestamp 1694700623
transform 1 0 39536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_345
timestamp 1694700623
transform 1 0 39984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_378
timestamp 1694700623
transform 1 0 43680 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_416
timestamp 1694700623
transform 1 0 47936 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_432
timestamp 1694700623
transform 1 0 49728 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_436
timestamp 1694700623
transform 1 0 50176 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_452
timestamp 1694700623
transform 1 0 51968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_454
timestamp 1694700623
transform 1 0 52192 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_457
timestamp 1694700623
transform 1 0 52528 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_459
timestamp 1694700623
transform 1 0 52752 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_476
timestamp 1694700623
transform 1 0 54656 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_2
timestamp 1694700623
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_68
timestamp 1694700623
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_72
timestamp 1694700623
transform 1 0 9408 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_80
timestamp 1694700623
transform 1 0 10304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_84
timestamp 1694700623
transform 1 0 10752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_117
timestamp 1694700623
transform 1 0 14448 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_133
timestamp 1694700623
transform 1 0 16240 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_137
timestamp 1694700623
transform 1 0 16688 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_139
timestamp 1694700623
transform 1 0 16912 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_150
timestamp 1694700623
transform 1 0 18144 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_195
timestamp 1694700623
transform 1 0 23184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_199
timestamp 1694700623
transform 1 0 23632 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_207
timestamp 1694700623
transform 1 0 24528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_209
timestamp 1694700623
transform 1 0 24752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_212
timestamp 1694700623
transform 1 0 25088 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_266
timestamp 1694700623
transform 1 0 31136 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_306
timestamp 1694700623
transform 1 0 35616 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_338
timestamp 1694700623
transform 1 0 39200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_342
timestamp 1694700623
transform 1 0 39648 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_352
timestamp 1694700623
transform 1 0 40768 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_356
timestamp 1694700623
transform 1 0 41216 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_358
timestamp 1694700623
transform 1 0 41440 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_361
timestamp 1694700623
transform 1 0 41776 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_365
timestamp 1694700623
transform 1 0 42224 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_369
timestamp 1694700623
transform 1 0 42672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_377
timestamp 1694700623
transform 1 0 43568 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_381
timestamp 1694700623
transform 1 0 44016 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_410
timestamp 1694700623
transform 1 0 47264 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_418
timestamp 1694700623
transform 1 0 48160 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_422
timestamp 1694700623
transform 1 0 48608 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_426
timestamp 1694700623
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_442
timestamp 1694700623
transform 1 0 50848 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_444
timestamp 1694700623
transform 1 0 51072 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_479
timestamp 1694700623
transform 1 0 54992 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_489
timestamp 1694700623
transform 1 0 56112 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_492
timestamp 1694700623
transform 1 0 56448 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_508
timestamp 1694700623
transform 1 0 58240 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1694700623
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1694700623
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_136
timestamp 1694700623
transform 1 0 16576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_140
timestamp 1694700623
transform 1 0 17024 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_144
timestamp 1694700623
transform 1 0 17472 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_177
timestamp 1694700623
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_181
timestamp 1694700623
transform 1 0 21616 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_189
timestamp 1694700623
transform 1 0 22512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_193
timestamp 1694700623
transform 1 0 22960 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_238
timestamp 1694700623
transform 1 0 28000 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_242
timestamp 1694700623
transform 1 0 28448 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_255
timestamp 1694700623
transform 1 0 29904 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_267
timestamp 1694700623
transform 1 0 31248 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_271
timestamp 1694700623
transform 1 0 31696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_275
timestamp 1694700623
transform 1 0 32144 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_317
timestamp 1694700623
transform 1 0 36848 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_321
timestamp 1694700623
transform 1 0 37296 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_329
timestamp 1694700623
transform 1 0 38192 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_387
timestamp 1694700623
transform 1 0 44688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_391
timestamp 1694700623
transform 1 0 45136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_395
timestamp 1694700623
transform 1 0 45584 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_403
timestamp 1694700623
transform 1 0 46480 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_407
timestamp 1694700623
transform 1 0 46928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_439
timestamp 1694700623
transform 1 0 50512 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_447
timestamp 1694700623
transform 1 0 51408 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_452
timestamp 1694700623
transform 1 0 51968 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_454
timestamp 1694700623
transform 1 0 52192 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_457
timestamp 1694700623
transform 1 0 52528 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_461
timestamp 1694700623
transform 1 0 52976 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_477
timestamp 1694700623
transform 1 0 54768 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1694700623
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_66
timestamp 1694700623
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_72
timestamp 1694700623
transform 1 0 9408 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_88
timestamp 1694700623
transform 1 0 11200 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_96
timestamp 1694700623
transform 1 0 12096 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_98
timestamp 1694700623
transform 1 0 12320 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_101
timestamp 1694700623
transform 1 0 12656 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_107
timestamp 1694700623
transform 1 0 13328 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_139
timestamp 1694700623
transform 1 0 16912 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_171
timestamp 1694700623
transform 1 0 20496 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_175
timestamp 1694700623
transform 1 0 20944 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_179
timestamp 1694700623
transform 1 0 21392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_212
timestamp 1694700623
transform 1 0 25088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_216
timestamp 1694700623
transform 1 0 25536 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_224
timestamp 1694700623
transform 1 0 26432 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_228
timestamp 1694700623
transform 1 0 26880 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_255
timestamp 1694700623
transform 1 0 29904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_259
timestamp 1694700623
transform 1 0 30352 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_275
timestamp 1694700623
transform 1 0 32144 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_279
timestamp 1694700623
transform 1 0 32592 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_282
timestamp 1694700623
transform 1 0 32928 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_290
timestamp 1694700623
transform 1 0 33824 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_294
timestamp 1694700623
transform 1 0 34272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_296
timestamp 1694700623
transform 1 0 34496 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_303
timestamp 1694700623
transform 1 0 35280 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_307
timestamp 1694700623
transform 1 0 35728 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_311
timestamp 1694700623
transform 1 0 36176 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_313
timestamp 1694700623
transform 1 0 36400 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_343
timestamp 1694700623
transform 1 0 39760 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_347
timestamp 1694700623
transform 1 0 40208 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_349
timestamp 1694700623
transform 1 0 40432 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_352
timestamp 1694700623
transform 1 0 40768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_356
timestamp 1694700623
transform 1 0 41216 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1694700623
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_480
timestamp 1694700623
transform 1 0 55104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_484
timestamp 1694700623
transform 1 0 55552 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_488
timestamp 1694700623
transform 1 0 56000 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_492
timestamp 1694700623
transform 1 0 56448 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_500
timestamp 1694700623
transform 1 0 57344 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_2
timestamp 1694700623
transform 1 0 1568 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_10
timestamp 1694700623
transform 1 0 2464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_12
timestamp 1694700623
transform 1 0 2688 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_17
timestamp 1694700623
transform 1 0 3248 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_33
timestamp 1694700623
transform 1 0 5040 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_40
timestamp 1694700623
transform 1 0 5824 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_48
timestamp 1694700623
transform 1 0 6720 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_53
timestamp 1694700623
transform 1 0 7280 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_61
timestamp 1694700623
transform 1 0 8176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_65
timestamp 1694700623
transform 1 0 8624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_67
timestamp 1694700623
transform 1 0 8848 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_74
timestamp 1694700623
transform 1 0 9632 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_82
timestamp 1694700623
transform 1 0 10528 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_84
timestamp 1694700623
transform 1 0 10752 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_89
timestamp 1694700623
transform 1 0 11312 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_97
timestamp 1694700623
transform 1 0 12208 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_101
timestamp 1694700623
transform 1 0 12656 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_108
timestamp 1694700623
transform 1 0 13440 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_116
timestamp 1694700623
transform 1 0 14336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_120
timestamp 1694700623
transform 1 0 14784 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_125
timestamp 1694700623
transform 1 0 15344 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_133
timestamp 1694700623
transform 1 0 16240 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_135
timestamp 1694700623
transform 1 0 16464 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_138
timestamp 1694700623
transform 1 0 16800 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_143
timestamp 1694700623
transform 1 0 17360 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_172
timestamp 1694700623
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_176
timestamp 1694700623
transform 1 0 21056 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_206
timestamp 1694700623
transform 1 0 24416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_210
timestamp 1694700623
transform 1 0 24864 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_237
timestamp 1694700623
transform 1 0 27888 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_240
timestamp 1694700623
transform 1 0 28224 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_244
timestamp 1694700623
transform 1 0 28672 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_246
timestamp 1694700623
transform 1 0 28896 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_251
timestamp 1694700623
transform 1 0 29456 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_259
timestamp 1694700623
transform 1 0 30352 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_263
timestamp 1694700623
transform 1 0 30800 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_269
timestamp 1694700623
transform 1 0 31472 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_271
timestamp 1694700623
transform 1 0 31696 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_274
timestamp 1694700623
transform 1 0 32032 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_282
timestamp 1694700623
transform 1 0 32928 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_287
timestamp 1694700623
transform 1 0 33488 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_295
timestamp 1694700623
transform 1 0 34384 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_299
timestamp 1694700623
transform 1 0 34832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_305
timestamp 1694700623
transform 1 0 35504 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_308
timestamp 1694700623
transform 1 0 35840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_312
timestamp 1694700623
transform 1 0 36288 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_368
timestamp 1694700623
transform 1 0 42560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_402
timestamp 1694700623
transform 1 0 46368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_406
timestamp 1694700623
transform 1 0 46816 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_436
timestamp 1694700623
transform 1 0 50176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_440
timestamp 1694700623
transform 1 0 50624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_470
timestamp 1694700623
transform 1 0 53984 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_474
timestamp 1694700623
transform 1 0 54432 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_504
timestamp 1694700623
transform 1 0 57792 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_508
timestamp 1694700623
transform 1 0 58240 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1694700623
transform -1 0 58352 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1694700623
transform -1 0 58352 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1694700623
transform -1 0 58352 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1694700623
transform -1 0 58352 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1694700623
transform -1 0 58352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1694700623
transform -1 0 58352 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1694700623
transform -1 0 58352 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1694700623
transform -1 0 58352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1694700623
transform -1 0 58352 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1694700623
transform -1 0 58352 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1694700623
transform 1 0 1568 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1694700623
transform 1 0 1568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 24192 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1694700623
transform 1 0 24976 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1694700623
transform -1 0 29904 0 -1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1694700623
transform -1 0 39424 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1694700623
transform 1 0 39648 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1694700623
transform 1 0 41552 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1694700623
transform -1 0 46368 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1694700623
transform 1 0 47264 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1694700623
transform -1 0 50064 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1694700623
transform 1 0 51072 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1694700623
transform 1 0 51184 0 -1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1694700623
transform 1 0 54880 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1694700623
transform 1 0 55216 0 1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1694700623
transform 1 0 53312 0 -1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1694700623
transform 1 0 17472 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1694700623
transform 1 0 21168 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_81 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_82
timestamp 1694700623
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_83
timestamp 1694700623
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_84
timestamp 1694700623
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_85
timestamp 1694700623
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_86
timestamp 1694700623
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_87
timestamp 1694700623
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_88
timestamp 1694700623
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_89
timestamp 1694700623
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_90
timestamp 1694700623
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_91
timestamp 1694700623
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_92
timestamp 1694700623
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_93
timestamp 1694700623
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_94
timestamp 1694700623
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_95
timestamp 1694700623
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_96
timestamp 1694700623
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_97
timestamp 1694700623
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_98
timestamp 1694700623
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_99
timestamp 1694700623
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_100
timestamp 1694700623
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_101
timestamp 1694700623
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_102
timestamp 1694700623
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_103
timestamp 1694700623
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_104
timestamp 1694700623
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_105
timestamp 1694700623
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_106
timestamp 1694700623
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_107
timestamp 1694700623
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_108
timestamp 1694700623
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_109
timestamp 1694700623
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1694700623
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_110
timestamp 1694700623
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1694700623
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_111
timestamp 1694700623
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1694700623
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_112
timestamp 1694700623
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1694700623
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_113
timestamp 1694700623
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1694700623
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_114
timestamp 1694700623
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1694700623
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_115
timestamp 1694700623
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1694700623
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_116
timestamp 1694700623
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1694700623
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_117
timestamp 1694700623
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1694700623
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_118
timestamp 1694700623
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1694700623
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_119
timestamp 1694700623
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1694700623
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_120
timestamp 1694700623
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1694700623
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_121
timestamp 1694700623
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1694700623
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_122
timestamp 1694700623
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1694700623
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_123
timestamp 1694700623
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1694700623
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_124
timestamp 1694700623
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1694700623
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_125
timestamp 1694700623
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1694700623
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_126
timestamp 1694700623
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1694700623
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_127
timestamp 1694700623
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1694700623
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_128
timestamp 1694700623
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1694700623
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_129
timestamp 1694700623
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1694700623
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_130
timestamp 1694700623
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1694700623
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_131
timestamp 1694700623
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1694700623
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_132
timestamp 1694700623
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1694700623
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_133
timestamp 1694700623
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1694700623
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_134
timestamp 1694700623
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1694700623
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_135
timestamp 1694700623
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1694700623
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_136
timestamp 1694700623
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1694700623
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_137
timestamp 1694700623
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1694700623
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_138
timestamp 1694700623
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1694700623
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_139
timestamp 1694700623
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1694700623
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_140
timestamp 1694700623
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1694700623
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_141
timestamp 1694700623
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1694700623
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_142
timestamp 1694700623
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1694700623
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_143
timestamp 1694700623
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1694700623
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_144
timestamp 1694700623
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1694700623
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_145
timestamp 1694700623
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1694700623
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_146
timestamp 1694700623
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1694700623
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_147
timestamp 1694700623
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1694700623
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_148
timestamp 1694700623
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1694700623
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_149
timestamp 1694700623
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1694700623
transform -1 0 58576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_150
timestamp 1694700623
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1694700623
transform -1 0 58576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_151
timestamp 1694700623
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1694700623
transform -1 0 58576 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_152
timestamp 1694700623
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1694700623
transform -1 0 58576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_153
timestamp 1694700623
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1694700623
transform -1 0 58576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_154
timestamp 1694700623
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1694700623
transform -1 0 58576 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_155
timestamp 1694700623
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1694700623
transform -1 0 58576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_156
timestamp 1694700623
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1694700623
transform -1 0 58576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_157
timestamp 1694700623
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1694700623
transform -1 0 58576 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_158
timestamp 1694700623
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1694700623
transform -1 0 58576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_159
timestamp 1694700623
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1694700623
transform -1 0 58576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_160
timestamp 1694700623
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1694700623
transform -1 0 58576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_161
timestamp 1694700623
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1694700623
transform -1 0 58576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1694700623
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1694700623
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1694700623
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_166
timestamp 1694700623
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_167
timestamp 1694700623
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_168
timestamp 1694700623
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_169
timestamp 1694700623
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_170
timestamp 1694700623
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_171
timestamp 1694700623
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_172
timestamp 1694700623
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_173
timestamp 1694700623
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_174
timestamp 1694700623
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_175
timestamp 1694700623
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_176
timestamp 1694700623
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_177
timestamp 1694700623
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_178
timestamp 1694700623
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_179
timestamp 1694700623
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_180
timestamp 1694700623
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_181
timestamp 1694700623
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_182
timestamp 1694700623
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_183
timestamp 1694700623
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_184
timestamp 1694700623
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_185
timestamp 1694700623
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_186
timestamp 1694700623
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_187
timestamp 1694700623
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_188
timestamp 1694700623
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_189
timestamp 1694700623
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_190
timestamp 1694700623
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_191
timestamp 1694700623
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_192
timestamp 1694700623
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_193
timestamp 1694700623
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_194
timestamp 1694700623
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_195
timestamp 1694700623
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_196
timestamp 1694700623
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_197
timestamp 1694700623
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_198
timestamp 1694700623
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_199
timestamp 1694700623
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_200
timestamp 1694700623
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_201
timestamp 1694700623
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_202
timestamp 1694700623
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_203
timestamp 1694700623
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_204
timestamp 1694700623
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_205
timestamp 1694700623
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_206
timestamp 1694700623
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_207
timestamp 1694700623
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_208
timestamp 1694700623
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_209
timestamp 1694700623
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_210
timestamp 1694700623
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_211
timestamp 1694700623
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_212
timestamp 1694700623
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_213
timestamp 1694700623
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_214
timestamp 1694700623
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_215
timestamp 1694700623
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_216
timestamp 1694700623
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_217
timestamp 1694700623
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_218
timestamp 1694700623
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_219
timestamp 1694700623
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_220
timestamp 1694700623
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_221
timestamp 1694700623
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_222
timestamp 1694700623
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_223
timestamp 1694700623
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_224
timestamp 1694700623
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_225
timestamp 1694700623
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_226
timestamp 1694700623
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_227
timestamp 1694700623
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_228
timestamp 1694700623
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_229
timestamp 1694700623
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_230
timestamp 1694700623
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_231
timestamp 1694700623
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_232
timestamp 1694700623
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_233
timestamp 1694700623
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_234
timestamp 1694700623
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_235
timestamp 1694700623
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_236
timestamp 1694700623
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_237
timestamp 1694700623
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_238
timestamp 1694700623
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_239
timestamp 1694700623
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_240
timestamp 1694700623
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_241
timestamp 1694700623
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_242
timestamp 1694700623
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_243
timestamp 1694700623
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_244
timestamp 1694700623
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_245
timestamp 1694700623
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_246
timestamp 1694700623
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_247
timestamp 1694700623
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_248
timestamp 1694700623
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_249
timestamp 1694700623
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_250
timestamp 1694700623
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_251
timestamp 1694700623
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_252
timestamp 1694700623
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_253
timestamp 1694700623
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_254
timestamp 1694700623
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_255
timestamp 1694700623
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_256
timestamp 1694700623
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_257
timestamp 1694700623
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_258
timestamp 1694700623
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_259
timestamp 1694700623
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_260
timestamp 1694700623
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_261
timestamp 1694700623
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_262
timestamp 1694700623
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_263
timestamp 1694700623
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_264
timestamp 1694700623
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_265
timestamp 1694700623
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_266
timestamp 1694700623
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_267
timestamp 1694700623
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_268
timestamp 1694700623
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_269
timestamp 1694700623
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_270
timestamp 1694700623
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_271
timestamp 1694700623
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_272
timestamp 1694700623
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_273
timestamp 1694700623
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_274
timestamp 1694700623
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_275
timestamp 1694700623
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_276
timestamp 1694700623
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_277
timestamp 1694700623
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_278
timestamp 1694700623
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_279
timestamp 1694700623
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_280
timestamp 1694700623
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_281
timestamp 1694700623
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_282
timestamp 1694700623
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_283
timestamp 1694700623
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_284
timestamp 1694700623
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_285
timestamp 1694700623
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_286
timestamp 1694700623
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_287
timestamp 1694700623
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_288
timestamp 1694700623
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_289
timestamp 1694700623
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_290
timestamp 1694700623
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_291
timestamp 1694700623
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_292
timestamp 1694700623
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_293
timestamp 1694700623
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_294
timestamp 1694700623
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_295
timestamp 1694700623
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_296
timestamp 1694700623
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_297
timestamp 1694700623
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_298
timestamp 1694700623
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_299
timestamp 1694700623
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_300
timestamp 1694700623
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_301
timestamp 1694700623
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_302
timestamp 1694700623
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_303
timestamp 1694700623
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_304
timestamp 1694700623
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_305
timestamp 1694700623
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_306
timestamp 1694700623
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_307
timestamp 1694700623
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_308
timestamp 1694700623
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_309
timestamp 1694700623
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_310
timestamp 1694700623
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_311
timestamp 1694700623
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_312
timestamp 1694700623
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_313
timestamp 1694700623
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_314
timestamp 1694700623
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_315
timestamp 1694700623
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_316
timestamp 1694700623
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_317
timestamp 1694700623
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_318
timestamp 1694700623
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_319
timestamp 1694700623
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_320
timestamp 1694700623
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_321
timestamp 1694700623
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_322
timestamp 1694700623
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_323
timestamp 1694700623
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_324
timestamp 1694700623
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_325
timestamp 1694700623
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_326
timestamp 1694700623
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_327
timestamp 1694700623
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_328
timestamp 1694700623
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_329
timestamp 1694700623
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_330
timestamp 1694700623
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_331
timestamp 1694700623
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_332
timestamp 1694700623
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_333
timestamp 1694700623
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_334
timestamp 1694700623
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_335
timestamp 1694700623
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_336
timestamp 1694700623
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_337
timestamp 1694700623
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_338
timestamp 1694700623
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_339
timestamp 1694700623
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_340
timestamp 1694700623
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_341
timestamp 1694700623
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_342
timestamp 1694700623
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_343
timestamp 1694700623
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_344
timestamp 1694700623
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_345
timestamp 1694700623
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_346
timestamp 1694700623
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_347
timestamp 1694700623
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_348
timestamp 1694700623
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_349
timestamp 1694700623
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_350
timestamp 1694700623
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_351
timestamp 1694700623
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_352
timestamp 1694700623
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_353
timestamp 1694700623
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_354
timestamp 1694700623
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_355
timestamp 1694700623
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_356
timestamp 1694700623
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_357
timestamp 1694700623
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_358
timestamp 1694700623
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_359
timestamp 1694700623
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_360
timestamp 1694700623
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_361
timestamp 1694700623
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_362
timestamp 1694700623
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_363
timestamp 1694700623
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_364
timestamp 1694700623
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_365
timestamp 1694700623
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_366
timestamp 1694700623
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_367
timestamp 1694700623
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1694700623
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1694700623
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1694700623
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1694700623
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_372
timestamp 1694700623
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1694700623
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1694700623
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1694700623
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1694700623
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_377
timestamp 1694700623
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_378
timestamp 1694700623
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_379
timestamp 1694700623
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_380
timestamp 1694700623
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1694700623
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_382
timestamp 1694700623
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_383
timestamp 1694700623
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_384
timestamp 1694700623
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1694700623
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_386
timestamp 1694700623
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_387
timestamp 1694700623
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_388
timestamp 1694700623
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_389
timestamp 1694700623
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_390
timestamp 1694700623
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1694700623
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1694700623
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_393
timestamp 1694700623
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_394
timestamp 1694700623
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_395
timestamp 1694700623
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_396
timestamp 1694700623
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_397
timestamp 1694700623
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_398
timestamp 1694700623
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_399
timestamp 1694700623
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_400
timestamp 1694700623
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_401
timestamp 1694700623
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_402
timestamp 1694700623
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_403
timestamp 1694700623
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_404
timestamp 1694700623
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_405
timestamp 1694700623
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_406
timestamp 1694700623
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_407
timestamp 1694700623
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_408
timestamp 1694700623
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_409
timestamp 1694700623
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_410
timestamp 1694700623
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_411
timestamp 1694700623
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_412
timestamp 1694700623
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_413
timestamp 1694700623
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_414
timestamp 1694700623
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_415
timestamp 1694700623
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_416
timestamp 1694700623
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_417
timestamp 1694700623
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_418
timestamp 1694700623
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_419
timestamp 1694700623
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_420
timestamp 1694700623
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_421
timestamp 1694700623
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_422
timestamp 1694700623
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_423
timestamp 1694700623
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_424
timestamp 1694700623
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_425
timestamp 1694700623
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_426
timestamp 1694700623
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_427
timestamp 1694700623
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_428
timestamp 1694700623
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_429
timestamp 1694700623
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_430
timestamp 1694700623
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_431
timestamp 1694700623
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_432
timestamp 1694700623
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_433
timestamp 1694700623
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_434
timestamp 1694700623
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_435
timestamp 1694700623
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_436
timestamp 1694700623
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_437
timestamp 1694700623
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_438
timestamp 1694700623
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_439
timestamp 1694700623
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_440
timestamp 1694700623
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_441
timestamp 1694700623
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_442
timestamp 1694700623
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_443
timestamp 1694700623
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_444
timestamp 1694700623
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_445
timestamp 1694700623
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_446
timestamp 1694700623
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_447
timestamp 1694700623
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_448
timestamp 1694700623
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_449
timestamp 1694700623
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_450
timestamp 1694700623
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_451
timestamp 1694700623
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_452
timestamp 1694700623
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_453
timestamp 1694700623
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_454
timestamp 1694700623
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_455
timestamp 1694700623
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_456
timestamp 1694700623
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_457
timestamp 1694700623
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_458
timestamp 1694700623
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_459
timestamp 1694700623
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_460
timestamp 1694700623
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_461
timestamp 1694700623
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_462
timestamp 1694700623
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_463
timestamp 1694700623
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_464
timestamp 1694700623
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_465
timestamp 1694700623
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_466
timestamp 1694700623
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_467
timestamp 1694700623
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_468
timestamp 1694700623
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_469
timestamp 1694700623
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_470
timestamp 1694700623
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_471
timestamp 1694700623
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_472
timestamp 1694700623
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_473
timestamp 1694700623
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_474
timestamp 1694700623
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_475
timestamp 1694700623
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_476
timestamp 1694700623
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_477
timestamp 1694700623
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_478
timestamp 1694700623
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_479
timestamp 1694700623
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_480
timestamp 1694700623
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_481
timestamp 1694700623
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_482
timestamp 1694700623
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_483
timestamp 1694700623
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_484
timestamp 1694700623
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_485
timestamp 1694700623
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_486
timestamp 1694700623
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_487
timestamp 1694700623
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_488
timestamp 1694700623
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_489
timestamp 1694700623
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_490
timestamp 1694700623
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_491
timestamp 1694700623
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_492
timestamp 1694700623
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_493
timestamp 1694700623
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_494
timestamp 1694700623
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_495
timestamp 1694700623
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_496
timestamp 1694700623
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_497
timestamp 1694700623
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_498
timestamp 1694700623
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_499
timestamp 1694700623
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_500
timestamp 1694700623
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_501
timestamp 1694700623
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_502
timestamp 1694700623
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_503
timestamp 1694700623
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_504
timestamp 1694700623
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_505
timestamp 1694700623
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_506
timestamp 1694700623
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_507
timestamp 1694700623
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_508
timestamp 1694700623
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_509
timestamp 1694700623
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_510
timestamp 1694700623
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_511
timestamp 1694700623
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_512
timestamp 1694700623
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_513
timestamp 1694700623
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_514
timestamp 1694700623
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_515
timestamp 1694700623
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_516
timestamp 1694700623
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_517
timestamp 1694700623
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_518
timestamp 1694700623
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_519
timestamp 1694700623
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_520
timestamp 1694700623
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_521
timestamp 1694700623
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_522
timestamp 1694700623
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_523
timestamp 1694700623
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_524
timestamp 1694700623
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_525
timestamp 1694700623
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_526
timestamp 1694700623
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_527
timestamp 1694700623
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_528
timestamp 1694700623
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_529
timestamp 1694700623
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_530
timestamp 1694700623
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_531
timestamp 1694700623
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_532
timestamp 1694700623
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_533
timestamp 1694700623
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_534
timestamp 1694700623
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_535
timestamp 1694700623
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_536
timestamp 1694700623
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_537
timestamp 1694700623
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_538
timestamp 1694700623
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_539
timestamp 1694700623
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_540
timestamp 1694700623
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_541
timestamp 1694700623
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_542
timestamp 1694700623
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_543
timestamp 1694700623
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_544
timestamp 1694700623
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_545
timestamp 1694700623
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_546
timestamp 1694700623
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_547
timestamp 1694700623
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_548
timestamp 1694700623
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_549
timestamp 1694700623
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_550
timestamp 1694700623
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_551
timestamp 1694700623
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_552
timestamp 1694700623
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_553
timestamp 1694700623
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_554
timestamp 1694700623
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_555
timestamp 1694700623
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_556
timestamp 1694700623
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_557
timestamp 1694700623
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_558
timestamp 1694700623
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_559
timestamp 1694700623
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_560
timestamp 1694700623
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_561
timestamp 1694700623
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_562
timestamp 1694700623
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_563
timestamp 1694700623
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_564
timestamp 1694700623
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_565
timestamp 1694700623
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_566
timestamp 1694700623
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_567
timestamp 1694700623
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_568
timestamp 1694700623
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_569
timestamp 1694700623
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_570
timestamp 1694700623
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_571
timestamp 1694700623
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_572
timestamp 1694700623
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_573
timestamp 1694700623
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_574
timestamp 1694700623
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_575
timestamp 1694700623
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_576
timestamp 1694700623
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_577
timestamp 1694700623
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_578
timestamp 1694700623
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_579
timestamp 1694700623
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_580
timestamp 1694700623
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_581
timestamp 1694700623
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_582
timestamp 1694700623
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_583
timestamp 1694700623
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_584
timestamp 1694700623
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_585
timestamp 1694700623
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_586
timestamp 1694700623
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_587
timestamp 1694700623
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_588
timestamp 1694700623
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_589
timestamp 1694700623
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_590
timestamp 1694700623
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_591
timestamp 1694700623
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_592
timestamp 1694700623
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_593
timestamp 1694700623
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_594
timestamp 1694700623
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_595
timestamp 1694700623
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_596
timestamp 1694700623
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_597
timestamp 1694700623
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_598
timestamp 1694700623
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_599
timestamp 1694700623
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_600
timestamp 1694700623
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_601
timestamp 1694700623
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_602
timestamp 1694700623
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_603
timestamp 1694700623
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_604
timestamp 1694700623
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_605
timestamp 1694700623
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_606
timestamp 1694700623
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_607
timestamp 1694700623
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_608
timestamp 1694700623
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_609
timestamp 1694700623
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_610
timestamp 1694700623
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_611
timestamp 1694700623
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_612
timestamp 1694700623
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_613
timestamp 1694700623
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_614
timestamp 1694700623
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_615
timestamp 1694700623
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_616
timestamp 1694700623
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_617
timestamp 1694700623
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_618
timestamp 1694700623
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_619
timestamp 1694700623
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_620
timestamp 1694700623
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_621
timestamp 1694700623
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_622
timestamp 1694700623
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_623
timestamp 1694700623
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_624
timestamp 1694700623
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_625
timestamp 1694700623
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_626
timestamp 1694700623
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_627
timestamp 1694700623
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_628
timestamp 1694700623
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_629
timestamp 1694700623
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_630
timestamp 1694700623
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_631
timestamp 1694700623
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_632
timestamp 1694700623
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_633
timestamp 1694700623
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_634
timestamp 1694700623
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_635
timestamp 1694700623
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_636
timestamp 1694700623
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_637
timestamp 1694700623
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_638
timestamp 1694700623
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_639
timestamp 1694700623
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_640
timestamp 1694700623
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_641
timestamp 1694700623
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_642
timestamp 1694700623
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_643
timestamp 1694700623
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_644
timestamp 1694700623
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_645
timestamp 1694700623
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_646
timestamp 1694700623
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_647
timestamp 1694700623
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_648
timestamp 1694700623
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_649
timestamp 1694700623
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_650
timestamp 1694700623
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_651
timestamp 1694700623
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_652
timestamp 1694700623
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_653
timestamp 1694700623
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_654
timestamp 1694700623
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_655
timestamp 1694700623
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_656
timestamp 1694700623
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_657
timestamp 1694700623
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_658
timestamp 1694700623
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_659
timestamp 1694700623
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_660
timestamp 1694700623
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_661
timestamp 1694700623
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_662
timestamp 1694700623
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_663
timestamp 1694700623
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_664
timestamp 1694700623
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_665
timestamp 1694700623
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_666
timestamp 1694700623
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_667
timestamp 1694700623
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_668
timestamp 1694700623
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_669
timestamp 1694700623
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_670
timestamp 1694700623
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_671
timestamp 1694700623
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_672
timestamp 1694700623
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_673
timestamp 1694700623
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_674
timestamp 1694700623
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_675
timestamp 1694700623
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_676
timestamp 1694700623
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_677
timestamp 1694700623
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_678
timestamp 1694700623
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_679
timestamp 1694700623
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_680
timestamp 1694700623
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_681
timestamp 1694700623
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_682
timestamp 1694700623
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_683
timestamp 1694700623
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_684
timestamp 1694700623
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_685
timestamp 1694700623
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_686
timestamp 1694700623
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_687
timestamp 1694700623
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_688
timestamp 1694700623
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_689
timestamp 1694700623
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_690
timestamp 1694700623
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_691
timestamp 1694700623
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_692
timestamp 1694700623
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_693
timestamp 1694700623
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_694
timestamp 1694700623
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_695
timestamp 1694700623
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_696
timestamp 1694700623
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_697
timestamp 1694700623
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_698
timestamp 1694700623
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_699
timestamp 1694700623
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_700
timestamp 1694700623
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_701
timestamp 1694700623
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_702
timestamp 1694700623
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_703
timestamp 1694700623
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_704
timestamp 1694700623
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_705
timestamp 1694700623
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_706
timestamp 1694700623
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_707
timestamp 1694700623
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_708
timestamp 1694700623
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_709
timestamp 1694700623
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_710
timestamp 1694700623
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_711
timestamp 1694700623
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_712
timestamp 1694700623
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_713
timestamp 1694700623
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_714
timestamp 1694700623
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_715
timestamp 1694700623
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_716
timestamp 1694700623
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_717
timestamp 1694700623
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_718
timestamp 1694700623
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_719
timestamp 1694700623
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_720
timestamp 1694700623
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_721
timestamp 1694700623
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_722
timestamp 1694700623
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_723
timestamp 1694700623
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_724
timestamp 1694700623
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_725
timestamp 1694700623
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_726
timestamp 1694700623
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_727
timestamp 1694700623
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_728
timestamp 1694700623
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_729
timestamp 1694700623
transform 1 0 5152 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_730
timestamp 1694700623
transform 1 0 8960 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_731
timestamp 1694700623
transform 1 0 12768 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_732
timestamp 1694700623
transform 1 0 16576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_733
timestamp 1694700623
transform 1 0 20384 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_734
timestamp 1694700623
transform 1 0 24192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_735
timestamp 1694700623
transform 1 0 28000 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_736
timestamp 1694700623
transform 1 0 31808 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_737
timestamp 1694700623
transform 1 0 35616 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_738
timestamp 1694700623
transform 1 0 39424 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_739
timestamp 1694700623
transform 1 0 43232 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_740
timestamp 1694700623
transform 1 0 47040 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_741
timestamp 1694700623
transform 1 0 50848 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_742
timestamp 1694700623
transform 1 0 54656 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1694700623
transform -1 0 3248 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_30
timestamp 1694700623
transform -1 0 5824 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_31
timestamp 1694700623
transform -1 0 7280 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_32
timestamp 1694700623
transform -1 0 9632 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_33
timestamp 1694700623
transform -1 0 11312 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_34
timestamp 1694700623
transform -1 0 13440 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_35
timestamp 1694700623
transform -1 0 15344 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_36
timestamp 1694700623
transform -1 0 17360 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_37
timestamp 1694700623
transform -1 0 29456 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_38
timestamp 1694700623
transform -1 0 31472 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_39
timestamp 1694700623
transform -1 0 33488 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_40
timestamp 1694700623
transform -1 0 35504 0 1 65856
box -86 -86 534 870
<< labels >>
flabel metal3 s 59200 59136 60000 59248 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 59200 66080 60000 66192 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 59200 3584 60000 3696 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 59200 10528 60000 10640 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 59200 17472 60000 17584 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 59200 24416 60000 24528 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 59200 31360 60000 31472 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 59200 38304 60000 38416 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 59200 45248 60000 45360 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 59200 52192 60000 52304 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 io_in_2
port 10 nsew signal input
flabel metal2 s 2688 69200 2800 70000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 22848 69200 22960 70000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 24864 69200 24976 70000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 26880 69200 26992 70000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 28896 69200 29008 70000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 30912 69200 31024 70000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 32928 69200 33040 70000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 34944 69200 35056 70000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 36960 69200 37072 70000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 38976 69200 39088 70000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 40992 69200 41104 70000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 4704 69200 4816 70000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 43008 69200 43120 70000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 45024 69200 45136 70000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 47040 69200 47152 70000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 49056 69200 49168 70000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 51072 69200 51184 70000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 53088 69200 53200 70000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 55104 69200 55216 70000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 57120 69200 57232 70000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 6720 69200 6832 70000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 8736 69200 8848 70000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 10752 69200 10864 70000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 12768 69200 12880 70000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 14784 69200 14896 70000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 16800 69200 16912 70000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 18816 69200 18928 70000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 20832 69200 20944 70000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 rst_n
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 66700 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 66700 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 66700 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 66700 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal3 s 0 11648 800 11760 0 FreeSans 448 0 0 0 wb_clk_i
port 42 nsew signal input
rlabel metal1 29960 66640 29960 66640 0 vdd
rlabel metal1 29960 65856 29960 65856 0 vss
rlabel metal2 47600 64344 47600 64344 0 _0000_
rlabel metal2 29624 10192 29624 10192 0 _0001_
rlabel metal2 29848 7784 29848 7784 0 _0002_
rlabel metal2 31080 5264 31080 5264 0 _0003_
rlabel metal2 31528 5264 31528 5264 0 _0004_
rlabel metal2 47768 5488 47768 5488 0 _0005_
rlabel metal2 45528 8456 45528 8456 0 _0006_
rlabel metal2 45080 4424 45080 4424 0 _0007_
rlabel metal2 43736 6048 43736 6048 0 _0008_
rlabel metal2 47544 22288 47544 22288 0 _0009_
rlabel metal2 47880 19600 47880 19600 0 _0010_
rlabel metal2 45864 18760 45864 18760 0 _0011_
rlabel metal2 45864 22736 45864 22736 0 _0012_
rlabel metal2 41160 40824 41160 40824 0 _0013_
rlabel metal2 41272 36904 41272 36904 0 _0014_
rlabel metal3 21056 43400 21056 43400 0 _0015_
rlabel metal2 23688 49392 23688 49392 0 _0016_
rlabel metal3 18760 49112 18760 49112 0 _0017_
rlabel metal2 18200 53256 18200 53256 0 _0018_
rlabel metal2 21336 53032 21336 53032 0 _0019_
rlabel metal2 22120 57288 22120 57288 0 _0020_
rlabel metal2 22624 60200 22624 60200 0 _0021_
rlabel metal2 17864 56336 17864 56336 0 _0022_
rlabel metal2 20552 59248 20552 59248 0 _0023_
rlabel metal2 2520 36680 2520 36680 0 _0024_
rlabel metal2 2520 40488 2520 40488 0 _0025_
rlabel metal2 2632 44072 2632 44072 0 _0026_
rlabel metal2 2632 47096 2632 47096 0 _0027_
rlabel metal2 2520 50232 2520 50232 0 _0028_
rlabel metal2 2520 54656 2520 54656 0 _0029_
rlabel metal2 2520 57960 2520 57960 0 _0030_
rlabel metal3 5600 59416 5600 59416 0 _0031_
rlabel metal2 6664 63896 6664 63896 0 _0032_
rlabel metal2 21000 61320 21000 61320 0 _0033_
rlabel metal2 19656 63952 19656 63952 0 _0034_
rlabel metal2 5320 37576 5320 37576 0 _0035_
rlabel metal2 6104 42224 6104 42224 0 _0036_
rlabel metal2 7336 44688 7336 44688 0 _0037_
rlabel metal2 12152 46816 12152 46816 0 _0038_
rlabel metal3 8064 48888 8064 48888 0 _0039_
rlabel metal2 5992 53256 5992 53256 0 _0040_
rlabel metal2 7448 57064 7448 57064 0 _0041_
rlabel metal2 11816 60032 11816 60032 0 _0042_
rlabel metal3 11480 64792 11480 64792 0 _0043_
rlabel metal2 14952 63560 14952 63560 0 _0044_
rlabel metal2 17640 64736 17640 64736 0 _0045_
rlabel metal2 54264 39088 54264 39088 0 _0046_
rlabel metal2 53592 47096 53592 47096 0 _0047_
rlabel metal2 57176 45472 57176 45472 0 _0048_
rlabel metal2 53816 42112 53816 42112 0 _0049_
rlabel metal2 50848 45192 50848 45192 0 _0050_
rlabel metal2 49896 41608 49896 41608 0 _0051_
rlabel metal2 51016 39312 51016 39312 0 _0052_
rlabel metal3 48496 31640 48496 31640 0 _0053_
rlabel metal2 49112 29848 49112 29848 0 _0054_
rlabel metal2 52808 27440 52808 27440 0 _0055_
rlabel metal2 50232 25032 50232 25032 0 _0056_
rlabel metal2 51464 23464 51464 23464 0 _0057_
rlabel metal2 54376 21728 54376 21728 0 _0058_
rlabel metal2 56056 20944 56056 20944 0 _0059_
rlabel metal2 57288 24472 57288 24472 0 _0060_
rlabel metal3 56560 26488 56560 26488 0 _0061_
rlabel metal2 56056 30744 56056 30744 0 _0062_
rlabel metal2 56112 31864 56112 31864 0 _0063_
rlabel metal3 56616 36232 56616 36232 0 _0064_
rlabel metal2 55160 36120 55160 36120 0 _0065_
rlabel metal3 52752 33208 52752 33208 0 _0066_
rlabel metal2 49112 32984 49112 32984 0 _0067_
rlabel metal2 49112 25816 49112 25816 0 _0068_
rlabel metal2 43288 25928 43288 25928 0 _0069_
rlabel metal2 41832 28560 41832 28560 0 _0070_
rlabel metal2 43064 31696 43064 31696 0 _0071_
rlabel metal2 39592 32088 39592 32088 0 _0072_
rlabel metal2 44856 35840 44856 35840 0 _0073_
rlabel metal2 47320 34384 47320 34384 0 _0074_
rlabel metal2 46648 37688 46648 37688 0 _0075_
rlabel metal2 45864 40880 45864 40880 0 _0076_
rlabel metal2 33992 44520 33992 44520 0 _0077_
rlabel metal3 32648 45752 32648 45752 0 _0078_
rlabel metal3 28448 50456 28448 50456 0 _0079_
rlabel metal2 26040 53872 26040 53872 0 _0080_
rlabel metal3 33096 56952 33096 56952 0 _0081_
rlabel metal3 25536 63224 25536 63224 0 _0082_
rlabel metal2 29064 63168 29064 63168 0 _0083_
rlabel metal2 35672 65072 35672 65072 0 _0084_
rlabel metal3 23072 64904 23072 64904 0 _0085_
rlabel metal2 51800 11200 51800 11200 0 _0086_
rlabel metal2 56504 17976 56504 17976 0 _0087_
rlabel metal2 57400 16464 57400 16464 0 _0088_
rlabel metal2 56504 14840 56504 14840 0 _0089_
rlabel metal3 54040 13608 54040 13608 0 _0090_
rlabel metal3 48384 11480 48384 11480 0 _0091_
rlabel metal3 44296 10696 44296 10696 0 _0092_
rlabel metal2 42504 14532 42504 14532 0 _0093_
rlabel metal2 40208 11480 40208 11480 0 _0094_
rlabel metal2 38584 22288 38584 22288 0 _0095_
rlabel metal2 27944 33712 27944 33712 0 _0096_
rlabel metal2 54488 9352 54488 9352 0 _0097_
rlabel metal3 53704 6664 53704 6664 0 _0098_
rlabel metal2 52696 4648 52696 4648 0 _0099_
rlabel metal3 41272 4424 41272 4424 0 _0100_
rlabel metal2 38248 4816 38248 4816 0 _0101_
rlabel metal2 36456 5040 36456 5040 0 _0102_
rlabel metal2 33544 5432 33544 5432 0 _0103_
rlabel metal2 30296 12320 30296 12320 0 _0104_
rlabel metal2 36008 12320 36008 12320 0 _0105_
rlabel metal2 35784 15792 35784 15792 0 _0106_
rlabel metal2 8344 25872 8344 25872 0 _0107_
rlabel metal2 26824 11928 26824 11928 0 _0108_
rlabel metal2 26040 4648 26040 4648 0 _0109_
rlabel metal2 22456 4648 22456 4648 0 _0110_
rlabel metal2 19208 4648 19208 4648 0 _0111_
rlabel metal2 17416 6328 17416 6328 0 _0112_
rlabel metal2 14728 9352 14728 9352 0 _0113_
rlabel metal2 15848 11032 15848 11032 0 _0114_
rlabel metal2 14728 13888 14728 13888 0 _0115_
rlabel metal2 23800 11704 23800 11704 0 _0116_
rlabel metal2 24584 15484 24584 15484 0 _0117_
rlabel metal3 17304 33208 17304 33208 0 _0118_
rlabel metal2 46648 43876 46648 43876 0 _0119_
rlabel metal2 41496 43932 41496 43932 0 _0120_
rlabel metal2 45528 45640 45528 45640 0 _0121_
rlabel metal2 39592 46200 39592 46200 0 _0122_
rlabel metal2 40712 50904 40712 50904 0 _0123_
rlabel metal2 39592 54936 39592 54936 0 _0124_
rlabel metal3 46144 58520 46144 58520 0 _0125_
rlabel metal2 39256 58800 39256 58800 0 _0126_
rlabel metal2 43624 64512 43624 64512 0 _0127_
rlabel metal2 46144 62216 46144 62216 0 _0128_
rlabel metal2 57400 63448 57400 63448 0 _0129_
rlabel metal3 57064 59416 57064 59416 0 _0130_
rlabel metal2 57344 64568 57344 64568 0 _0131_
rlabel metal3 52528 54712 52528 54712 0 _0132_
rlabel metal2 55944 48664 55944 48664 0 _0133_
rlabel metal2 56056 51296 56056 51296 0 _0134_
rlabel metal2 55384 55412 55384 55412 0 _0135_
rlabel metal2 56000 53816 56000 53816 0 _0136_
rlabel metal2 51240 52640 51240 52640 0 _0137_
rlabel metal2 53032 48552 53032 48552 0 _0138_
rlabel metal2 48888 49336 48888 49336 0 _0139_
rlabel metal2 44968 50960 44968 50960 0 _0140_
rlabel metal2 48888 51800 48888 51800 0 _0141_
rlabel metal2 43288 52528 43288 52528 0 _0142_
rlabel metal2 45640 55608 45640 55608 0 _0143_
rlabel metal2 48888 56504 48888 56504 0 _0144_
rlabel metal2 48104 59640 48104 59640 0 _0145_
rlabel metal2 49392 62216 49392 62216 0 _0146_
rlabel metal2 50232 65128 50232 65128 0 _0147_
rlabel metal2 51800 65128 51800 65128 0 _0148_
rlabel metal2 52136 58856 52136 58856 0 _0149_
rlabel metal2 51632 56168 51632 56168 0 _0150_
rlabel metal3 50176 36344 50176 36344 0 _0151_
rlabel metal2 41496 22008 41496 22008 0 _0152_
rlabel metal3 41832 19880 41832 19880 0 _0153_
rlabel metal2 42224 17752 42224 17752 0 _0154_
rlabel metal2 38528 17640 38528 17640 0 _0155_
rlabel metal2 36008 18480 36008 18480 0 _0156_
rlabel metal2 34440 22008 34440 22008 0 _0157_
rlabel metal2 27384 15456 27384 15456 0 _0158_
rlabel metal2 28000 13832 28000 13832 0 _0159_
rlabel metal2 29288 20356 29288 20356 0 _0160_
rlabel metal2 26040 18592 26040 18592 0 _0161_
rlabel metal2 30408 17024 30408 17024 0 _0162_
rlabel metal2 31360 20216 31360 20216 0 _0163_
rlabel metal2 16632 16576 16632 16576 0 _0164_
rlabel metal2 14728 17192 14728 17192 0 _0165_
rlabel metal3 17136 20664 17136 20664 0 _0166_
rlabel metal3 16632 18424 16632 18424 0 _0167_
rlabel metal2 20664 17024 20664 17024 0 _0168_
rlabel metal2 20272 20104 20272 20104 0 _0169_
rlabel metal2 31752 27440 31752 27440 0 _0170_
rlabel metal2 31864 28728 31864 28728 0 _0171_
rlabel metal2 29176 30576 29176 30576 0 _0172_
rlabel metal2 26488 29680 26488 29680 0 _0173_
rlabel metal2 25032 30968 25032 30968 0 _0174_
rlabel metal2 21560 30352 21560 30352 0 _0175_
rlabel metal2 22120 33264 22120 33264 0 _0176_
rlabel metal2 20328 28616 20328 28616 0 _0177_
rlabel metal3 9912 29288 9912 29288 0 _0178_
rlabel metal2 5544 28168 5544 28168 0 _0179_
rlabel metal3 12824 25368 12824 25368 0 _0180_
rlabel metal3 12432 24584 12432 24584 0 _0181_
rlabel metal2 16464 29288 16464 29288 0 _0182_
rlabel metal2 17584 25368 17584 25368 0 _0183_
rlabel metal2 17528 28280 17528 28280 0 _0184_
rlabel metal2 16128 23240 16128 23240 0 _0185_
rlabel metal2 20552 24864 20552 24864 0 _0186_
rlabel metal2 22512 21672 22512 21672 0 _0187_
rlabel metal2 30072 23464 30072 23464 0 _0188_
rlabel metal3 43960 26376 43960 26376 0 _0189_
rlabel metal2 36120 25032 36120 25032 0 _0190_
rlabel metal2 37240 29848 37240 29848 0 _0191_
rlabel metal2 39480 28112 39480 28112 0 _0192_
rlabel metal2 8680 56952 8680 56952 0 _0193_
rlabel metal2 47656 46480 47656 46480 0 _0194_
rlabel metal2 10248 56840 10248 56840 0 _0195_
rlabel metal2 10472 56560 10472 56560 0 _0196_
rlabel metal2 11816 58352 11816 58352 0 _0197_
rlabel metal2 12040 59024 12040 59024 0 _0198_
rlabel metal2 11144 60704 11144 60704 0 _0199_
rlabel metal2 12936 60760 12936 60760 0 _0200_
rlabel metal2 11816 62328 11816 62328 0 _0201_
rlabel metal2 11368 64344 11368 64344 0 _0202_
rlabel metal3 13272 64008 13272 64008 0 _0203_
rlabel metal2 13720 63000 13720 63000 0 _0204_
rlabel metal2 12936 62776 12936 62776 0 _0205_
rlabel metal3 16408 63112 16408 63112 0 _0206_
rlabel metal2 14840 62720 14840 62720 0 _0207_
rlabel metal2 16744 63224 16744 63224 0 _0208_
rlabel metal2 39312 34104 39312 34104 0 _0209_
rlabel metal2 19544 52724 19544 52724 0 _0210_
rlabel metal2 17528 63336 17528 63336 0 _0211_
rlabel metal2 56840 39200 56840 39200 0 _0212_
rlabel metal3 52472 11368 52472 11368 0 _0213_
rlabel metal2 53928 46648 53928 46648 0 _0214_
rlabel metal2 57288 61488 57288 61488 0 _0215_
rlabel metal2 56840 45192 56840 45192 0 _0216_
rlabel metal2 56168 44800 56168 44800 0 _0217_
rlabel metal2 53704 43680 53704 43680 0 _0218_
rlabel metal2 53592 43288 53592 43288 0 _0219_
rlabel metal2 47936 26264 47936 26264 0 _0220_
rlabel metal2 51240 45136 51240 45136 0 _0221_
rlabel metal3 51184 41160 51184 41160 0 _0222_
rlabel metal2 48944 48104 48944 48104 0 _0223_
rlabel metal2 49672 48048 49672 48048 0 _0224_
rlabel metal2 51688 42728 51688 42728 0 _0225_
rlabel metal2 50344 42168 50344 42168 0 _0226_
rlabel metal2 51352 40040 51352 40040 0 _0227_
rlabel metal2 39144 33320 39144 33320 0 _0228_
rlabel metal2 50120 35112 50120 35112 0 _0229_
rlabel metal2 53256 35168 53256 35168 0 _0230_
rlabel metal2 53200 29624 53200 29624 0 _0231_
rlabel metal2 50232 30408 50232 30408 0 _0232_
rlabel metal2 49896 31416 49896 31416 0 _0233_
rlabel metal2 50120 28224 50120 28224 0 _0234_
rlabel metal2 50120 31808 50120 31808 0 _0235_
rlabel metal2 51240 29680 51240 29680 0 _0236_
rlabel metal2 52192 32648 52192 32648 0 _0237_
rlabel metal2 53480 24752 53480 24752 0 _0238_
rlabel metal2 53256 29008 53256 29008 0 _0239_
rlabel metal2 53144 25032 53144 25032 0 _0240_
rlabel metal2 53816 24696 53816 24696 0 _0241_
rlabel metal3 53256 26936 53256 26936 0 _0242_
rlabel metal2 52360 26684 52360 26684 0 _0243_
rlabel metal3 53256 25480 53256 25480 0 _0244_
rlabel metal2 52584 25200 52584 25200 0 _0245_
rlabel metal2 53088 23912 53088 23912 0 _0246_
rlabel metal2 53368 24192 53368 24192 0 _0247_
rlabel metal2 54936 22792 54936 22792 0 _0248_
rlabel metal2 56896 25368 56896 25368 0 _0249_
rlabel metal3 55832 22232 55832 22232 0 _0250_
rlabel metal2 57176 21840 57176 21840 0 _0251_
rlabel metal3 57288 23240 57288 23240 0 _0252_
rlabel metal2 56952 21896 56952 21896 0 _0253_
rlabel metal2 56504 21840 56504 21840 0 _0254_
rlabel metal2 56952 24024 56952 24024 0 _0255_
rlabel metal2 56448 24696 56448 24696 0 _0256_
rlabel metal3 57456 27608 57456 27608 0 _0257_
rlabel metal2 57288 26572 57288 26572 0 _0258_
rlabel metal2 56728 30296 56728 30296 0 _0259_
rlabel metal2 55048 33432 55048 33432 0 _0260_
rlabel metal2 57288 32256 57288 32256 0 _0261_
rlabel metal3 56000 30968 56000 30968 0 _0262_
rlabel metal3 53760 34664 53760 34664 0 _0263_
rlabel metal2 57064 33824 57064 33824 0 _0264_
rlabel metal2 56728 34440 56728 34440 0 _0265_
rlabel metal2 58072 36176 58072 36176 0 _0266_
rlabel metal2 57512 36176 57512 36176 0 _0267_
rlabel metal3 55944 35672 55944 35672 0 _0268_
rlabel metal2 54712 35000 54712 35000 0 _0269_
rlabel metal2 53872 32312 53872 32312 0 _0270_
rlabel metal2 51800 32816 51800 32816 0 _0271_
rlabel metal2 46536 31416 46536 31416 0 _0272_
rlabel metal3 48216 32536 48216 32536 0 _0273_
rlabel metal3 50064 32536 50064 32536 0 _0274_
rlabel metal2 57624 40320 57624 40320 0 _0275_
rlabel metal2 55944 40768 55944 40768 0 _0276_
rlabel metal2 57064 40096 57064 40096 0 _0277_
rlabel metal2 55720 40880 55720 40880 0 _0278_
rlabel metal2 57064 42448 57064 42448 0 _0279_
rlabel metal2 49784 12712 49784 12712 0 _0280_
rlabel metal2 40040 14336 40040 14336 0 _0281_
rlabel metal3 46984 25592 46984 25592 0 _0282_
rlabel metal2 50288 46536 50288 46536 0 _0283_
rlabel metal4 57512 41104 57512 41104 0 _0284_
rlabel metal2 45864 25592 45864 25592 0 _0285_
rlabel metal3 35392 15848 35392 15848 0 _0286_
rlabel metal2 38696 11480 38696 11480 0 _0287_
rlabel metal2 46872 10360 46872 10360 0 _0288_
rlabel metal2 44184 14280 44184 14280 0 _0289_
rlabel metal2 43960 25872 43960 25872 0 _0290_
rlabel metal3 44688 26936 44688 26936 0 _0291_
rlabel metal2 44128 26824 44128 26824 0 _0292_
rlabel metal2 44016 31976 44016 31976 0 _0293_
rlabel metal2 43456 28728 43456 28728 0 _0294_
rlabel metal2 43904 33320 43904 33320 0 _0295_
rlabel metal2 43736 33768 43736 33768 0 _0296_
rlabel metal2 44744 32536 44744 32536 0 _0297_
rlabel metal3 43848 32424 43848 32424 0 _0298_
rlabel metal2 44296 34552 44296 34552 0 _0299_
rlabel metal2 41664 33320 41664 33320 0 _0300_
rlabel metal2 44072 35224 44072 35224 0 _0301_
rlabel metal3 45192 34104 45192 34104 0 _0302_
rlabel metal2 44968 35728 44968 35728 0 _0303_
rlabel metal2 46816 33992 46816 33992 0 _0304_
rlabel metal2 45864 39144 45864 39144 0 _0305_
rlabel metal2 46536 37408 46536 37408 0 _0306_
rlabel metal3 45640 39592 45640 39592 0 _0307_
rlabel metal3 44688 39480 44688 39480 0 _0308_
rlabel metal2 45304 40320 45304 40320 0 _0309_
rlabel metal2 44632 40096 44632 40096 0 _0310_
rlabel metal2 44184 41328 44184 41328 0 _0311_
rlabel metal2 44184 41944 44184 41944 0 _0312_
rlabel metal3 33432 44296 33432 44296 0 _0313_
rlabel metal2 34552 44296 34552 44296 0 _0314_
rlabel metal2 37240 22288 37240 22288 0 _0315_
rlabel metal2 31752 44800 31752 44800 0 _0316_
rlabel metal2 32480 43736 32480 43736 0 _0317_
rlabel metal2 31080 46480 31080 46480 0 _0318_
rlabel metal3 31584 46536 31584 46536 0 _0319_
rlabel metal2 29736 47432 29736 47432 0 _0320_
rlabel metal2 29008 46648 29008 46648 0 _0321_
rlabel metal2 29288 47936 29288 47936 0 _0322_
rlabel metal2 28504 50204 28504 50204 0 _0323_
rlabel metal2 29568 50008 29568 50008 0 _0324_
rlabel metal3 30184 50680 30184 50680 0 _0325_
rlabel metal3 29288 50008 29288 50008 0 _0326_
rlabel metal2 30184 50204 30184 50204 0 _0327_
rlabel metal2 29400 54824 29400 54824 0 _0328_
rlabel metal3 26796 54600 26796 54600 0 _0329_
rlabel metal2 28560 62888 28560 62888 0 _0330_
rlabel metal2 27272 54376 27272 54376 0 _0331_
rlabel metal2 29736 54152 29736 54152 0 _0332_
rlabel metal2 29512 54992 29512 54992 0 _0333_
rlabel metal2 30184 57232 30184 57232 0 _0334_
rlabel metal2 31864 57512 31864 57512 0 _0335_
rlabel metal2 29960 57568 29960 57568 0 _0336_
rlabel metal2 30856 57512 30856 57512 0 _0337_
rlabel metal2 27272 62552 27272 62552 0 _0338_
rlabel metal2 27048 63336 27048 63336 0 _0339_
rlabel metal3 26936 63112 26936 63112 0 _0340_
rlabel metal2 27832 63448 27832 63448 0 _0341_
rlabel metal2 27440 64008 27440 64008 0 _0342_
rlabel metal3 29960 64680 29960 64680 0 _0343_
rlabel metal2 29512 62944 29512 62944 0 _0344_
rlabel metal2 29400 62832 29400 62832 0 _0345_
rlabel metal2 32872 63616 32872 63616 0 _0346_
rlabel metal2 32648 63560 32648 63560 0 _0347_
rlabel metal2 34664 64176 34664 64176 0 _0348_
rlabel metal2 35168 64008 35168 64008 0 _0349_
rlabel metal2 32312 63504 32312 63504 0 _0350_
rlabel metal2 32088 63560 32088 63560 0 _0351_
rlabel metal2 23688 64176 23688 64176 0 _0352_
rlabel metal2 50344 12880 50344 12880 0 _0353_
rlabel metal2 51912 11760 51912 11760 0 _0354_
rlabel metal2 50904 10080 50904 10080 0 _0355_
rlabel metal2 51688 16464 51688 16464 0 _0356_
rlabel metal2 47768 15680 47768 15680 0 _0357_
rlabel metal2 49336 16520 49336 16520 0 _0358_
rlabel metal2 51296 14280 51296 14280 0 _0359_
rlabel metal2 51464 11256 51464 11256 0 _0360_
rlabel metal2 49560 10416 49560 10416 0 _0361_
rlabel metal2 51744 14392 51744 14392 0 _0362_
rlabel metal2 51520 17864 51520 17864 0 _0363_
rlabel metal3 52976 18200 52976 18200 0 _0364_
rlabel metal2 39144 14168 39144 14168 0 _0365_
rlabel metal2 20888 12712 20888 12712 0 _0366_
rlabel metal3 51912 18424 51912 18424 0 _0367_
rlabel metal3 53872 18312 53872 18312 0 _0368_
rlabel metal2 52136 17472 52136 17472 0 _0369_
rlabel metal3 53480 17864 53480 17864 0 _0370_
rlabel metal2 52024 16912 52024 16912 0 _0371_
rlabel metal2 53424 17416 53424 17416 0 _0372_
rlabel metal3 46480 15848 46480 15848 0 _0373_
rlabel metal2 52584 15232 52584 15232 0 _0374_
rlabel metal3 51800 14616 51800 14616 0 _0375_
rlabel metal2 52584 14728 52584 14728 0 _0376_
rlabel metal3 52360 14280 52360 14280 0 _0377_
rlabel metal2 53704 14868 53704 14868 0 _0378_
rlabel metal3 49952 14728 49952 14728 0 _0379_
rlabel metal3 50736 14504 50736 14504 0 _0380_
rlabel metal2 50120 8036 50120 8036 0 _0381_
rlabel metal2 50848 13944 50848 13944 0 _0382_
rlabel metal3 52304 13720 52304 13720 0 _0383_
rlabel metal2 51072 6664 51072 6664 0 _0384_
rlabel metal2 47656 14616 47656 14616 0 _0385_
rlabel metal2 47544 13664 47544 13664 0 _0386_
rlabel metal2 48216 13216 48216 13216 0 _0387_
rlabel metal2 47768 12320 47768 12320 0 _0388_
rlabel metal2 45080 15624 45080 15624 0 _0389_
rlabel metal2 45136 14504 45136 14504 0 _0390_
rlabel metal2 44968 13384 44968 13384 0 _0391_
rlabel metal2 44072 14112 44072 14112 0 _0392_
rlabel metal2 44856 13440 44856 13440 0 _0393_
rlabel metal2 44744 12488 44744 12488 0 _0394_
rlabel metal2 42560 13720 42560 13720 0 _0395_
rlabel metal2 41160 13328 41160 13328 0 _0396_
rlabel metal2 41496 14840 41496 14840 0 _0397_
rlabel metal3 40264 14392 40264 14392 0 _0398_
rlabel metal2 41272 12432 41272 12432 0 _0399_
rlabel metal2 41496 14056 41496 14056 0 _0400_
rlabel metal2 39648 13720 39648 13720 0 _0401_
rlabel metal2 39872 12152 39872 12152 0 _0402_
rlabel metal2 51016 12096 51016 12096 0 _0403_
rlabel metal2 39256 12040 39256 12040 0 _0404_
rlabel metal2 39592 12264 39592 12264 0 _0405_
rlabel metal2 28896 26152 28896 26152 0 _0406_
rlabel metal2 38360 22288 38360 22288 0 _0407_
rlabel metal2 37464 21952 37464 21952 0 _0408_
rlabel metal2 28392 33488 28392 33488 0 _0409_
rlabel metal3 52304 9800 52304 9800 0 _0410_
rlabel metal3 45696 8008 45696 8008 0 _0411_
rlabel metal3 38472 9688 38472 9688 0 _0412_
rlabel metal2 47320 8176 47320 8176 0 _0413_
rlabel metal3 50680 8344 50680 8344 0 _0414_
rlabel metal2 52584 9744 52584 9744 0 _0415_
rlabel metal3 49000 8120 49000 8120 0 _0416_
rlabel metal3 51184 7448 51184 7448 0 _0417_
rlabel metal2 50456 7448 50456 7448 0 _0418_
rlabel metal2 50792 7056 50792 7056 0 _0419_
rlabel metal3 52024 7336 52024 7336 0 _0420_
rlabel metal2 49280 6776 49280 6776 0 _0421_
rlabel metal3 49448 6608 49448 6608 0 _0422_
rlabel metal2 50344 7112 50344 7112 0 _0423_
rlabel metal2 51184 5208 51184 5208 0 _0424_
rlabel metal2 39368 7672 39368 7672 0 _0425_
rlabel metal3 39816 9184 39816 9184 0 _0426_
rlabel metal3 40768 7672 40768 7672 0 _0427_
rlabel metal2 40768 6888 40768 6888 0 _0428_
rlabel metal2 38920 7784 38920 7784 0 _0429_
rlabel metal2 40936 6944 40936 6944 0 _0430_
rlabel metal2 40712 5488 40712 5488 0 _0431_
rlabel metal2 37744 7448 37744 7448 0 _0432_
rlabel metal2 38808 6944 38808 6944 0 _0433_
rlabel metal2 38920 7056 38920 7056 0 _0434_
rlabel metal2 38136 5432 38136 5432 0 _0435_
rlabel metal2 35448 8456 35448 8456 0 _0436_
rlabel metal2 35000 7616 35000 7616 0 _0437_
rlabel metal2 36064 7448 36064 7448 0 _0438_
rlabel metal3 25200 6440 25200 6440 0 _0439_
rlabel metal2 35504 5992 35504 5992 0 _0440_
rlabel metal2 32536 15624 32536 15624 0 _0441_
rlabel metal2 33544 9352 33544 9352 0 _0442_
rlabel metal2 33768 7728 33768 7728 0 _0443_
rlabel metal2 33544 12656 33544 12656 0 _0444_
rlabel metal3 33152 7448 33152 7448 0 _0445_
rlabel metal2 33880 6272 33880 6272 0 _0446_
rlabel metal2 31640 11984 31640 11984 0 _0447_
rlabel metal2 33656 13104 33656 13104 0 _0448_
rlabel metal2 34832 13160 34832 13160 0 _0449_
rlabel metal2 32312 11760 32312 11760 0 _0450_
rlabel metal2 32704 11368 32704 11368 0 _0451_
rlabel metal2 34776 13832 34776 13832 0 _0452_
rlabel metal2 35000 13440 35000 13440 0 _0453_
rlabel metal2 34776 12432 34776 12432 0 _0454_
rlabel metal2 34552 12600 34552 12600 0 _0455_
rlabel metal3 41384 46536 41384 46536 0 _0456_
rlabel metal2 9576 26208 9576 26208 0 _0457_
rlabel metal2 33992 15512 33992 15512 0 _0458_
rlabel metal2 35336 15680 35336 15680 0 _0459_
rlabel metal2 46200 46200 46200 46200 0 _0460_
rlabel metal2 8792 25704 8792 25704 0 _0461_
rlabel metal2 27496 12096 27496 12096 0 _0462_
rlabel metal2 24808 8736 24808 8736 0 _0463_
rlabel metal2 19880 10024 19880 10024 0 _0464_
rlabel metal2 26712 9856 26712 9856 0 _0465_
rlabel metal3 26628 7448 26628 7448 0 _0466_
rlabel metal2 27272 11480 27272 11480 0 _0467_
rlabel metal3 20496 6552 20496 6552 0 _0468_
rlabel metal2 26768 7560 26768 7560 0 _0469_
rlabel metal2 23800 6832 23800 6832 0 _0470_
rlabel metal2 26824 7896 26824 7896 0 _0471_
rlabel metal2 26152 5824 26152 5824 0 _0472_
rlabel metal2 23576 5936 23576 5936 0 _0473_
rlabel metal2 21336 7224 21336 7224 0 _0474_
rlabel metal2 20328 6384 20328 6384 0 _0475_
rlabel metal2 23576 6104 23576 6104 0 _0476_
rlabel metal2 23240 5992 23240 5992 0 _0477_
rlabel metal2 21560 11032 21560 11032 0 _0478_
rlabel metal2 20776 6272 20776 6272 0 _0479_
rlabel metal2 20216 7168 20216 7168 0 _0480_
rlabel metal3 21000 6664 21000 6664 0 _0481_
rlabel metal2 19320 6496 19320 6496 0 _0482_
rlabel metal2 20216 5992 20216 5992 0 _0483_
rlabel metal2 18984 7672 18984 7672 0 _0484_
rlabel metal3 18592 9128 18592 9128 0 _0485_
rlabel metal2 18984 5712 18984 5712 0 _0486_
rlabel metal2 17584 5992 17584 5992 0 _0487_
rlabel metal2 18088 10024 18088 10024 0 _0488_
rlabel metal3 18648 12712 18648 12712 0 _0489_
rlabel metal2 18872 9296 18872 9296 0 _0490_
rlabel metal3 17304 9912 17304 9912 0 _0491_
rlabel metal2 18872 12992 18872 12992 0 _0492_
rlabel metal3 18984 12824 18984 12824 0 _0493_
rlabel metal2 19544 12320 19544 12320 0 _0494_
rlabel metal2 19992 12936 19992 12936 0 _0495_
rlabel metal2 19656 12376 19656 12376 0 _0496_
rlabel metal2 15960 10920 15960 10920 0 _0497_
rlabel metal2 20552 13440 20552 13440 0 _0498_
rlabel metal2 18984 13608 18984 13608 0 _0499_
rlabel metal2 21280 13160 21280 13160 0 _0500_
rlabel metal2 21448 13384 21448 13384 0 _0501_
rlabel metal3 20328 13720 20328 13720 0 _0502_
rlabel metal2 23352 13776 23352 13776 0 _0503_
rlabel metal2 24472 13272 24472 13272 0 _0504_
rlabel metal2 23016 12768 23016 12768 0 _0505_
rlabel metal3 23408 12936 23408 12936 0 _0506_
rlabel metal3 21448 16184 21448 16184 0 _0507_
rlabel metal2 23688 15512 23688 15512 0 _0508_
rlabel metal2 24248 15680 24248 15680 0 _0509_
rlabel metal2 19544 33040 19544 33040 0 _0510_
rlabel metal2 46536 44408 46536 44408 0 _0511_
rlabel metal2 46872 44408 46872 44408 0 _0512_
rlabel metal2 44184 42896 44184 42896 0 _0513_
rlabel metal2 34888 41496 34888 41496 0 _0514_
rlabel metal2 39256 42392 39256 42392 0 _0515_
rlabel metal2 43960 43932 43960 43932 0 _0516_
rlabel metal2 41888 42616 41888 42616 0 _0517_
rlabel metal2 43904 41720 43904 41720 0 _0518_
rlabel metal2 44520 44296 44520 44296 0 _0519_
rlabel metal2 45976 46928 45976 46928 0 _0520_
rlabel metal3 44100 46648 44100 46648 0 _0521_
rlabel metal3 45584 46648 45584 46648 0 _0522_
rlabel metal2 45080 46200 45080 46200 0 _0523_
rlabel metal2 42560 49000 42560 49000 0 _0524_
rlabel metal2 42392 48552 42392 48552 0 _0525_
rlabel metal2 42504 47712 42504 47712 0 _0526_
rlabel metal3 42784 49672 42784 49672 0 _0527_
rlabel metal2 41216 46760 41216 46760 0 _0528_
rlabel metal2 41944 49448 41944 49448 0 _0529_
rlabel metal2 41272 49672 41272 49672 0 _0530_
rlabel metal3 41608 50008 41608 50008 0 _0531_
rlabel metal3 41888 49784 41888 49784 0 _0532_
rlabel metal3 41440 50792 41440 50792 0 _0533_
rlabel metal2 41384 50204 41384 50204 0 _0534_
rlabel metal3 41496 51128 41496 51128 0 _0535_
rlabel metal2 41272 54152 41272 54152 0 _0536_
rlabel metal2 40040 54208 40040 54208 0 _0537_
rlabel metal3 40152 54600 40152 54600 0 _0538_
rlabel metal2 39648 43680 39648 43680 0 _0539_
rlabel metal2 39928 54152 39928 54152 0 _0540_
rlabel metal3 43624 63896 43624 63896 0 _0541_
rlabel metal2 42504 54768 42504 54768 0 _0542_
rlabel metal2 42728 57008 42728 57008 0 _0543_
rlabel metal2 42952 56392 42952 56392 0 _0544_
rlabel metal2 43624 57344 43624 57344 0 _0545_
rlabel metal2 44968 58408 44968 58408 0 _0546_
rlabel metal3 42728 59304 42728 59304 0 _0547_
rlabel metal2 42616 58744 42616 58744 0 _0548_
rlabel metal3 42280 59192 42280 59192 0 _0549_
rlabel metal3 40712 60536 40712 60536 0 _0550_
rlabel metal2 40936 59528 40936 59528 0 _0551_
rlabel metal2 41496 59528 41496 59528 0 _0552_
rlabel metal3 43820 62328 43820 62328 0 _0553_
rlabel metal3 42896 61432 42896 61432 0 _0554_
rlabel metal2 43008 62328 43008 62328 0 _0555_
rlabel metal2 42504 62272 42504 62272 0 _0556_
rlabel metal2 43288 63056 43288 63056 0 _0557_
rlabel metal2 45528 62664 45528 62664 0 _0558_
rlabel metal2 44744 62720 44744 62720 0 _0559_
rlabel metal2 44744 62328 44744 62328 0 _0560_
rlabel metal3 45360 62328 45360 62328 0 _0561_
rlabel metal2 46536 62384 46536 62384 0 _0562_
rlabel metal2 45192 63560 45192 63560 0 _0563_
rlabel metal2 47096 62552 47096 62552 0 _0564_
rlabel metal3 52528 64120 52528 64120 0 _0565_
rlabel metal2 55048 62104 55048 62104 0 _0566_
rlabel metal2 54656 63336 54656 63336 0 _0567_
rlabel metal2 53592 63616 53592 63616 0 _0568_
rlabel metal2 54376 62216 54376 62216 0 _0569_
rlabel metal2 56616 59976 56616 59976 0 _0570_
rlabel metal2 56952 61544 56952 61544 0 _0571_
rlabel metal3 57512 60648 57512 60648 0 _0572_
rlabel metal2 52864 51576 52864 51576 0 _0573_
rlabel metal2 51688 54208 51688 54208 0 _0574_
rlabel metal2 54488 51688 54488 51688 0 _0575_
rlabel metal3 55160 48328 55160 48328 0 _0576_
rlabel metal2 56728 51968 56728 51968 0 _0577_
rlabel metal2 55160 55720 55160 55720 0 _0578_
rlabel metal2 55608 56280 55608 56280 0 _0579_
rlabel metal2 56056 54320 56056 54320 0 _0580_
rlabel metal2 50736 51912 50736 51912 0 _0581_
rlabel metal2 53032 49280 53032 49280 0 _0582_
rlabel metal2 54488 53592 54488 53592 0 _0583_
rlabel metal3 53648 50792 53648 50792 0 _0584_
rlabel metal2 47656 50960 47656 50960 0 _0585_
rlabel metal2 47320 49952 47320 49952 0 _0586_
rlabel metal2 44576 46424 44576 46424 0 _0587_
rlabel metal2 45528 51408 45528 51408 0 _0588_
rlabel metal3 51688 53648 51688 53648 0 _0589_
rlabel metal2 51240 53984 51240 53984 0 _0590_
rlabel metal2 48776 51520 48776 51520 0 _0591_
rlabel metal2 43848 52472 43848 52472 0 _0592_
rlabel metal2 47208 55776 47208 55776 0 _0593_
rlabel metal2 46648 55328 46648 55328 0 _0594_
rlabel metal3 48496 56168 48496 56168 0 _0595_
rlabel metal2 51464 62104 51464 62104 0 _0596_
rlabel metal3 50232 63112 50232 63112 0 _0597_
rlabel metal3 48888 59304 48888 59304 0 _0598_
rlabel metal2 49672 61208 49672 61208 0 _0599_
rlabel metal2 50400 64120 50400 64120 0 _0600_
rlabel metal2 51688 63896 51688 63896 0 _0601_
rlabel metal2 52024 59136 52024 59136 0 _0602_
rlabel metal3 52416 56504 52416 56504 0 _0603_
rlabel metal2 31360 24920 31360 24920 0 _0604_
rlabel metal2 31864 24528 31864 24528 0 _0605_
rlabel metal2 27888 22232 27888 22232 0 _0606_
rlabel metal2 26936 21952 26936 21952 0 _0607_
rlabel metal3 23912 25368 23912 25368 0 _0608_
rlabel metal2 25424 22232 25424 22232 0 _0609_
rlabel metal2 28504 21952 28504 21952 0 _0610_
rlabel metal2 37128 20440 37128 20440 0 _0611_
rlabel metal2 33992 21616 33992 21616 0 _0612_
rlabel metal2 41832 22064 41832 22064 0 _0613_
rlabel metal2 33656 18704 33656 18704 0 _0614_
rlabel metal3 36680 18984 36680 18984 0 _0615_
rlabel metal2 42168 19656 42168 19656 0 _0616_
rlabel metal2 35952 21560 35952 21560 0 _0617_
rlabel metal3 42000 18424 42000 18424 0 _0618_
rlabel metal2 39704 18872 39704 18872 0 _0619_
rlabel metal2 30968 17696 30968 17696 0 _0620_
rlabel metal2 37800 19208 37800 19208 0 _0621_
rlabel via2 33656 25256 33656 25256 0 _0622_
rlabel metal3 30968 23352 30968 23352 0 _0623_
rlabel metal2 30408 18816 30408 18816 0 _0624_
rlabel metal3 35280 21560 35280 21560 0 _0625_
rlabel metal2 25368 23408 25368 23408 0 _0626_
rlabel metal2 27216 26488 27216 26488 0 _0627_
rlabel metal2 28056 22120 28056 22120 0 _0628_
rlabel metal2 29064 20468 29064 20468 0 _0629_
rlabel metal3 29680 19992 29680 19992 0 _0630_
rlabel metal3 28896 15960 28896 15960 0 _0631_
rlabel metal2 28168 17024 28168 17024 0 _0632_
rlabel metal2 28280 16800 28280 16800 0 _0633_
rlabel metal2 29400 20832 29400 20832 0 _0634_
rlabel metal3 28000 18648 28000 18648 0 _0635_
rlabel metal2 29904 20552 29904 20552 0 _0636_
rlabel metal2 19432 24472 19432 24472 0 _0637_
rlabel metal2 29064 18368 29064 18368 0 _0638_
rlabel metal3 27888 18424 27888 18424 0 _0639_
rlabel metal3 31416 17640 31416 17640 0 _0640_
rlabel metal3 31864 20104 31864 20104 0 _0641_
rlabel metal3 22680 21784 22680 21784 0 _0642_
rlabel metal2 18312 21224 18312 21224 0 _0643_
rlabel metal2 20104 21224 20104 21224 0 _0644_
rlabel metal2 19208 16968 19208 16968 0 _0645_
rlabel metal2 22344 18368 22344 18368 0 _0646_
rlabel metal2 18200 17640 18200 17640 0 _0647_
rlabel metal2 21896 20356 21896 20356 0 _0648_
rlabel metal2 18536 20272 18536 20272 0 _0649_
rlabel metal2 18536 18648 18536 18648 0 _0650_
rlabel metal2 21896 17976 21896 17976 0 _0651_
rlabel metal3 28168 25200 28168 25200 0 _0652_
rlabel metal3 21392 20664 21392 20664 0 _0653_
rlabel metal2 31024 25368 31024 25368 0 _0654_
rlabel metal2 25368 26656 25368 26656 0 _0655_
rlabel metal2 32424 25704 32424 25704 0 _0656_
rlabel metal3 27440 26264 27440 26264 0 _0657_
rlabel metal2 26152 26040 26152 26040 0 _0658_
rlabel metal2 26488 26684 26488 26684 0 _0659_
rlabel metal2 28168 27552 28168 27552 0 _0660_
rlabel metal2 30632 29120 30632 29120 0 _0661_
rlabel metal2 28840 29008 28840 29008 0 _0662_
rlabel metal2 31304 28336 31304 28336 0 _0663_
rlabel metal2 31080 29568 31080 29568 0 _0664_
rlabel metal2 25256 29456 25256 29456 0 _0665_
rlabel metal2 29624 30184 29624 30184 0 _0666_
rlabel metal3 28112 29512 28112 29512 0 _0667_
rlabel metal2 27888 26040 27888 26040 0 _0668_
rlabel metal2 25648 23352 25648 23352 0 _0669_
rlabel metal2 26208 25592 26208 25592 0 _0670_
rlabel metal2 24584 28336 24584 28336 0 _0671_
rlabel metal2 22344 30576 22344 30576 0 _0672_
rlabel metal3 23072 29512 23072 29512 0 _0673_
rlabel metal2 24584 30520 24584 30520 0 _0674_
rlabel metal2 22008 30240 22008 30240 0 _0675_
rlabel metal2 21112 29512 21112 29512 0 _0676_
rlabel metal3 22288 30968 22288 30968 0 _0677_
rlabel metal3 21840 29512 21840 29512 0 _0678_
rlabel metal2 27496 26320 27496 26320 0 _0679_
rlabel metal2 25704 26600 25704 26600 0 _0680_
rlabel metal3 20552 26376 20552 26376 0 _0681_
rlabel metal2 13832 25256 13832 25256 0 _0682_
rlabel metal2 14672 27832 14672 27832 0 _0683_
rlabel metal2 15008 27608 15008 27608 0 _0684_
rlabel metal2 14224 28056 14224 28056 0 _0685_
rlabel metal2 14504 25984 14504 25984 0 _0686_
rlabel metal2 14280 25704 14280 25704 0 _0687_
rlabel metal2 14392 24640 14392 24640 0 _0688_
rlabel metal2 27272 25816 27272 25816 0 _0689_
rlabel metal2 17752 25872 17752 25872 0 _0690_
rlabel metal3 16408 24920 16408 24920 0 _0691_
rlabel metal2 17416 25928 17416 25928 0 _0692_
rlabel metal3 16912 29512 16912 29512 0 _0693_
rlabel metal3 18032 24696 18032 24696 0 _0694_
rlabel metal2 39144 27776 39144 27776 0 _0695_
rlabel metal2 17752 28168 17752 28168 0 _0696_
rlabel metal2 16520 24976 16520 24976 0 _0697_
rlabel metal2 28280 24248 28280 24248 0 _0698_
rlabel metal2 22344 24696 22344 24696 0 _0699_
rlabel metal3 23632 23128 23632 23128 0 _0700_
rlabel metal2 29120 24024 29120 24024 0 _0701_
rlabel metal2 38472 25984 38472 25984 0 _0702_
rlabel metal2 37016 26180 37016 26180 0 _0703_
rlabel metal2 38192 25592 38192 25592 0 _0704_
rlabel metal2 37912 29064 37912 29064 0 _0705_
rlabel metal2 38920 28616 38920 28616 0 _0706_
rlabel metal3 38752 27944 38752 27944 0 _0707_
rlabel metal2 22792 36176 22792 36176 0 _0708_
rlabel metal2 26152 38248 26152 38248 0 _0709_
rlabel metal2 24136 38724 24136 38724 0 _0710_
rlabel metal2 26040 37576 26040 37576 0 _0711_
rlabel metal2 27160 37632 27160 37632 0 _0712_
rlabel metal2 26600 37632 26600 37632 0 _0713_
rlabel metal2 27608 40320 27608 40320 0 _0714_
rlabel metal2 23352 40880 23352 40880 0 _0715_
rlabel metal2 25592 39144 25592 39144 0 _0716_
rlabel metal2 22680 39872 22680 39872 0 _0717_
rlabel metal2 25032 39592 25032 39592 0 _0718_
rlabel metal2 24472 41272 24472 41272 0 _0719_
rlabel metal3 23520 37912 23520 37912 0 _0720_
rlabel metal2 31304 41496 31304 41496 0 _0721_
rlabel metal2 31192 40376 31192 40376 0 _0722_
rlabel metal2 23688 39200 23688 39200 0 _0723_
rlabel metal2 24696 37688 24696 37688 0 _0724_
rlabel metal2 24248 37744 24248 37744 0 _0725_
rlabel metal2 23464 41160 23464 41160 0 _0726_
rlabel metal3 23912 40432 23912 40432 0 _0727_
rlabel metal3 31584 40936 31584 40936 0 _0728_
rlabel metal3 38248 31752 38248 31752 0 _0729_
rlabel metal3 37408 34104 37408 34104 0 _0730_
rlabel metal3 33264 35672 33264 35672 0 _0731_
rlabel metal2 33880 33656 33880 33656 0 _0732_
rlabel metal2 34664 30072 34664 30072 0 _0733_
rlabel metal2 38920 32312 38920 32312 0 _0734_
rlabel metal2 34104 35728 34104 35728 0 _0735_
rlabel metal2 39256 36176 39256 36176 0 _0736_
rlabel metal3 36064 33096 36064 33096 0 _0737_
rlabel metal2 39424 35672 39424 35672 0 _0738_
rlabel metal2 37688 32480 37688 32480 0 _0739_
rlabel metal3 34608 37240 34608 37240 0 _0740_
rlabel metal2 37352 32984 37352 32984 0 _0741_
rlabel metal2 33040 39368 33040 39368 0 _0742_
rlabel metal3 33992 41048 33992 41048 0 _0743_
rlabel metal3 31304 31752 31304 31752 0 _0744_
rlabel metal2 31976 35056 31976 35056 0 _0745_
rlabel metal2 36232 36400 36232 36400 0 _0746_
rlabel metal3 32368 38696 32368 38696 0 _0747_
rlabel metal2 34888 39144 34888 39144 0 _0748_
rlabel metal2 35896 41104 35896 41104 0 _0749_
rlabel metal2 19600 35000 19600 35000 0 _0750_
rlabel metal2 17584 40376 17584 40376 0 _0751_
rlabel metal2 20440 37632 20440 37632 0 _0752_
rlabel metal3 18032 37912 18032 37912 0 _0753_
rlabel metal2 18872 36064 18872 36064 0 _0754_
rlabel metal2 16464 34888 16464 34888 0 _0755_
rlabel metal2 15960 35224 15960 35224 0 _0756_
rlabel metal3 17304 38136 17304 38136 0 _0757_
rlabel metal2 18872 38864 18872 38864 0 _0758_
rlabel metal2 16800 38248 16800 38248 0 _0759_
rlabel metal2 15232 40936 15232 40936 0 _0760_
rlabel metal2 12936 39536 12936 39536 0 _0761_
rlabel metal2 18704 38136 18704 38136 0 _0762_
rlabel metal3 18200 38696 18200 38696 0 _0763_
rlabel metal2 15848 38752 15848 38752 0 _0764_
rlabel metal2 17360 37240 17360 37240 0 _0765_
rlabel metal2 12264 39256 12264 39256 0 _0766_
rlabel metal2 11032 28448 11032 28448 0 _0767_
rlabel metal3 9912 28056 9912 28056 0 _0768_
rlabel metal2 7952 30072 7952 30072 0 _0769_
rlabel metal2 9352 32256 9352 32256 0 _0770_
rlabel metal3 8680 30296 8680 30296 0 _0771_
rlabel metal2 9912 31808 9912 31808 0 _0772_
rlabel metal2 11144 30800 11144 30800 0 _0773_
rlabel metal2 10472 29344 10472 29344 0 _0774_
rlabel metal2 11368 34496 11368 34496 0 _0775_
rlabel metal2 10920 32928 10920 32928 0 _0776_
rlabel metal2 14840 26852 14840 26852 0 _0777_
rlabel metal2 11256 29120 11256 29120 0 _0778_
rlabel metal3 11256 38696 11256 38696 0 _0779_
rlabel metal2 12936 30576 12936 30576 0 _0780_
rlabel metal2 11928 28896 11928 28896 0 _0781_
rlabel metal2 12264 32816 12264 32816 0 _0782_
rlabel metal2 12824 32088 12824 32088 0 _0783_
rlabel metal3 12880 38808 12880 38808 0 _0784_
rlabel metal2 13944 42840 13944 42840 0 _0785_
rlabel metal3 24024 39312 24024 39312 0 _0786_
rlabel metal2 36904 41832 36904 41832 0 _0787_
rlabel metal2 40376 40824 40376 40824 0 _0788_
rlabel metal2 37128 40432 37128 40432 0 _0789_
rlabel metal2 37240 42224 37240 42224 0 _0790_
rlabel metal2 37128 43232 37128 43232 0 _0791_
rlabel metal3 25144 38808 25144 38808 0 _0792_
rlabel metal2 25704 39200 25704 39200 0 _0793_
rlabel metal2 26824 38472 26824 38472 0 _0794_
rlabel metal2 34888 28672 34888 28672 0 _0795_
rlabel metal2 37688 36680 37688 36680 0 _0796_
rlabel metal2 39032 36288 39032 36288 0 _0797_
rlabel metal2 38136 36960 38136 36960 0 _0798_
rlabel metal2 37464 37464 37464 37464 0 _0799_
rlabel metal2 36848 36456 36848 36456 0 _0800_
rlabel metal2 43400 40096 43400 40096 0 _0801_
rlabel metal2 38808 41216 38808 41216 0 _0802_
rlabel metal2 21504 40600 21504 40600 0 _0803_
rlabel metal3 19096 41160 19096 41160 0 _0804_
rlabel metal3 18424 41272 18424 41272 0 _0805_
rlabel metal2 15960 41048 15960 41048 0 _0806_
rlabel metal2 21112 40432 21112 40432 0 _0807_
rlabel metal2 14000 41048 14000 41048 0 _0808_
rlabel metal2 21448 41776 21448 41776 0 _0809_
rlabel metal2 17416 42616 17416 42616 0 _0810_
rlabel metal2 11704 42056 11704 42056 0 _0811_
rlabel metal2 14392 27832 14392 27832 0 _0812_
rlabel metal2 13944 33768 13944 33768 0 _0813_
rlabel metal2 12824 29680 12824 29680 0 _0814_
rlabel metal2 14280 26992 14280 26992 0 _0815_
rlabel metal2 14280 30632 14280 30632 0 _0816_
rlabel metal2 12264 32088 12264 32088 0 _0817_
rlabel metal2 11032 41104 11032 41104 0 _0818_
rlabel metal2 38920 41888 38920 41888 0 _0819_
rlabel metal2 39480 42280 39480 42280 0 _0820_
rlabel metal2 39144 46984 39144 46984 0 _0821_
rlabel metal2 38864 37016 38864 37016 0 _0822_
rlabel metal2 37464 42728 37464 42728 0 _0823_
rlabel metal2 37464 45136 37464 45136 0 _0824_
rlabel metal2 10024 29064 10024 29064 0 _0825_
rlabel metal3 13832 41944 13832 41944 0 _0826_
rlabel metal2 14056 42056 14056 42056 0 _0827_
rlabel metal2 14504 42448 14504 42448 0 _0828_
rlabel metal2 14672 47208 14672 47208 0 _0829_
rlabel metal2 17864 46256 17864 46256 0 _0830_
rlabel metal2 8568 32984 8568 32984 0 _0831_
rlabel metal2 8904 35112 8904 35112 0 _0832_
rlabel metal2 9800 26684 9800 26684 0 _0833_
rlabel metal2 9632 33880 9632 33880 0 _0834_
rlabel metal3 10024 35672 10024 35672 0 _0835_
rlabel metal2 11088 36456 11088 36456 0 _0836_
rlabel metal3 11760 36232 11760 36232 0 _0837_
rlabel metal2 12152 35784 12152 35784 0 _0838_
rlabel metal3 15316 44296 15316 44296 0 _0839_
rlabel metal2 18872 40376 18872 40376 0 _0840_
rlabel metal3 16968 39592 16968 39592 0 _0841_
rlabel metal3 19376 34104 19376 34104 0 _0842_
rlabel metal2 20776 42168 20776 42168 0 _0843_
rlabel metal3 16016 41160 16016 41160 0 _0844_
rlabel metal2 16520 39368 16520 39368 0 _0845_
rlabel metal3 16968 40152 16968 40152 0 _0846_
rlabel metal3 16856 44296 16856 44296 0 _0847_
rlabel metal2 17752 45864 17752 45864 0 _0848_
rlabel metal2 35112 37016 35112 37016 0 _0849_
rlabel metal2 37464 34048 37464 34048 0 _0850_
rlabel metal2 32536 41216 32536 41216 0 _0851_
rlabel metal2 31304 37352 31304 37352 0 _0852_
rlabel metal2 32088 34552 32088 34552 0 _0853_
rlabel metal2 32984 37128 32984 37128 0 _0854_
rlabel metal2 25816 44688 25816 44688 0 _0855_
rlabel metal2 25256 41664 25256 41664 0 _0856_
rlabel metal2 25480 41048 25480 41048 0 _0857_
rlabel metal2 25592 41216 25592 41216 0 _0858_
rlabel metal2 25928 41552 25928 41552 0 _0859_
rlabel metal2 27944 40544 27944 40544 0 _0860_
rlabel metal3 28168 42728 28168 42728 0 _0861_
rlabel metal3 25088 44296 25088 44296 0 _0862_
rlabel metal2 25256 45920 25256 45920 0 _0863_
rlabel metal3 20160 46368 20160 46368 0 _0864_
rlabel metal2 39032 47264 39032 47264 0 _0865_
rlabel metal2 36456 47152 36456 47152 0 _0866_
rlabel metal2 37688 47320 37688 47320 0 _0867_
rlabel metal3 23688 47208 23688 47208 0 _0868_
rlabel metal2 25592 44576 25592 44576 0 _0869_
rlabel metal2 24472 44520 24472 44520 0 _0870_
rlabel metal2 24136 45976 24136 45976 0 _0871_
rlabel metal2 34776 46816 34776 46816 0 _0872_
rlabel metal2 35112 34048 35112 34048 0 _0873_
rlabel metal2 32424 34328 32424 34328 0 _0874_
rlabel metal2 33656 34440 33656 34440 0 _0875_
rlabel metal2 29288 44968 29288 44968 0 _0876_
rlabel metal2 23912 41440 23912 41440 0 _0877_
rlabel metal2 26600 41440 26600 41440 0 _0878_
rlabel metal2 26040 38472 26040 38472 0 _0879_
rlabel metal2 26712 40040 26712 40040 0 _0880_
rlabel metal3 27160 45864 27160 45864 0 _0881_
rlabel metal2 26152 47768 26152 47768 0 _0882_
rlabel metal2 13160 33320 13160 33320 0 _0883_
rlabel metal3 13384 34776 13384 34776 0 _0884_
rlabel metal2 14616 43008 14616 43008 0 _0885_
rlabel metal3 16240 42728 16240 42728 0 _0886_
rlabel metal2 18480 39928 18480 39928 0 _0887_
rlabel metal2 19432 41664 19432 41664 0 _0888_
rlabel metal2 14952 43960 14952 43960 0 _0889_
rlabel metal2 26040 46592 26040 46592 0 _0890_
rlabel metal2 15624 44800 15624 44800 0 _0891_
rlabel metal2 9744 45080 9744 45080 0 _0892_
rlabel metal3 16464 45864 16464 45864 0 _0893_
rlabel metal2 26264 46144 26264 46144 0 _0894_
rlabel metal2 34664 47488 34664 47488 0 _0895_
rlabel metal2 36680 47880 36680 47880 0 _0896_
rlabel metal2 35336 47040 35336 47040 0 _0897_
rlabel metal2 37240 49000 37240 49000 0 _0898_
rlabel metal2 26824 46928 26824 46928 0 _0899_
rlabel metal2 29400 46928 29400 46928 0 _0900_
rlabel metal3 24304 48104 24304 48104 0 _0901_
rlabel metal2 28168 47656 28168 47656 0 _0902_
rlabel metal2 34888 49560 34888 49560 0 _0903_
rlabel metal2 28392 42784 28392 42784 0 _0904_
rlabel metal3 31360 49000 31360 49000 0 _0905_
rlabel metal3 31528 39368 31528 39368 0 _0906_
rlabel metal2 32200 45192 32200 45192 0 _0907_
rlabel metal2 32760 49448 32760 49448 0 _0908_
rlabel metal2 14280 48608 14280 48608 0 _0909_
rlabel metal2 13888 50344 13888 50344 0 _0910_
rlabel metal2 15624 49280 15624 49280 0 _0911_
rlabel metal2 15400 47096 15400 47096 0 _0912_
rlabel metal2 13720 47600 13720 47600 0 _0913_
rlabel metal2 11144 48552 11144 48552 0 _0914_
rlabel metal2 15960 47824 15960 47824 0 _0915_
rlabel metal2 15680 47544 15680 47544 0 _0916_
rlabel metal2 16296 49168 16296 49168 0 _0917_
rlabel metal2 35168 49784 35168 49784 0 _0918_
rlabel metal2 38696 50512 38696 50512 0 _0919_
rlabel metal2 38696 51800 38696 51800 0 _0920_
rlabel metal2 35504 50008 35504 50008 0 _0921_
rlabel metal2 36008 53424 36008 53424 0 _0922_
rlabel metal2 19208 49560 19208 49560 0 _0923_
rlabel metal2 32424 50036 32424 50036 0 _0924_
rlabel metal2 33320 49896 33320 49896 0 _0925_
rlabel metal3 34552 52136 34552 52136 0 _0926_
rlabel metal2 28056 42056 28056 42056 0 _0927_
rlabel metal2 30408 44408 30408 44408 0 _0928_
rlabel metal2 30408 38976 30408 38976 0 _0929_
rlabel metal2 31528 52528 31528 52528 0 _0930_
rlabel metal2 33768 52472 33768 52472 0 _0931_
rlabel metal2 15064 51072 15064 51072 0 _0932_
rlabel metal2 15288 49840 15288 49840 0 _0933_
rlabel metal2 15512 37744 15512 37744 0 _0934_
rlabel metal2 13552 44520 13552 44520 0 _0935_
rlabel metal2 9072 37240 9072 37240 0 _0936_
rlabel metal2 9688 34832 9688 34832 0 _0937_
rlabel metal2 8904 37352 8904 37352 0 _0938_
rlabel metal2 12096 40936 12096 40936 0 _0939_
rlabel metal2 14560 51352 14560 51352 0 _0940_
rlabel metal2 15176 51632 15176 51632 0 _0941_
rlabel metal2 15960 52360 15960 52360 0 _0942_
rlabel metal2 32536 51968 32536 51968 0 _0943_
rlabel metal3 36400 52920 36400 52920 0 _0944_
rlabel metal2 36232 53424 36232 53424 0 _0945_
rlabel metal2 42056 54152 42056 54152 0 _0946_
rlabel metal2 30968 32312 30968 32312 0 _0947_
rlabel metal2 30072 34496 30072 34496 0 _0948_
rlabel metal2 29736 35336 29736 35336 0 _0949_
rlabel metal2 31416 34944 31416 34944 0 _0950_
rlabel metal2 31752 44296 31752 44296 0 _0951_
rlabel metal2 26824 37296 26824 37296 0 _0952_
rlabel metal2 29232 40936 29232 40936 0 _0953_
rlabel metal2 29064 41552 29064 41552 0 _0954_
rlabel metal2 28616 42056 28616 42056 0 _0955_
rlabel metal2 29008 42504 29008 42504 0 _0956_
rlabel metal2 29120 47656 29120 47656 0 _0957_
rlabel metal2 32312 55216 32312 55216 0 _0958_
rlabel metal2 17304 43624 17304 43624 0 _0959_
rlabel metal2 20552 42112 20552 42112 0 _0960_
rlabel metal2 17864 43232 17864 43232 0 _0961_
rlabel metal2 16856 44856 16856 44856 0 _0962_
rlabel metal3 11928 37352 11928 37352 0 _0963_
rlabel metal2 8232 35448 8232 35448 0 _0964_
rlabel metal2 9464 37184 9464 37184 0 _0965_
rlabel metal3 10416 37352 10416 37352 0 _0966_
rlabel metal2 12600 53760 12600 53760 0 _0967_
rlabel metal2 12936 52584 12936 52584 0 _0968_
rlabel metal2 14784 54488 14784 54488 0 _0969_
rlabel metal3 20160 54320 20160 54320 0 _0970_
rlabel metal2 34328 55272 34328 55272 0 _0971_
rlabel metal3 20664 53648 20664 53648 0 _0972_
rlabel metal3 28840 54376 28840 54376 0 _0973_
rlabel metal2 32760 52416 32760 52416 0 _0974_
rlabel metal2 33712 56056 33712 56056 0 _0975_
rlabel metal3 35672 56728 35672 56728 0 _0976_
rlabel metal2 36120 53088 36120 53088 0 _0977_
rlabel metal2 36456 53424 36456 53424 0 _0978_
rlabel metal3 38836 56056 38836 56056 0 _0979_
rlabel metal2 42168 57232 42168 57232 0 _0980_
rlabel metal2 36008 56168 36008 56168 0 _0981_
rlabel metal2 36344 57344 36344 57344 0 _0982_
rlabel metal3 31136 55160 31136 55160 0 _0983_
rlabel metal2 24808 53816 24808 53816 0 _0984_
rlabel metal2 31752 55720 31752 55720 0 _0985_
rlabel metal2 32312 55776 32312 55776 0 _0986_
rlabel metal3 34104 56168 34104 56168 0 _0987_
rlabel metal2 11704 36960 11704 36960 0 _0988_
rlabel metal2 13328 47096 13328 47096 0 _0989_
rlabel metal2 15064 38920 15064 38920 0 _0990_
rlabel metal2 13664 46200 13664 46200 0 _0991_
rlabel metal3 13720 56168 13720 56168 0 _0992_
rlabel metal2 11256 56504 11256 56504 0 _0993_
rlabel metal3 12096 60760 12096 60760 0 _0994_
rlabel metal2 13944 56672 13944 56672 0 _0995_
rlabel metal3 14728 56056 14728 56056 0 _0996_
rlabel metal2 11144 54880 11144 54880 0 _0997_
rlabel metal2 11032 55384 11032 55384 0 _0998_
rlabel metal2 13496 55720 13496 55720 0 _0999_
rlabel metal2 14280 54768 14280 54768 0 _1000_
rlabel metal2 15288 55692 15288 55692 0 _1001_
rlabel metal2 27048 56728 27048 56728 0 _1002_
rlabel metal2 24976 41944 24976 41944 0 _1003_
rlabel metal2 25816 56840 25816 56840 0 _1004_
rlabel metal2 30576 38248 30576 38248 0 _1005_
rlabel metal2 26264 57232 26264 57232 0 _1006_
rlabel metal3 26992 56728 26992 56728 0 _1007_
rlabel metal2 27608 58072 27608 58072 0 _1008_
rlabel metal2 36008 58016 36008 58016 0 _1009_
rlabel metal2 39480 59024 39480 59024 0 _1010_
rlabel metal2 36232 59920 36232 59920 0 _1011_
rlabel metal2 36904 58912 36904 58912 0 _1012_
rlabel metal3 38808 62328 38808 62328 0 _1013_
rlabel metal2 25144 56952 25144 56952 0 _1014_
rlabel metal2 25760 57736 25760 57736 0 _1015_
rlabel metal2 25256 58128 25256 58128 0 _1016_
rlabel metal2 34776 61264 34776 61264 0 _1017_
rlabel metal2 31080 62216 31080 62216 0 _1018_
rlabel metal2 27888 60088 27888 60088 0 _1019_
rlabel metal2 27272 58520 27272 58520 0 _1020_
rlabel metal2 28392 60480 28392 60480 0 _1021_
rlabel metal2 25928 60704 25928 60704 0 _1022_
rlabel metal3 28448 59976 28448 59976 0 _1023_
rlabel metal3 28448 60760 28448 60760 0 _1024_
rlabel metal2 15456 44968 15456 44968 0 _1025_
rlabel metal2 12600 63448 12600 63448 0 _1026_
rlabel metal2 12040 43960 12040 43960 0 _1027_
rlabel metal2 10136 52640 10136 52640 0 _1028_
rlabel metal2 10304 52696 10304 52696 0 _1029_
rlabel metal2 12376 52864 12376 52864 0 _1030_
rlabel metal3 9632 49784 9632 49784 0 _1031_
rlabel metal2 3304 51296 3304 51296 0 _1032_
rlabel metal2 12544 52248 12544 52248 0 _1033_
rlabel metal2 14112 56616 14112 56616 0 _1034_
rlabel metal2 13720 56504 13720 56504 0 _1035_
rlabel metal2 15288 59080 15288 59080 0 _1036_
rlabel metal2 15736 60424 15736 60424 0 _1037_
rlabel metal2 34664 61264 34664 61264 0 _1038_
rlabel metal3 38920 62216 38920 62216 0 _1039_
rlabel metal2 41944 62664 41944 62664 0 _1040_
rlabel metal2 35672 61656 35672 61656 0 _1041_
rlabel metal2 35448 59696 35448 59696 0 _1042_
rlabel metal3 36456 61432 36456 61432 0 _1043_
rlabel metal2 34216 60256 34216 60256 0 _1044_
rlabel metal3 32872 59080 32872 59080 0 _1045_
rlabel metal2 31080 44296 31080 44296 0 _1046_
rlabel metal2 33096 60368 33096 60368 0 _1047_
rlabel metal2 15848 49896 15848 49896 0 _1048_
rlabel metal2 16576 43680 16576 43680 0 _1049_
rlabel metal2 16296 60368 16296 60368 0 _1050_
rlabel metal2 18144 60872 18144 60872 0 _1051_
rlabel metal2 16408 61992 16408 61992 0 _1052_
rlabel metal3 17864 59304 17864 59304 0 _1053_
rlabel metal2 16744 59976 16744 59976 0 _1054_
rlabel metal2 7896 62776 7896 62776 0 _1055_
rlabel metal2 13832 57064 13832 57064 0 _1056_
rlabel metal2 14168 58072 14168 58072 0 _1057_
rlabel metal2 17080 59920 17080 59920 0 _1058_
rlabel metal3 22260 60200 22260 60200 0 _1059_
rlabel metal2 34328 60648 34328 60648 0 _1060_
rlabel metal2 37408 62216 37408 62216 0 _1061_
rlabel metal2 45304 62664 45304 62664 0 _1062_
rlabel metal2 32536 63224 32536 63224 0 _1063_
rlabel metal2 20384 56840 20384 56840 0 _1064_
rlabel metal2 32536 60760 32536 60760 0 _1065_
rlabel metal2 32872 60704 32872 60704 0 _1066_
rlabel metal3 38892 60872 38892 60872 0 _1067_
rlabel metal2 17752 59976 17752 59976 0 _1068_
rlabel metal3 20160 59024 20160 59024 0 _1069_
rlabel metal2 38752 62328 38752 62328 0 _1070_
rlabel metal2 34776 60368 34776 60368 0 _1071_
rlabel metal2 38416 62216 38416 62216 0 _1072_
rlabel metal3 50568 62440 50568 62440 0 _1073_
rlabel metal3 39928 60872 39928 60872 0 _1074_
rlabel metal2 51632 57848 51632 57848 0 _1075_
rlabel metal2 52192 51352 52192 51352 0 _1076_
rlabel metal2 54264 51996 54264 51996 0 _1077_
rlabel metal3 51464 51128 51464 51128 0 _1078_
rlabel metal2 51688 53704 51688 53704 0 _1079_
rlabel metal3 30352 9576 30352 9576 0 _1080_
rlabel metal2 34664 25424 34664 25424 0 _1081_
rlabel metal2 33320 25928 33320 25928 0 _1082_
rlabel metal2 29512 25704 29512 25704 0 _1083_
rlabel metal2 26936 25816 26936 25816 0 _1084_
rlabel metal2 27944 24472 27944 24472 0 _1085_
rlabel metal2 29176 24640 29176 24640 0 _1086_
rlabel metal2 32984 22428 32984 22428 0 _1087_
rlabel metal2 30968 5824 30968 5824 0 _1088_
rlabel metal2 31528 10136 31528 10136 0 _1089_
rlabel metal2 30744 10136 30744 10136 0 _1090_
rlabel metal2 35784 24584 35784 24584 0 _1091_
rlabel metal3 24416 29624 24416 29624 0 _1092_
rlabel metal2 46480 6776 46480 6776 0 _1093_
rlabel metal2 36008 17080 36008 17080 0 _1094_
rlabel metal2 33768 19320 33768 19320 0 _1095_
rlabel metal3 45304 8232 45304 8232 0 _1096_
rlabel metal3 24696 19208 24696 19208 0 _1097_
rlabel metal3 35000 18144 35000 18144 0 _1098_
rlabel metal2 45864 7728 45864 7728 0 _1099_
rlabel metal3 31416 8008 31416 8008 0 _1100_
rlabel metal2 14168 25200 14168 25200 0 _1101_
rlabel metal2 44968 5432 44968 5432 0 _1102_
rlabel metal2 30744 5432 30744 5432 0 _1103_
rlabel metal2 14224 24808 14224 24808 0 _1104_
rlabel metal2 44128 6664 44128 6664 0 _1105_
rlabel metal2 31640 6104 31640 6104 0 _1106_
rlabel metal3 47880 4536 47880 4536 0 _1107_
rlabel metal3 39928 25368 39928 25368 0 _1108_
rlabel metal3 40320 26264 40320 26264 0 _1109_
rlabel metal3 41720 9240 41720 9240 0 _1110_
rlabel metal3 45920 5880 45920 5880 0 _1111_
rlabel metal2 46200 7840 46200 7840 0 _1112_
rlabel metal3 46816 5992 46816 5992 0 _1113_
rlabel metal2 46088 8232 46088 8232 0 _1114_
rlabel metal3 45976 5096 45976 5096 0 _1115_
rlabel metal2 45864 4872 45864 4872 0 _1116_
rlabel metal2 43736 7112 43736 7112 0 _1117_
rlabel metal3 48328 21784 48328 21784 0 _1118_
rlabel metal2 39816 25872 39816 25872 0 _1119_
rlabel metal2 44632 23688 44632 23688 0 _1120_
rlabel metal2 45640 22792 45640 22792 0 _1121_
rlabel metal2 47544 19880 47544 19880 0 _1122_
rlabel metal2 47096 22008 47096 22008 0 _1123_
rlabel metal2 47096 18872 47096 18872 0 _1124_
rlabel metal2 46200 19320 46200 19320 0 _1125_
rlabel metal2 21336 38136 21336 38136 0 _1126_
rlabel metal2 22008 48720 22008 48720 0 _1127_
rlabel metal2 46480 22344 46480 22344 0 _1128_
rlabel metal2 41384 40488 41384 40488 0 _1129_
rlabel metal3 49672 45752 49672 45752 0 _1130_
rlabel metal2 49000 39312 49000 39312 0 _1131_
rlabel metal3 25032 12936 25032 12936 0 _1132_
rlabel metal3 39984 38584 39984 38584 0 _1133_
rlabel metal2 40880 36680 40880 36680 0 _1134_
rlabel metal2 39144 37688 39144 37688 0 _1135_
rlabel metal2 39984 37464 39984 37464 0 _1136_
rlabel metal2 23688 44016 23688 44016 0 _1137_
rlabel metal2 22288 44184 22288 44184 0 _1138_
rlabel metal2 22792 43848 22792 43848 0 _1139_
rlabel metal3 49560 46648 49560 46648 0 _1140_
rlabel metal2 25480 47096 25480 47096 0 _1141_
rlabel metal2 23912 49784 23912 49784 0 _1142_
rlabel metal2 22008 45024 22008 45024 0 _1143_
rlabel metal2 23352 45192 23352 45192 0 _1144_
rlabel metal2 22904 46760 22904 46760 0 _1145_
rlabel metal2 22120 49000 22120 49000 0 _1146_
rlabel metal2 24360 47768 24360 47768 0 _1147_
rlabel metal3 24136 47432 24136 47432 0 _1148_
rlabel metal2 21560 48216 21560 48216 0 _1149_
rlabel metal2 20216 49112 20216 49112 0 _1150_
rlabel metal2 20440 48552 20440 48552 0 _1151_
rlabel metal3 21000 48888 21000 48888 0 _1152_
rlabel metal3 20496 49784 20496 49784 0 _1153_
rlabel metal2 21224 49672 21224 49672 0 _1154_
rlabel metal2 20328 50960 20328 50960 0 _1155_
rlabel metal2 18592 53480 18592 53480 0 _1156_
rlabel metal3 17080 54488 17080 54488 0 _1157_
rlabel metal2 17864 53760 17864 53760 0 _1158_
rlabel metal2 20216 52864 20216 52864 0 _1159_
rlabel metal2 20440 53032 20440 53032 0 _1160_
rlabel metal2 23128 52528 23128 52528 0 _1161_
rlabel metal2 22568 52752 22568 52752 0 _1162_
rlabel metal2 23912 53256 23912 53256 0 _1163_
rlabel metal2 24024 53424 24024 53424 0 _1164_
rlabel metal2 23016 56112 23016 56112 0 _1165_
rlabel metal2 22680 56840 22680 56840 0 _1166_
rlabel metal2 23800 56448 23800 56448 0 _1167_
rlabel metal2 24696 57344 24696 57344 0 _1168_
rlabel metal2 24024 59920 24024 59920 0 _1169_
rlabel metal2 23184 59864 23184 59864 0 _1170_
rlabel metal2 2968 46032 2968 46032 0 _1171_
rlabel metal2 25480 61152 25480 61152 0 _1172_
rlabel metal2 26264 60368 26264 60368 0 _1173_
rlabel metal2 25928 60088 25928 60088 0 _1174_
rlabel metal2 20776 57680 20776 57680 0 _1175_
rlabel metal2 18480 55944 18480 55944 0 _1176_
rlabel metal3 19880 57624 19880 57624 0 _1177_
rlabel metal2 20104 57288 20104 57288 0 _1178_
rlabel metal2 2744 37408 2744 37408 0 _1179_
rlabel metal3 3472 37240 3472 37240 0 _1180_
rlabel metal2 3080 40432 3080 40432 0 _1181_
rlabel metal2 2856 40600 2856 40600 0 _1182_
rlabel metal2 4984 40768 4984 40768 0 _1183_
rlabel metal3 5376 41160 5376 41160 0 _1184_
rlabel metal2 3640 41888 3640 41888 0 _1185_
rlabel metal2 4536 44352 4536 44352 0 _1186_
rlabel metal2 5096 44072 5096 44072 0 _1187_
rlabel metal2 3528 44464 3528 44464 0 _1188_
rlabel metal2 2912 42840 2912 42840 0 _1189_
rlabel metal2 4984 44016 4984 44016 0 _1190_
rlabel metal2 4088 45528 4088 45528 0 _1191_
rlabel metal3 3080 46536 3080 46536 0 _1192_
rlabel metal2 5656 47880 5656 47880 0 _1193_
rlabel metal2 5712 48328 5712 48328 0 _1194_
rlabel metal2 4760 49672 4760 49672 0 _1195_
rlabel metal2 5096 51072 5096 51072 0 _1196_
rlabel metal2 4312 50064 4312 50064 0 _1197_
rlabel metal2 4872 50092 4872 50092 0 _1198_
rlabel metal3 4648 50568 4648 50568 0 _1199_
rlabel metal2 5768 51072 5768 51072 0 _1200_
rlabel metal2 3192 54880 3192 54880 0 _1201_
rlabel metal2 2856 55104 2856 55104 0 _1202_
rlabel metal2 6776 39704 6776 39704 0 _1203_
rlabel metal2 3640 55272 3640 55272 0 _1204_
rlabel metal2 4648 53816 4648 53816 0 _1205_
rlabel metal2 5096 54936 5096 54936 0 _1206_
rlabel metal3 4312 56840 4312 56840 0 _1207_
rlabel metal3 4424 57736 4424 57736 0 _1208_
rlabel metal2 4368 56952 4368 56952 0 _1209_
rlabel metal3 21112 45640 21112 45640 0 _1210_
rlabel metal3 20216 47040 20216 47040 0 _1211_
rlabel metal2 6328 57904 6328 57904 0 _1212_
rlabel metal2 6104 57176 6104 57176 0 _1213_
rlabel metal2 7112 59864 7112 59864 0 _1214_
rlabel metal2 7840 59304 7840 59304 0 _1215_
rlabel metal2 6552 60536 6552 60536 0 _1216_
rlabel metal2 7448 60648 7448 60648 0 _1217_
rlabel metal3 6944 62328 6944 62328 0 _1218_
rlabel metal2 8008 62384 8008 62384 0 _1219_
rlabel metal3 7112 63000 7112 63000 0 _1220_
rlabel metal2 7224 62776 7224 62776 0 _1221_
rlabel metal2 8344 62328 8344 62328 0 _1222_
rlabel metal2 9128 62328 9128 62328 0 _1223_
rlabel metal3 14952 62440 14952 62440 0 _1224_
rlabel metal2 18984 60816 18984 60816 0 _1225_
rlabel metal2 19432 62832 19432 62832 0 _1226_
rlabel metal2 43736 12992 43736 12992 0 _1227_
rlabel metal2 29960 25032 29960 25032 0 _1228_
rlabel metal2 19824 62552 19824 62552 0 _1229_
rlabel metal2 7896 38976 7896 38976 0 _1230_
rlabel metal2 6496 38024 6496 38024 0 _1231_
rlabel metal3 9408 41160 9408 41160 0 _1232_
rlabel metal2 8344 41776 8344 41776 0 _1233_
rlabel metal2 8904 42112 8904 42112 0 _1234_
rlabel metal2 9912 42056 9912 42056 0 _1235_
rlabel metal2 10136 44016 10136 44016 0 _1236_
rlabel metal2 8064 44408 8064 44408 0 _1237_
rlabel metal2 8400 45640 8400 45640 0 _1238_
rlabel metal2 7784 45080 7784 45080 0 _1239_
rlabel metal2 9128 46312 9128 46312 0 _1240_
rlabel metal2 9632 45304 9632 45304 0 _1241_
rlabel metal3 10416 47432 10416 47432 0 _1242_
rlabel metal2 12488 47880 12488 47880 0 _1243_
rlabel metal2 11256 48160 11256 48160 0 _1244_
rlabel metal2 12600 46984 12600 46984 0 _1245_
rlabel metal2 9576 48272 9576 48272 0 _1246_
rlabel metal2 8680 49616 8680 49616 0 _1247_
rlabel metal2 8568 48720 8568 48720 0 _1248_
rlabel metal2 8456 48608 8456 48608 0 _1249_
rlabel metal2 9912 49784 9912 49784 0 _1250_
rlabel metal2 9464 50064 9464 50064 0 _1251_
rlabel metal2 8624 52920 8624 52920 0 _1252_
rlabel metal2 7336 52528 7336 52528 0 _1253_
rlabel metal3 8120 53144 8120 53144 0 _1254_
rlabel metal2 8792 52752 8792 52752 0 _1255_
rlabel metal2 8680 53704 8680 53704 0 _1256_
rlabel metal2 8568 54992 8568 54992 0 _1257_
rlabel metal3 8512 56280 8512 56280 0 _1258_
rlabel metal2 29680 26152 29680 26152 0 clknet_0_wb_clk_i
rlabel metal2 14392 10192 14392 10192 0 clknet_4_0_0_wb_clk_i
rlabel metal2 2856 60424 2856 60424 0 clknet_4_10_0_wb_clk_i
rlabel metal2 20664 53088 20664 53088 0 clknet_4_11_0_wb_clk_i
rlabel metal2 44856 47488 44856 47488 0 clknet_4_12_0_wb_clk_i
rlabel metal2 49672 49336 49672 49336 0 clknet_4_13_0_wb_clk_i
rlabel metal2 44408 65408 44408 65408 0 clknet_4_14_0_wb_clk_i
rlabel metal2 55272 53424 55272 53424 0 clknet_4_15_0_wb_clk_i
rlabel metal2 30856 20776 30856 20776 0 clknet_4_1_0_wb_clk_i
rlabel metal2 10136 24976 10136 24976 0 clknet_4_2_0_wb_clk_i
rlabel metal2 30744 23240 30744 23240 0 clknet_4_3_0_wb_clk_i
rlabel metal2 44072 5544 44072 5544 0 clknet_4_4_0_wb_clk_i
rlabel metal3 48720 5096 48720 5096 0 clknet_4_5_0_wb_clk_i
rlabel metal2 38472 24360 38472 24360 0 clknet_4_6_0_wb_clk_i
rlabel metal2 47992 22736 47992 22736 0 clknet_4_7_0_wb_clk_i
rlabel metal2 1848 49000 1848 49000 0 clknet_4_8_0_wb_clk_i
rlabel metal3 22792 49000 22792 49000 0 clknet_4_9_0_wb_clk_i
rlabel metal3 58730 59192 58730 59192 0 custom_settings[0]
rlabel metal2 58184 65800 58184 65800 0 custom_settings[1]
rlabel metal2 58184 3976 58184 3976 0 io_in_1[0]
rlabel metal3 58730 10584 58730 10584 0 io_in_1[1]
rlabel metal3 58730 17528 58730 17528 0 io_in_1[2]
rlabel metal2 58184 24920 58184 24920 0 io_in_1[3]
rlabel metal2 58184 31248 58184 31248 0 io_in_1[4]
rlabel metal3 57848 38808 57848 38808 0 io_in_1[5]
rlabel metal3 58730 45304 58730 45304 0 io_in_1[6]
rlabel metal2 58184 52584 58184 52584 0 io_in_1[7]
rlabel metal3 1246 58296 1246 58296 0 io_in_2
rlabel metal2 22904 67802 22904 67802 0 io_out[10]
rlabel metal3 25536 66472 25536 66472 0 io_out[11]
rlabel metal2 26936 68222 26936 68222 0 io_out[12]
rlabel metal2 37016 67802 37016 67802 0 io_out[17]
rlabel metal3 39928 66472 39928 66472 0 io_out[18]
rlabel metal3 41888 65464 41888 65464 0 io_out[19]
rlabel metal2 43848 66808 43848 66808 0 io_out[20]
rlabel metal3 46760 66472 46760 66472 0 io_out[21]
rlabel metal2 47096 68222 47096 68222 0 io_out[22]
rlabel metal3 50680 66472 50680 66472 0 io_out[23]
rlabel metal3 51128 65520 51128 65520 0 io_out[24]
rlabel metal2 53144 67858 53144 67858 0 io_out[25]
rlabel metal2 55160 66514 55160 66514 0 io_out[26]
rlabel metal2 55384 63672 55384 63672 0 io_out[27]
rlabel metal2 18872 67802 18872 67802 0 io_out[8]
rlabel metal2 20888 68222 20888 68222 0 io_out[9]
rlabel metal2 57792 59080 57792 59080 0 net1
rlabel metal3 29288 26264 29288 26264 0 net10
rlabel metal2 2296 29204 2296 29204 0 net11
rlabel metal3 49336 47208 49336 47208 0 net12
rlabel metal2 23016 64624 23016 64624 0 net13
rlabel metal2 24696 65800 24696 65800 0 net14
rlabel metal2 30296 65128 30296 65128 0 net15
rlabel metal2 39424 63896 39424 63896 0 net16
rlabel metal2 39592 65800 39592 65800 0 net17
rlabel metal2 41384 64736 41384 64736 0 net18
rlabel metal2 46200 64848 46200 64848 0 net19
rlabel metal2 57680 60984 57680 60984 0 net2
rlabel metal2 47432 64204 47432 64204 0 net20
rlabel metal2 49448 63504 49448 63504 0 net21
rlabel metal2 51016 63056 51016 63056 0 net22
rlabel metal3 50456 63896 50456 63896 0 net23
rlabel metal2 50680 63280 50680 63280 0 net24
rlabel metal2 52808 61152 52808 61152 0 net25
rlabel metal2 54712 60648 54712 60648 0 net26
rlabel metal2 17416 65800 17416 65800 0 net27
rlabel metal2 20776 64400 20776 64400 0 net28
rlabel metal2 2744 68222 2744 68222 0 net29
rlabel metal2 31640 23184 31640 23184 0 net3
rlabel metal2 5544 66472 5544 66472 0 net30
rlabel metal2 6776 68222 6776 68222 0 net31
rlabel metal2 9352 66472 9352 66472 0 net32
rlabel metal2 10808 68222 10808 68222 0 net33
rlabel metal2 12824 68222 12824 68222 0 net34
rlabel metal2 14840 68222 14840 68222 0 net35
rlabel metal2 16856 68222 16856 68222 0 net36
rlabel metal2 28952 68222 28952 68222 0 net37
rlabel metal2 30968 68222 30968 68222 0 net38
rlabel metal2 32984 68222 32984 68222 0 net39
rlabel metal2 57624 11256 57624 11256 0 net4
rlabel metal2 35000 68222 35000 68222 0 net40
rlabel metal2 34440 26656 34440 26656 0 net5
rlabel metal2 57848 25032 57848 25032 0 net6
rlabel metal2 40152 26208 40152 26208 0 net7
rlabel metal2 36232 25648 36232 25648 0 net8
rlabel metal3 31360 26488 31360 26488 0 net9
rlabel metal3 1302 35000 1302 35000 0 rst_n
rlabel metal2 18648 32088 18648 32088 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
rlabel metal2 19208 25984 19208 25984 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
rlabel metal2 19992 35280 19992 35280 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
rlabel metal2 13944 23856 13944 23856 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
rlabel metal3 18256 34776 18256 34776 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.in
rlabel metal2 7672 30128 7672 30128 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
rlabel metal3 8624 27720 8624 27720 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
rlabel metal2 11816 25928 11816 25928 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
rlabel metal2 12936 26208 12936 26208 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
rlabel metal2 8904 26488 8904 26488 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.in
rlabel metal2 24136 32984 24136 32984 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
rlabel metal2 24024 35336 24024 35336 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
rlabel metal3 24080 37128 24080 37128 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
rlabel metal2 22736 40488 22736 40488 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
rlabel metal2 25480 34776 25480 34776 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.in
rlabel metal2 34440 27776 34440 27776 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
rlabel metal2 31864 32592 31864 32592 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
rlabel metal2 36568 35112 36568 35112 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
rlabel metal2 38360 34776 38360 34776 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
rlabel metal2 37576 31808 37576 31808 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.in
rlabel metal2 57008 39592 57008 39592 0 tt_um_rejunity_sn76489.clk_counter\[0\]
rlabel metal2 56728 43456 56728 43456 0 tt_um_rejunity_sn76489.clk_counter\[1\]
rlabel metal2 55440 45080 55440 45080 0 tt_um_rejunity_sn76489.clk_counter\[2\]
rlabel metal2 55944 42280 55944 42280 0 tt_um_rejunity_sn76489.clk_counter\[3\]
rlabel metal2 51912 44632 51912 44632 0 tt_um_rejunity_sn76489.clk_counter\[4\]
rlabel metal2 52024 42168 52024 42168 0 tt_um_rejunity_sn76489.clk_counter\[5\]
rlabel metal2 53144 39928 53144 39928 0 tt_um_rejunity_sn76489.clk_counter\[6\]
rlabel metal2 38416 25256 38416 25256 0 tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
rlabel metal2 39872 30296 39872 30296 0 tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
rlabel metal2 41496 29008 41496 29008 0 tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
rlabel metal3 29288 9688 29288 9688 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
rlabel metal3 29736 7336 29736 7336 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
rlabel metal3 25956 6552 25956 6552 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
rlabel metal2 29400 5376 29400 5376 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
rlabel metal3 19096 16184 19096 16184 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
rlabel metal2 16856 16912 16856 16912 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
rlabel metal2 18704 19992 18704 19992 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
rlabel metal3 17920 18984 17920 18984 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
rlabel metal2 22792 16800 22792 16800 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
rlabel metal2 22400 19880 22400 19880 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
rlabel metal2 49896 6048 49896 6048 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
rlabel metal3 47040 8232 47040 8232 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
rlabel metal3 47824 4200 47824 4200 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
rlabel metal3 40992 7560 40992 7560 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
rlabel metal2 29512 15512 29512 15512 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
rlabel metal2 30072 13720 30072 13720 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
rlabel metal2 30240 18984 30240 18984 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
rlabel metal2 28728 17864 28728 17864 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
rlabel metal2 31752 16856 31752 16856 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
rlabel metal2 33656 18200 33656 18200 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
rlabel metal2 50848 22456 50848 22456 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
rlabel metal2 50008 18480 50008 18480 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
rlabel metal2 47768 19656 47768 19656 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
rlabel metal2 48216 22736 48216 22736 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
rlabel metal2 44184 19600 44184 19600 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
rlabel metal2 46816 15064 46816 15064 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
rlabel metal2 44296 17808 44296 17808 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
rlabel metal2 40712 16520 40712 16520 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
rlabel metal2 38136 16856 38136 16856 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
rlabel metal2 36456 22792 36456 22792 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
rlabel metal3 7224 38584 7224 38584 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
rlabel metal2 9688 41552 9688 41552 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
rlabel metal2 8904 45864 8904 45864 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
rlabel metal2 10584 47152 10584 47152 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
rlabel metal2 8904 48720 8904 48720 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
rlabel metal2 8176 52808 8176 52808 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
rlabel metal2 10248 57848 10248 57848 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
rlabel metal2 11256 60032 11256 60032 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
rlabel metal2 12936 63952 12936 63952 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
rlabel metal2 16408 63896 16408 63896 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
rlabel metal2 3864 36904 3864 36904 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
rlabel metal2 5096 40768 5096 40768 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
rlabel metal2 4928 45192 4928 45192 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
rlabel metal2 5768 47432 5768 47432 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
rlabel metal2 4984 50624 4984 50624 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
rlabel metal2 4648 54432 4648 54432 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
rlabel metal2 5656 57232 5656 57232 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
rlabel metal2 6328 60760 6328 60760 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
rlabel metal2 8904 64792 8904 64792 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
rlabel metal2 20216 60144 20216 60144 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
rlabel metal3 41384 40376 41384 40376 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
rlabel metal2 39704 37240 39704 37240 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
rlabel metal2 21784 45136 21784 45136 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
rlabel metal2 24472 48776 24472 48776 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
rlabel metal2 19600 49112 19600 49112 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
rlabel metal2 20328 52528 20328 52528 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
rlabel metal3 23744 53592 23744 53592 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
rlabel metal2 24248 56560 24248 56560 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
rlabel metal2 24920 60648 24920 60648 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
rlabel metal2 20216 56392 20216 56392 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
rlabel metal2 45808 38024 45808 38024 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
rlabel metal2 47544 39984 47544 39984 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
rlabel metal2 32424 44632 32424 44632 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
rlabel metal2 29848 46368 29848 46368 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
rlabel metal2 28392 51044 28392 51044 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
rlabel metal2 28952 54096 28952 54096 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
rlabel metal2 30632 57736 30632 57736 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
rlabel metal2 27496 64344 27496 64344 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
rlabel metal2 31304 63056 31304 63056 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
rlabel metal2 33544 64344 33544 64344 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
rlabel metal2 22680 24640 22680 24640 0 tt_um_rejunity_sn76489.latch_control_reg\[0\]
rlabel metal3 25200 22344 25200 22344 0 tt_um_rejunity_sn76489.latch_control_reg\[1\]
rlabel metal2 27664 24808 27664 24808 0 tt_um_rejunity_sn76489.latch_control_reg\[2\]
rlabel metal2 45136 25368 45136 25368 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
rlabel metal2 45304 25760 45304 25760 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
rlabel metal3 43736 28392 43736 28392 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
rlabel metal3 44744 31752 44744 31752 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
rlabel metal2 41272 33712 41272 33712 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
rlabel metal2 42728 35000 42728 35000 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
rlabel metal2 45976 33600 45976 33600 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
rlabel metal3 57848 33096 57848 33096 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
rlabel metal2 57848 37016 57848 37016 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
rlabel metal2 56672 35896 56672 35896 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
rlabel metal2 55608 33096 55608 33096 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
rlabel metal2 51240 33096 51240 33096 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
rlabel metal2 50344 30184 50344 30184 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
rlabel metal2 54264 27328 54264 27328 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
rlabel metal2 52528 26376 52528 26376 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
rlabel metal3 53704 23744 53704 23744 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
rlabel metal3 53200 23240 53200 23240 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
rlabel metal2 57848 21504 57848 21504 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
rlabel metal3 55944 23352 55944 23352 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
rlabel metal2 56616 25480 56616 25480 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
rlabel metal3 57568 29624 57568 29624 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
rlabel metal3 49168 28728 49168 28728 0 tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
rlabel metal2 52080 35784 52080 35784 0 tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
rlabel metal3 47544 43400 47544 43400 0 tt_um_rejunity_sn76489.pwm.accumulator\[0\]
rlabel metal3 54600 63224 54600 63224 0 tt_um_rejunity_sn76489.pwm.accumulator\[10\]
rlabel metal2 55272 60536 55272 60536 0 tt_um_rejunity_sn76489.pwm.accumulator\[11\]
rlabel metal2 44072 44296 44072 44296 0 tt_um_rejunity_sn76489.pwm.accumulator\[1\]
rlabel metal2 44856 46928 44856 46928 0 tt_um_rejunity_sn76489.pwm.accumulator\[2\]
rlabel metal2 42616 47712 42616 47712 0 tt_um_rejunity_sn76489.pwm.accumulator\[3\]
rlabel metal3 38136 49896 38136 49896 0 tt_um_rejunity_sn76489.pwm.accumulator\[4\]
rlabel metal2 41496 55160 41496 55160 0 tt_um_rejunity_sn76489.pwm.accumulator\[5\]
rlabel metal2 43176 58352 43176 58352 0 tt_um_rejunity_sn76489.pwm.accumulator\[6\]
rlabel metal2 41384 59640 41384 59640 0 tt_um_rejunity_sn76489.pwm.accumulator\[7\]
rlabel metal3 44632 63000 44632 63000 0 tt_um_rejunity_sn76489.pwm.accumulator\[8\]
rlabel via2 46536 64232 46536 64232 0 tt_um_rejunity_sn76489.pwm.accumulator\[9\]
rlabel metal2 53704 53144 53704 53144 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
rlabel metal2 55384 51296 55384 51296 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
rlabel metal2 57064 51464 57064 51464 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
rlabel metal2 55160 54264 55160 54264 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
rlabel metal2 54936 53984 54936 53984 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
rlabel metal2 46816 49112 46816 49112 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 54264 59528 54264 59528 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 53984 52920 53984 52920 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 46928 51352 46928 51352 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 47712 52248 47712 52248 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 46648 53816 46648 53816 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 47768 54880 47768 54880 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 48104 56728 48104 56728 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 49896 59640 49896 59640 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal3 50904 62216 50904 62216 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 50792 63896 50792 63896 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 51800 61544 51800 61544 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 24696 9464 24696 9464 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
rlabel metal2 25928 6944 25928 6944 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
rlabel metal2 24472 5432 24472 5432 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
rlabel metal2 22344 6552 22344 6552 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
rlabel metal2 18760 7728 18760 7728 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
rlabel metal3 17752 9688 17752 9688 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
rlabel metal2 18760 11088 18760 11088 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
rlabel metal3 17808 13832 17808 13832 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
rlabel metal2 21672 10416 21672 10416 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
rlabel metal2 23296 15960 23296 15960 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
rlabel metal3 51408 8232 51408 8232 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
rlabel metal2 51464 7112 51464 7112 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
rlabel metal2 51240 6496 51240 6496 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
rlabel metal2 48328 7112 48328 7112 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
rlabel metal2 37128 9464 37128 9464 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
rlabel metal2 35112 5824 35112 5824 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
rlabel metal2 34664 6328 34664 6328 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
rlabel metal2 33320 11592 33320 11592 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
rlabel metal2 38136 11984 38136 11984 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
rlabel metal2 37856 15176 37856 15176 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
rlabel metal2 52136 13272 52136 13272 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
rlabel metal2 53144 18088 53144 18088 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
rlabel metal3 52248 17528 52248 17528 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
rlabel metal2 53592 14784 53592 14784 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
rlabel metal3 52584 14504 52584 14504 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
rlabel metal2 46984 12936 46984 12936 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
rlabel metal2 45976 12936 45976 12936 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
rlabel metal2 42840 14784 42840 14784 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
rlabel metal3 46620 12488 46620 12488 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
rlabel metal4 40712 19208 40712 19208 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
rlabel metal3 1862 11704 1862 11704 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 60000 70000
<< end >>
