VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_pdp11
  CLASS BLOCK ;
  FOREIGN wrapped_pdp11 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 800.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 452.480 4.000 453.040 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 488.320 4.000 488.880 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 667.520 4.000 668.080 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 703.360 4.000 703.920 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 739.200 4.000 739.760 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 775.040 4.000 775.600 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.920 4.000 130.480 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.440 4.000 238.000 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.960 4.000 345.520 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END custom_settings[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 0.000 295.120 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 0.000 456.400 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 0.000 483.280 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 0.000 563.920 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 0.000 617.680 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 644.000 0.000 644.560 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 697.760 0.000 698.320 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 724.640 0.000 725.200 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 778.400 0.000 778.960 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 805.280 0.000 805.840 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 859.040 0.000 859.600 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 885.920 0.000 886.480 4.000 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 22.400 1800.000 22.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 257.600 1800.000 258.160 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 281.120 1800.000 281.680 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 304.640 1800.000 305.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 328.160 1800.000 328.720 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 351.680 1800.000 352.240 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 375.200 1800.000 375.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 398.720 1800.000 399.280 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 422.240 1800.000 422.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 445.760 1800.000 446.320 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 469.280 1800.000 469.840 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 45.920 1800.000 46.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 492.800 1800.000 493.360 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 516.320 1800.000 516.880 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 539.840 1800.000 540.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 563.360 1800.000 563.920 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 586.880 1800.000 587.440 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 610.400 1800.000 610.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 633.920 1800.000 634.480 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 657.440 1800.000 658.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 680.960 1800.000 681.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 704.480 1800.000 705.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 69.440 1800.000 70.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 728.000 1800.000 728.560 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 751.520 1800.000 752.080 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 775.040 1800.000 775.600 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 92.960 1800.000 93.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 116.480 1800.000 117.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 140.000 1800.000 140.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 163.520 1800.000 164.080 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 187.040 1800.000 187.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 210.560 1800.000 211.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1796.000 234.080 1800.000 234.640 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 912.800 0.000 913.360 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1181.600 0.000 1182.160 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1208.480 0.000 1209.040 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1235.360 0.000 1235.920 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1262.240 0.000 1262.800 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1289.120 0.000 1289.680 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1316.000 0.000 1316.560 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1342.880 0.000 1343.440 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1369.760 0.000 1370.320 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1396.640 0.000 1397.200 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 1423.520 0.000 1424.080 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 0.000 940.240 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1450.400 0.000 1450.960 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1477.280 0.000 1477.840 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1504.160 0.000 1504.720 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1531.040 0.000 1531.600 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1557.920 0.000 1558.480 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1584.800 0.000 1585.360 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1611.680 0.000 1612.240 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1638.560 0.000 1639.120 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1665.440 0.000 1666.000 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1692.320 0.000 1692.880 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 966.560 0.000 967.120 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1719.200 0.000 1719.760 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1746.080 0.000 1746.640 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1772.960 0.000 1773.520 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 993.440 0.000 994.000 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1020.320 0.000 1020.880 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1047.200 0.000 1047.760 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1074.080 0.000 1074.640 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1100.960 0.000 1101.520 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1127.840 0.000 1128.400 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1154.720 0.000 1155.280 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 4.000 58.800 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 4.000 22.960 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1793.120 784.300 ;
      LAYER Metal2 ;
        RECT 5.740 4.300 1790.740 793.430 ;
        RECT 5.740 3.450 25.460 4.300 ;
        RECT 26.620 3.450 52.340 4.300 ;
        RECT 53.500 3.450 79.220 4.300 ;
        RECT 80.380 3.450 106.100 4.300 ;
        RECT 107.260 3.450 132.980 4.300 ;
        RECT 134.140 3.450 159.860 4.300 ;
        RECT 161.020 3.450 186.740 4.300 ;
        RECT 187.900 3.450 213.620 4.300 ;
        RECT 214.780 3.450 240.500 4.300 ;
        RECT 241.660 3.450 267.380 4.300 ;
        RECT 268.540 3.450 294.260 4.300 ;
        RECT 295.420 3.450 321.140 4.300 ;
        RECT 322.300 3.450 348.020 4.300 ;
        RECT 349.180 3.450 374.900 4.300 ;
        RECT 376.060 3.450 401.780 4.300 ;
        RECT 402.940 3.450 428.660 4.300 ;
        RECT 429.820 3.450 455.540 4.300 ;
        RECT 456.700 3.450 482.420 4.300 ;
        RECT 483.580 3.450 509.300 4.300 ;
        RECT 510.460 3.450 536.180 4.300 ;
        RECT 537.340 3.450 563.060 4.300 ;
        RECT 564.220 3.450 589.940 4.300 ;
        RECT 591.100 3.450 616.820 4.300 ;
        RECT 617.980 3.450 643.700 4.300 ;
        RECT 644.860 3.450 670.580 4.300 ;
        RECT 671.740 3.450 697.460 4.300 ;
        RECT 698.620 3.450 724.340 4.300 ;
        RECT 725.500 3.450 751.220 4.300 ;
        RECT 752.380 3.450 778.100 4.300 ;
        RECT 779.260 3.450 804.980 4.300 ;
        RECT 806.140 3.450 831.860 4.300 ;
        RECT 833.020 3.450 858.740 4.300 ;
        RECT 859.900 3.450 885.620 4.300 ;
        RECT 886.780 3.450 912.500 4.300 ;
        RECT 913.660 3.450 939.380 4.300 ;
        RECT 940.540 3.450 966.260 4.300 ;
        RECT 967.420 3.450 993.140 4.300 ;
        RECT 994.300 3.450 1020.020 4.300 ;
        RECT 1021.180 3.450 1046.900 4.300 ;
        RECT 1048.060 3.450 1073.780 4.300 ;
        RECT 1074.940 3.450 1100.660 4.300 ;
        RECT 1101.820 3.450 1127.540 4.300 ;
        RECT 1128.700 3.450 1154.420 4.300 ;
        RECT 1155.580 3.450 1181.300 4.300 ;
        RECT 1182.460 3.450 1208.180 4.300 ;
        RECT 1209.340 3.450 1235.060 4.300 ;
        RECT 1236.220 3.450 1261.940 4.300 ;
        RECT 1263.100 3.450 1288.820 4.300 ;
        RECT 1289.980 3.450 1315.700 4.300 ;
        RECT 1316.860 3.450 1342.580 4.300 ;
        RECT 1343.740 3.450 1369.460 4.300 ;
        RECT 1370.620 3.450 1396.340 4.300 ;
        RECT 1397.500 3.450 1423.220 4.300 ;
        RECT 1424.380 3.450 1450.100 4.300 ;
        RECT 1451.260 3.450 1476.980 4.300 ;
        RECT 1478.140 3.450 1503.860 4.300 ;
        RECT 1505.020 3.450 1530.740 4.300 ;
        RECT 1531.900 3.450 1557.620 4.300 ;
        RECT 1558.780 3.450 1584.500 4.300 ;
        RECT 1585.660 3.450 1611.380 4.300 ;
        RECT 1612.540 3.450 1638.260 4.300 ;
        RECT 1639.420 3.450 1665.140 4.300 ;
        RECT 1666.300 3.450 1692.020 4.300 ;
        RECT 1693.180 3.450 1718.900 4.300 ;
        RECT 1720.060 3.450 1745.780 4.300 ;
        RECT 1746.940 3.450 1772.660 4.300 ;
        RECT 1773.820 3.450 1790.740 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 775.900 1796.340 793.380 ;
        RECT 4.300 774.740 1795.700 775.900 ;
        RECT 4.000 752.380 1796.340 774.740 ;
        RECT 4.000 751.220 1795.700 752.380 ;
        RECT 4.000 740.060 1796.340 751.220 ;
        RECT 4.300 738.900 1796.340 740.060 ;
        RECT 4.000 728.860 1796.340 738.900 ;
        RECT 4.000 727.700 1795.700 728.860 ;
        RECT 4.000 705.340 1796.340 727.700 ;
        RECT 4.000 704.220 1795.700 705.340 ;
        RECT 4.300 704.180 1795.700 704.220 ;
        RECT 4.300 703.060 1796.340 704.180 ;
        RECT 4.000 681.820 1796.340 703.060 ;
        RECT 4.000 680.660 1795.700 681.820 ;
        RECT 4.000 668.380 1796.340 680.660 ;
        RECT 4.300 667.220 1796.340 668.380 ;
        RECT 4.000 658.300 1796.340 667.220 ;
        RECT 4.000 657.140 1795.700 658.300 ;
        RECT 4.000 634.780 1796.340 657.140 ;
        RECT 4.000 633.620 1795.700 634.780 ;
        RECT 4.000 632.540 1796.340 633.620 ;
        RECT 4.300 631.380 1796.340 632.540 ;
        RECT 4.000 611.260 1796.340 631.380 ;
        RECT 4.000 610.100 1795.700 611.260 ;
        RECT 4.000 596.700 1796.340 610.100 ;
        RECT 4.300 595.540 1796.340 596.700 ;
        RECT 4.000 587.740 1796.340 595.540 ;
        RECT 4.000 586.580 1795.700 587.740 ;
        RECT 4.000 564.220 1796.340 586.580 ;
        RECT 4.000 563.060 1795.700 564.220 ;
        RECT 4.000 560.860 1796.340 563.060 ;
        RECT 4.300 559.700 1796.340 560.860 ;
        RECT 4.000 540.700 1796.340 559.700 ;
        RECT 4.000 539.540 1795.700 540.700 ;
        RECT 4.000 525.020 1796.340 539.540 ;
        RECT 4.300 523.860 1796.340 525.020 ;
        RECT 4.000 517.180 1796.340 523.860 ;
        RECT 4.000 516.020 1795.700 517.180 ;
        RECT 4.000 493.660 1796.340 516.020 ;
        RECT 4.000 492.500 1795.700 493.660 ;
        RECT 4.000 489.180 1796.340 492.500 ;
        RECT 4.300 488.020 1796.340 489.180 ;
        RECT 4.000 470.140 1796.340 488.020 ;
        RECT 4.000 468.980 1795.700 470.140 ;
        RECT 4.000 453.340 1796.340 468.980 ;
        RECT 4.300 452.180 1796.340 453.340 ;
        RECT 4.000 446.620 1796.340 452.180 ;
        RECT 4.000 445.460 1795.700 446.620 ;
        RECT 4.000 423.100 1796.340 445.460 ;
        RECT 4.000 421.940 1795.700 423.100 ;
        RECT 4.000 417.500 1796.340 421.940 ;
        RECT 4.300 416.340 1796.340 417.500 ;
        RECT 4.000 399.580 1796.340 416.340 ;
        RECT 4.000 398.420 1795.700 399.580 ;
        RECT 4.000 381.660 1796.340 398.420 ;
        RECT 4.300 380.500 1796.340 381.660 ;
        RECT 4.000 376.060 1796.340 380.500 ;
        RECT 4.000 374.900 1795.700 376.060 ;
        RECT 4.000 352.540 1796.340 374.900 ;
        RECT 4.000 351.380 1795.700 352.540 ;
        RECT 4.000 345.820 1796.340 351.380 ;
        RECT 4.300 344.660 1796.340 345.820 ;
        RECT 4.000 329.020 1796.340 344.660 ;
        RECT 4.000 327.860 1795.700 329.020 ;
        RECT 4.000 309.980 1796.340 327.860 ;
        RECT 4.300 308.820 1796.340 309.980 ;
        RECT 4.000 305.500 1796.340 308.820 ;
        RECT 4.000 304.340 1795.700 305.500 ;
        RECT 4.000 281.980 1796.340 304.340 ;
        RECT 4.000 280.820 1795.700 281.980 ;
        RECT 4.000 274.140 1796.340 280.820 ;
        RECT 4.300 272.980 1796.340 274.140 ;
        RECT 4.000 258.460 1796.340 272.980 ;
        RECT 4.000 257.300 1795.700 258.460 ;
        RECT 4.000 238.300 1796.340 257.300 ;
        RECT 4.300 237.140 1796.340 238.300 ;
        RECT 4.000 234.940 1796.340 237.140 ;
        RECT 4.000 233.780 1795.700 234.940 ;
        RECT 4.000 211.420 1796.340 233.780 ;
        RECT 4.000 210.260 1795.700 211.420 ;
        RECT 4.000 202.460 1796.340 210.260 ;
        RECT 4.300 201.300 1796.340 202.460 ;
        RECT 4.000 187.900 1796.340 201.300 ;
        RECT 4.000 186.740 1795.700 187.900 ;
        RECT 4.000 166.620 1796.340 186.740 ;
        RECT 4.300 165.460 1796.340 166.620 ;
        RECT 4.000 164.380 1796.340 165.460 ;
        RECT 4.000 163.220 1795.700 164.380 ;
        RECT 4.000 140.860 1796.340 163.220 ;
        RECT 4.000 139.700 1795.700 140.860 ;
        RECT 4.000 130.780 1796.340 139.700 ;
        RECT 4.300 129.620 1796.340 130.780 ;
        RECT 4.000 117.340 1796.340 129.620 ;
        RECT 4.000 116.180 1795.700 117.340 ;
        RECT 4.000 94.940 1796.340 116.180 ;
        RECT 4.300 93.820 1796.340 94.940 ;
        RECT 4.300 93.780 1795.700 93.820 ;
        RECT 4.000 92.660 1795.700 93.780 ;
        RECT 4.000 70.300 1796.340 92.660 ;
        RECT 4.000 69.140 1795.700 70.300 ;
        RECT 4.000 59.100 1796.340 69.140 ;
        RECT 4.300 57.940 1796.340 59.100 ;
        RECT 4.000 46.780 1796.340 57.940 ;
        RECT 4.000 45.620 1795.700 46.780 ;
        RECT 4.000 23.260 1796.340 45.620 ;
        RECT 4.300 22.100 1795.700 23.260 ;
        RECT 4.000 3.500 1796.340 22.100 ;
      LAYER Metal4 ;
        RECT 16.940 784.600 1777.300 786.150 ;
        RECT 16.940 15.080 21.940 784.600 ;
        RECT 24.140 15.080 98.740 784.600 ;
        RECT 100.940 15.080 175.540 784.600 ;
        RECT 177.740 15.080 252.340 784.600 ;
        RECT 254.540 15.080 329.140 784.600 ;
        RECT 331.340 15.080 405.940 784.600 ;
        RECT 408.140 15.080 482.740 784.600 ;
        RECT 484.940 15.080 559.540 784.600 ;
        RECT 561.740 15.080 636.340 784.600 ;
        RECT 638.540 15.080 713.140 784.600 ;
        RECT 715.340 15.080 789.940 784.600 ;
        RECT 792.140 15.080 866.740 784.600 ;
        RECT 868.940 15.080 943.540 784.600 ;
        RECT 945.740 15.080 1020.340 784.600 ;
        RECT 1022.540 15.080 1097.140 784.600 ;
        RECT 1099.340 15.080 1173.940 784.600 ;
        RECT 1176.140 15.080 1250.740 784.600 ;
        RECT 1252.940 15.080 1327.540 784.600 ;
        RECT 1329.740 15.080 1404.340 784.600 ;
        RECT 1406.540 15.080 1481.140 784.600 ;
        RECT 1483.340 15.080 1557.940 784.600 ;
        RECT 1560.140 15.080 1634.740 784.600 ;
        RECT 1636.940 15.080 1711.540 784.600 ;
        RECT 1713.740 15.080 1777.300 784.600 ;
        RECT 16.940 3.450 1777.300 15.080 ;
  END
END wrapped_pdp11
END LIBRARY

