VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN blinker_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 596.000 473.200 600.000 ;
    END
  END blinker_do[0]
  PIN blinker_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 596.000 478.800 600.000 ;
    END
  END blinker_do[1]
  PIN blinker_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 596.000 484.400 600.000 ;
    END
  END blinker_do[2]
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 200.480 600.000 201.040 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 245.280 600.000 245.840 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 249.760 600.000 250.320 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 254.240 600.000 254.800 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 258.720 600.000 259.280 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 263.200 600.000 263.760 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 267.680 600.000 268.240 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 272.160 600.000 272.720 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 276.640 600.000 277.200 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 281.120 600.000 281.680 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 285.600 600.000 286.160 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 204.960 600.000 205.520 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 290.080 600.000 290.640 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 294.560 600.000 295.120 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 299.040 600.000 299.600 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 303.520 600.000 304.080 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 308.000 600.000 308.560 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 312.480 600.000 313.040 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 316.960 600.000 317.520 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 321.440 600.000 322.000 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 325.920 600.000 326.480 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 330.400 600.000 330.960 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 209.440 600.000 210.000 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 334.880 600.000 335.440 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 339.360 600.000 339.920 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 213.920 600.000 214.480 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 218.400 600.000 218.960 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 222.880 600.000 223.440 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 227.360 600.000 227.920 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 231.840 600.000 232.400 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 236.320 600.000 236.880 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 240.800 600.000 241.360 ;
    END
  END custom_settings[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 596.000 25.200 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 596.000 81.200 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 596.000 86.800 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 596.000 92.400 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 596.000 98.000 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 596.000 103.600 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 596.000 109.200 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 596.000 114.800 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 596.000 120.400 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 596.000 126.000 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 596.000 131.600 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 596.000 30.800 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 596.000 137.200 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 596.000 142.800 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 596.000 148.400 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 596.000 154.000 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 596.000 159.600 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 596.000 165.200 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 596.000 170.800 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 596.000 176.400 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 596.000 182.000 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 596.000 187.600 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 596.000 36.400 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 596.000 193.200 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 596.000 198.800 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 596.000 204.400 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 596.000 210.000 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 596.000 215.600 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 596.000 221.200 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 596.000 226.800 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 596.000 232.400 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 596.000 42.000 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 596.000 47.600 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 596.000 53.200 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 596.000 58.800 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 596.000 64.400 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 596.000 70.000 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 596.000 75.600 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 4.000 95.760 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.400 4.000 50.960 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.600 4.000 90.160 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 596.000 238.000 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 596.000 294.000 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 596.000 299.600 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 596.000 305.200 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 596.000 310.800 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 596.000 316.400 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 596.000 322.000 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 596.000 327.600 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 596.000 333.200 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 596.000 338.800 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 596.000 344.400 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 596.000 243.600 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 596.000 350.000 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 596.000 355.600 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 596.000 361.200 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 596.000 366.800 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 596.000 372.400 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 596.000 378.000 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 596.000 383.600 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 596.000 389.200 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 596.000 394.800 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 596.000 400.400 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 596.000 249.200 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 596.000 406.000 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 596.000 411.600 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 596.000 417.200 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 596.000 422.800 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 596.000 428.400 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 596.000 434.000 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 596.000 439.600 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 596.000 445.200 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 596.000 254.800 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 596.000 260.400 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 596.000 266.000 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 596.000 271.600 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 596.000 277.200 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 596.000 282.800 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 596.000 288.400 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 596.000 450.800 600.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 596.000 456.400 600.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 596.000 462.000 600.000 ;
    END
  END irq[2]
  PIN mc14500_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END mc14500_do[0]
  PIN mc14500_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END mc14500_do[10]
  PIN mc14500_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END mc14500_do[11]
  PIN mc14500_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END mc14500_do[12]
  PIN mc14500_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 464.800 4.000 465.360 ;
    END
  END mc14500_do[13]
  PIN mc14500_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END mc14500_do[14]
  PIN mc14500_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END mc14500_do[15]
  PIN mc14500_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END mc14500_do[16]
  PIN mc14500_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 487.200 4.000 487.760 ;
    END
  END mc14500_do[17]
  PIN mc14500_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.800 4.000 493.360 ;
    END
  END mc14500_do[18]
  PIN mc14500_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 498.400 4.000 498.960 ;
    END
  END mc14500_do[19]
  PIN mc14500_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 397.600 4.000 398.160 ;
    END
  END mc14500_do[1]
  PIN mc14500_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END mc14500_do[20]
  PIN mc14500_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END mc14500_do[21]
  PIN mc14500_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.200 4.000 515.760 ;
    END
  END mc14500_do[22]
  PIN mc14500_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 520.800 4.000 521.360 ;
    END
  END mc14500_do[23]
  PIN mc14500_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.400 4.000 526.960 ;
    END
  END mc14500_do[24]
  PIN mc14500_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 532.000 4.000 532.560 ;
    END
  END mc14500_do[25]
  PIN mc14500_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END mc14500_do[26]
  PIN mc14500_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END mc14500_do[27]
  PIN mc14500_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END mc14500_do[28]
  PIN mc14500_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 554.400 4.000 554.960 ;
    END
  END mc14500_do[29]
  PIN mc14500_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END mc14500_do[2]
  PIN mc14500_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END mc14500_do[30]
  PIN mc14500_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END mc14500_do[3]
  PIN mc14500_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 414.400 4.000 414.960 ;
    END
  END mc14500_do[4]
  PIN mc14500_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 420.000 4.000 420.560 ;
    END
  END mc14500_do[5]
  PIN mc14500_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END mc14500_do[6]
  PIN mc14500_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 431.200 4.000 431.760 ;
    END
  END mc14500_do[7]
  PIN mc14500_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END mc14500_do[8]
  PIN mc14500_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END mc14500_do[9]
  PIN mc14500_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 596.000 495.600 600.000 ;
    END
  END mc14500_sram_addr[0]
  PIN mc14500_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 596.000 501.200 600.000 ;
    END
  END mc14500_sram_addr[1]
  PIN mc14500_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 506.240 596.000 506.800 600.000 ;
    END
  END mc14500_sram_addr[2]
  PIN mc14500_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 596.000 512.400 600.000 ;
    END
  END mc14500_sram_addr[3]
  PIN mc14500_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 596.000 518.000 600.000 ;
    END
  END mc14500_sram_addr[4]
  PIN mc14500_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 596.000 523.600 600.000 ;
    END
  END mc14500_sram_addr[5]
  PIN mc14500_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 573.440 596.000 574.000 600.000 ;
    END
  END mc14500_sram_gwe
  PIN mc14500_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 596.000 529.200 600.000 ;
    END
  END mc14500_sram_in[0]
  PIN mc14500_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 596.000 534.800 600.000 ;
    END
  END mc14500_sram_in[1]
  PIN mc14500_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 596.000 540.400 600.000 ;
    END
  END mc14500_sram_in[2]
  PIN mc14500_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 545.440 596.000 546.000 600.000 ;
    END
  END mc14500_sram_in[3]
  PIN mc14500_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 596.000 551.600 600.000 ;
    END
  END mc14500_sram_in[4]
  PIN mc14500_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 596.000 557.200 600.000 ;
    END
  END mc14500_sram_in[5]
  PIN mc14500_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 596.000 562.800 600.000 ;
    END
  END mc14500_sram_in[6]
  PIN mc14500_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 596.000 568.400 600.000 ;
    END
  END mc14500_sram_in[7]
  PIN qcpu_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 0.000 422.800 4.000 ;
    END
  END qcpu_do[0]
  PIN qcpu_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 0.000 467.600 4.000 ;
    END
  END qcpu_do[10]
  PIN qcpu_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 0.000 472.080 4.000 ;
    END
  END qcpu_do[11]
  PIN qcpu_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 0.000 476.560 4.000 ;
    END
  END qcpu_do[12]
  PIN qcpu_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END qcpu_do[13]
  PIN qcpu_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 0.000 485.520 4.000 ;
    END
  END qcpu_do[14]
  PIN qcpu_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END qcpu_do[15]
  PIN qcpu_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 0.000 494.480 4.000 ;
    END
  END qcpu_do[16]
  PIN qcpu_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END qcpu_do[17]
  PIN qcpu_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END qcpu_do[18]
  PIN qcpu_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END qcpu_do[19]
  PIN qcpu_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END qcpu_do[1]
  PIN qcpu_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 511.840 0.000 512.400 4.000 ;
    END
  END qcpu_do[20]
  PIN qcpu_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END qcpu_do[21]
  PIN qcpu_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 0.000 521.360 4.000 ;
    END
  END qcpu_do[22]
  PIN qcpu_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END qcpu_do[23]
  PIN qcpu_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END qcpu_do[24]
  PIN qcpu_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END qcpu_do[25]
  PIN qcpu_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 0.000 539.280 4.000 ;
    END
  END qcpu_do[26]
  PIN qcpu_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END qcpu_do[27]
  PIN qcpu_do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 0.000 548.240 4.000 ;
    END
  END qcpu_do[28]
  PIN qcpu_do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 0.000 552.720 4.000 ;
    END
  END qcpu_do[29]
  PIN qcpu_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 0.000 431.760 4.000 ;
    END
  END qcpu_do[2]
  PIN qcpu_do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 0.000 557.200 4.000 ;
    END
  END qcpu_do[30]
  PIN qcpu_do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END qcpu_do[31]
  PIN qcpu_do[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 0.000 566.160 4.000 ;
    END
  END qcpu_do[32]
  PIN qcpu_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END qcpu_do[3]
  PIN qcpu_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 0.000 440.720 4.000 ;
    END
  END qcpu_do[4]
  PIN qcpu_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 0.000 445.200 4.000 ;
    END
  END qcpu_do[5]
  PIN qcpu_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END qcpu_do[6]
  PIN qcpu_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END qcpu_do[7]
  PIN qcpu_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 4.000 ;
    END
  END qcpu_do[8]
  PIN qcpu_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 0.000 463.120 4.000 ;
    END
  END qcpu_do[9]
  PIN qcpu_oeb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 343.840 600.000 344.400 ;
    END
  END qcpu_oeb[0]
  PIN qcpu_oeb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 388.640 600.000 389.200 ;
    END
  END qcpu_oeb[10]
  PIN qcpu_oeb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 393.120 600.000 393.680 ;
    END
  END qcpu_oeb[11]
  PIN qcpu_oeb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 397.600 600.000 398.160 ;
    END
  END qcpu_oeb[12]
  PIN qcpu_oeb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 402.080 600.000 402.640 ;
    END
  END qcpu_oeb[13]
  PIN qcpu_oeb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 406.560 600.000 407.120 ;
    END
  END qcpu_oeb[14]
  PIN qcpu_oeb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 411.040 600.000 411.600 ;
    END
  END qcpu_oeb[15]
  PIN qcpu_oeb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 415.520 600.000 416.080 ;
    END
  END qcpu_oeb[16]
  PIN qcpu_oeb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 420.000 600.000 420.560 ;
    END
  END qcpu_oeb[17]
  PIN qcpu_oeb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 424.480 600.000 425.040 ;
    END
  END qcpu_oeb[18]
  PIN qcpu_oeb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 428.960 600.000 429.520 ;
    END
  END qcpu_oeb[19]
  PIN qcpu_oeb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 348.320 600.000 348.880 ;
    END
  END qcpu_oeb[1]
  PIN qcpu_oeb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 433.440 600.000 434.000 ;
    END
  END qcpu_oeb[20]
  PIN qcpu_oeb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 437.920 600.000 438.480 ;
    END
  END qcpu_oeb[21]
  PIN qcpu_oeb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 442.400 600.000 442.960 ;
    END
  END qcpu_oeb[22]
  PIN qcpu_oeb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 446.880 600.000 447.440 ;
    END
  END qcpu_oeb[23]
  PIN qcpu_oeb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 451.360 600.000 451.920 ;
    END
  END qcpu_oeb[24]
  PIN qcpu_oeb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 455.840 600.000 456.400 ;
    END
  END qcpu_oeb[25]
  PIN qcpu_oeb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 460.320 600.000 460.880 ;
    END
  END qcpu_oeb[26]
  PIN qcpu_oeb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 464.800 600.000 465.360 ;
    END
  END qcpu_oeb[27]
  PIN qcpu_oeb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 469.280 600.000 469.840 ;
    END
  END qcpu_oeb[28]
  PIN qcpu_oeb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 473.760 600.000 474.320 ;
    END
  END qcpu_oeb[29]
  PIN qcpu_oeb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 352.800 600.000 353.360 ;
    END
  END qcpu_oeb[2]
  PIN qcpu_oeb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 478.240 600.000 478.800 ;
    END
  END qcpu_oeb[30]
  PIN qcpu_oeb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 482.720 600.000 483.280 ;
    END
  END qcpu_oeb[31]
  PIN qcpu_oeb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 487.200 600.000 487.760 ;
    END
  END qcpu_oeb[32]
  PIN qcpu_oeb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 357.280 600.000 357.840 ;
    END
  END qcpu_oeb[3]
  PIN qcpu_oeb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 361.760 600.000 362.320 ;
    END
  END qcpu_oeb[4]
  PIN qcpu_oeb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 366.240 600.000 366.800 ;
    END
  END qcpu_oeb[5]
  PIN qcpu_oeb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 370.720 600.000 371.280 ;
    END
  END qcpu_oeb[6]
  PIN qcpu_oeb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 375.200 600.000 375.760 ;
    END
  END qcpu_oeb[7]
  PIN qcpu_oeb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 379.680 600.000 380.240 ;
    END
  END qcpu_oeb[8]
  PIN qcpu_oeb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 384.160 600.000 384.720 ;
    END
  END qcpu_oeb[9]
  PIN qcpu_sram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END qcpu_sram_addr[0]
  PIN qcpu_sram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END qcpu_sram_addr[1]
  PIN qcpu_sram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END qcpu_sram_addr[2]
  PIN qcpu_sram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 0.000 584.080 4.000 ;
    END
  END qcpu_sram_addr[3]
  PIN qcpu_sram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END qcpu_sram_addr[4]
  PIN qcpu_sram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 592.480 0.000 593.040 4.000 ;
    END
  END qcpu_sram_addr[5]
  PIN qcpu_sram_gwe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 0.000 597.520 4.000 ;
    END
  END qcpu_sram_gwe
  PIN qcpu_sram_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 491.680 600.000 492.240 ;
    END
  END qcpu_sram_in[0]
  PIN qcpu_sram_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 496.160 600.000 496.720 ;
    END
  END qcpu_sram_in[1]
  PIN qcpu_sram_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 500.640 600.000 501.200 ;
    END
  END qcpu_sram_in[2]
  PIN qcpu_sram_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 505.120 600.000 505.680 ;
    END
  END qcpu_sram_in[3]
  PIN qcpu_sram_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 509.600 600.000 510.160 ;
    END
  END qcpu_sram_in[4]
  PIN qcpu_sram_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 514.080 600.000 514.640 ;
    END
  END qcpu_sram_in[5]
  PIN qcpu_sram_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 518.560 600.000 519.120 ;
    END
  END qcpu_sram_in[6]
  PIN qcpu_sram_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 523.040 600.000 523.600 ;
    END
  END qcpu_sram_in[7]
  PIN qcpu_sram_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 527.520 600.000 528.080 ;
    END
  END qcpu_sram_out[0]
  PIN qcpu_sram_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 532.000 600.000 532.560 ;
    END
  END qcpu_sram_out[1]
  PIN qcpu_sram_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 536.480 600.000 537.040 ;
    END
  END qcpu_sram_out[2]
  PIN qcpu_sram_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 540.960 600.000 541.520 ;
    END
  END qcpu_sram_out[3]
  PIN qcpu_sram_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 545.440 600.000 546.000 ;
    END
  END qcpu_sram_out[4]
  PIN qcpu_sram_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 549.920 600.000 550.480 ;
    END
  END qcpu_sram_out[5]
  PIN qcpu_sram_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 554.400 600.000 554.960 ;
    END
  END qcpu_sram_out[6]
  PIN qcpu_sram_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 558.880 600.000 559.440 ;
    END
  END qcpu_sram_out[7]
  PIN rst_blinker
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 596.000 467.600 600.000 ;
    END
  END rst_blinker
  PIN rst_mc14500
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END rst_mc14500
  PIN rst_qcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.800 4.000 381.360 ;
    END
  END rst_qcpu
  PIN rst_sid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END rst_sid
  PIN rst_sn76489
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 596.000 490.000 600.000 ;
    END
  END rst_sn76489
  PIN sid_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END sid_do[0]
  PIN sid_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END sid_do[10]
  PIN sid_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END sid_do[11]
  PIN sid_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END sid_do[12]
  PIN sid_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.400 4.000 330.960 ;
    END
  END sid_do[13]
  PIN sid_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END sid_do[14]
  PIN sid_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END sid_do[15]
  PIN sid_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.200 4.000 347.760 ;
    END
  END sid_do[16]
  PIN sid_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.800 4.000 353.360 ;
    END
  END sid_do[17]
  PIN sid_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END sid_do[18]
  PIN sid_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END sid_do[19]
  PIN sid_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END sid_do[1]
  PIN sid_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END sid_do[20]
  PIN sid_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END sid_do[2]
  PIN sid_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END sid_do[3]
  PIN sid_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END sid_do[4]
  PIN sid_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END sid_do[5]
  PIN sid_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END sid_do[6]
  PIN sid_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END sid_do[7]
  PIN sid_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END sid_do[8]
  PIN sid_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END sid_do[9]
  PIN sid_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END sid_oeb
  PIN sn76489_do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 0.000 297.360 4.000 ;
    END
  END sn76489_do[0]
  PIN sn76489_do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 0.000 342.160 4.000 ;
    END
  END sn76489_do[10]
  PIN sn76489_do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END sn76489_do[11]
  PIN sn76489_do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 350.560 0.000 351.120 4.000 ;
    END
  END sn76489_do[12]
  PIN sn76489_do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 0.000 355.600 4.000 ;
    END
  END sn76489_do[13]
  PIN sn76489_do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END sn76489_do[14]
  PIN sn76489_do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END sn76489_do[15]
  PIN sn76489_do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END sn76489_do[16]
  PIN sn76489_do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END sn76489_do[17]
  PIN sn76489_do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 0.000 378.000 4.000 ;
    END
  END sn76489_do[18]
  PIN sn76489_do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 0.000 382.480 4.000 ;
    END
  END sn76489_do[19]
  PIN sn76489_do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END sn76489_do[1]
  PIN sn76489_do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END sn76489_do[20]
  PIN sn76489_do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END sn76489_do[21]
  PIN sn76489_do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 0.000 395.920 4.000 ;
    END
  END sn76489_do[22]
  PIN sn76489_do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END sn76489_do[23]
  PIN sn76489_do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 404.320 0.000 404.880 4.000 ;
    END
  END sn76489_do[24]
  PIN sn76489_do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END sn76489_do[25]
  PIN sn76489_do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 0.000 413.840 4.000 ;
    END
  END sn76489_do[26]
  PIN sn76489_do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 0.000 418.320 4.000 ;
    END
  END sn76489_do[27]
  PIN sn76489_do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 0.000 306.320 4.000 ;
    END
  END sn76489_do[2]
  PIN sn76489_do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END sn76489_do[3]
  PIN sn76489_do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 0.000 315.280 4.000 ;
    END
  END sn76489_do[4]
  PIN sn76489_do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END sn76489_do[5]
  PIN sn76489_do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 323.680 0.000 324.240 4.000 ;
    END
  END sn76489_do[6]
  PIN sn76489_do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END sn76489_do[7]
  PIN sn76489_do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 0.000 333.200 4.000 ;
    END
  END sn76489_do[8]
  PIN sn76489_do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 0.000 337.680 4.000 ;
    END
  END sn76489_do[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1.120 0.000 1.680 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 196.000 600.000 196.560 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 0.000 55.440 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 0.000 82.320 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 0.000 136.080 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 0.000 145.040 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 0.000 28.560 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 187.040 600.000 187.600 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 0.000 216.720 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 243.040 0.000 243.600 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 0.000 252.560 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 0.000 171.920 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 0.000 189.840 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 39.200 600.000 39.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 84.000 600.000 84.560 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 88.480 600.000 89.040 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 92.960 600.000 93.520 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 97.440 600.000 98.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 101.920 600.000 102.480 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 106.400 600.000 106.960 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 110.880 600.000 111.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 115.360 600.000 115.920 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 119.840 600.000 120.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 124.320 600.000 124.880 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 43.680 600.000 44.240 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 128.800 600.000 129.360 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 133.280 600.000 133.840 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 137.760 600.000 138.320 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 142.240 600.000 142.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 146.720 600.000 147.280 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 151.200 600.000 151.760 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 155.680 600.000 156.240 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 160.160 600.000 160.720 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 164.640 600.000 165.200 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 169.120 600.000 169.680 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 48.160 600.000 48.720 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 173.600 600.000 174.160 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 178.080 600.000 178.640 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 52.640 600.000 53.200 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 57.120 600.000 57.680 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 61.600 600.000 62.160 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 66.080 600.000 66.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 70.560 600.000 71.120 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 75.040 600.000 75.600 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 79.520 600.000 80.080 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 191.520 600.000 192.080 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 596.000 182.560 600.000 183.120 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 593.040 586.730 ;
      LAYER Metal2 ;
        RECT 1.260 595.700 24.340 596.820 ;
        RECT 25.500 595.700 29.940 596.820 ;
        RECT 31.100 595.700 35.540 596.820 ;
        RECT 36.700 595.700 41.140 596.820 ;
        RECT 42.300 595.700 46.740 596.820 ;
        RECT 47.900 595.700 52.340 596.820 ;
        RECT 53.500 595.700 57.940 596.820 ;
        RECT 59.100 595.700 63.540 596.820 ;
        RECT 64.700 595.700 69.140 596.820 ;
        RECT 70.300 595.700 74.740 596.820 ;
        RECT 75.900 595.700 80.340 596.820 ;
        RECT 81.500 595.700 85.940 596.820 ;
        RECT 87.100 595.700 91.540 596.820 ;
        RECT 92.700 595.700 97.140 596.820 ;
        RECT 98.300 595.700 102.740 596.820 ;
        RECT 103.900 595.700 108.340 596.820 ;
        RECT 109.500 595.700 113.940 596.820 ;
        RECT 115.100 595.700 119.540 596.820 ;
        RECT 120.700 595.700 125.140 596.820 ;
        RECT 126.300 595.700 130.740 596.820 ;
        RECT 131.900 595.700 136.340 596.820 ;
        RECT 137.500 595.700 141.940 596.820 ;
        RECT 143.100 595.700 147.540 596.820 ;
        RECT 148.700 595.700 153.140 596.820 ;
        RECT 154.300 595.700 158.740 596.820 ;
        RECT 159.900 595.700 164.340 596.820 ;
        RECT 165.500 595.700 169.940 596.820 ;
        RECT 171.100 595.700 175.540 596.820 ;
        RECT 176.700 595.700 181.140 596.820 ;
        RECT 182.300 595.700 186.740 596.820 ;
        RECT 187.900 595.700 192.340 596.820 ;
        RECT 193.500 595.700 197.940 596.820 ;
        RECT 199.100 595.700 203.540 596.820 ;
        RECT 204.700 595.700 209.140 596.820 ;
        RECT 210.300 595.700 214.740 596.820 ;
        RECT 215.900 595.700 220.340 596.820 ;
        RECT 221.500 595.700 225.940 596.820 ;
        RECT 227.100 595.700 231.540 596.820 ;
        RECT 232.700 595.700 237.140 596.820 ;
        RECT 238.300 595.700 242.740 596.820 ;
        RECT 243.900 595.700 248.340 596.820 ;
        RECT 249.500 595.700 253.940 596.820 ;
        RECT 255.100 595.700 259.540 596.820 ;
        RECT 260.700 595.700 265.140 596.820 ;
        RECT 266.300 595.700 270.740 596.820 ;
        RECT 271.900 595.700 276.340 596.820 ;
        RECT 277.500 595.700 281.940 596.820 ;
        RECT 283.100 595.700 287.540 596.820 ;
        RECT 288.700 595.700 293.140 596.820 ;
        RECT 294.300 595.700 298.740 596.820 ;
        RECT 299.900 595.700 304.340 596.820 ;
        RECT 305.500 595.700 309.940 596.820 ;
        RECT 311.100 595.700 315.540 596.820 ;
        RECT 316.700 595.700 321.140 596.820 ;
        RECT 322.300 595.700 326.740 596.820 ;
        RECT 327.900 595.700 332.340 596.820 ;
        RECT 333.500 595.700 337.940 596.820 ;
        RECT 339.100 595.700 343.540 596.820 ;
        RECT 344.700 595.700 349.140 596.820 ;
        RECT 350.300 595.700 354.740 596.820 ;
        RECT 355.900 595.700 360.340 596.820 ;
        RECT 361.500 595.700 365.940 596.820 ;
        RECT 367.100 595.700 371.540 596.820 ;
        RECT 372.700 595.700 377.140 596.820 ;
        RECT 378.300 595.700 382.740 596.820 ;
        RECT 383.900 595.700 388.340 596.820 ;
        RECT 389.500 595.700 393.940 596.820 ;
        RECT 395.100 595.700 399.540 596.820 ;
        RECT 400.700 595.700 405.140 596.820 ;
        RECT 406.300 595.700 410.740 596.820 ;
        RECT 411.900 595.700 416.340 596.820 ;
        RECT 417.500 595.700 421.940 596.820 ;
        RECT 423.100 595.700 427.540 596.820 ;
        RECT 428.700 595.700 433.140 596.820 ;
        RECT 434.300 595.700 438.740 596.820 ;
        RECT 439.900 595.700 444.340 596.820 ;
        RECT 445.500 595.700 449.940 596.820 ;
        RECT 451.100 595.700 455.540 596.820 ;
        RECT 456.700 595.700 461.140 596.820 ;
        RECT 462.300 595.700 466.740 596.820 ;
        RECT 467.900 595.700 472.340 596.820 ;
        RECT 473.500 595.700 477.940 596.820 ;
        RECT 479.100 595.700 483.540 596.820 ;
        RECT 484.700 595.700 489.140 596.820 ;
        RECT 490.300 595.700 494.740 596.820 ;
        RECT 495.900 595.700 500.340 596.820 ;
        RECT 501.500 595.700 505.940 596.820 ;
        RECT 507.100 595.700 511.540 596.820 ;
        RECT 512.700 595.700 517.140 596.820 ;
        RECT 518.300 595.700 522.740 596.820 ;
        RECT 523.900 595.700 528.340 596.820 ;
        RECT 529.500 595.700 533.940 596.820 ;
        RECT 535.100 595.700 539.540 596.820 ;
        RECT 540.700 595.700 545.140 596.820 ;
        RECT 546.300 595.700 550.740 596.820 ;
        RECT 551.900 595.700 556.340 596.820 ;
        RECT 557.500 595.700 561.940 596.820 ;
        RECT 563.100 595.700 567.540 596.820 ;
        RECT 568.700 595.700 573.140 596.820 ;
        RECT 574.300 595.700 597.380 596.820 ;
        RECT 1.260 4.300 597.380 595.700 ;
        RECT 1.980 3.500 5.300 4.300 ;
        RECT 6.460 3.500 9.780 4.300 ;
        RECT 10.940 3.500 14.260 4.300 ;
        RECT 15.420 3.500 18.740 4.300 ;
        RECT 19.900 3.500 23.220 4.300 ;
        RECT 24.380 3.500 27.700 4.300 ;
        RECT 28.860 3.500 32.180 4.300 ;
        RECT 33.340 3.500 36.660 4.300 ;
        RECT 37.820 3.500 41.140 4.300 ;
        RECT 42.300 3.500 45.620 4.300 ;
        RECT 46.780 3.500 50.100 4.300 ;
        RECT 51.260 3.500 54.580 4.300 ;
        RECT 55.740 3.500 59.060 4.300 ;
        RECT 60.220 3.500 63.540 4.300 ;
        RECT 64.700 3.500 68.020 4.300 ;
        RECT 69.180 3.500 72.500 4.300 ;
        RECT 73.660 3.500 76.980 4.300 ;
        RECT 78.140 3.500 81.460 4.300 ;
        RECT 82.620 3.500 85.940 4.300 ;
        RECT 87.100 3.500 90.420 4.300 ;
        RECT 91.580 3.500 94.900 4.300 ;
        RECT 96.060 3.500 99.380 4.300 ;
        RECT 100.540 3.500 103.860 4.300 ;
        RECT 105.020 3.500 108.340 4.300 ;
        RECT 109.500 3.500 112.820 4.300 ;
        RECT 113.980 3.500 117.300 4.300 ;
        RECT 118.460 3.500 121.780 4.300 ;
        RECT 122.940 3.500 126.260 4.300 ;
        RECT 127.420 3.500 130.740 4.300 ;
        RECT 131.900 3.500 135.220 4.300 ;
        RECT 136.380 3.500 139.700 4.300 ;
        RECT 140.860 3.500 144.180 4.300 ;
        RECT 145.340 3.500 148.660 4.300 ;
        RECT 149.820 3.500 153.140 4.300 ;
        RECT 154.300 3.500 157.620 4.300 ;
        RECT 158.780 3.500 162.100 4.300 ;
        RECT 163.260 3.500 166.580 4.300 ;
        RECT 167.740 3.500 171.060 4.300 ;
        RECT 172.220 3.500 175.540 4.300 ;
        RECT 176.700 3.500 180.020 4.300 ;
        RECT 181.180 3.500 184.500 4.300 ;
        RECT 185.660 3.500 188.980 4.300 ;
        RECT 190.140 3.500 193.460 4.300 ;
        RECT 194.620 3.500 197.940 4.300 ;
        RECT 199.100 3.500 202.420 4.300 ;
        RECT 203.580 3.500 206.900 4.300 ;
        RECT 208.060 3.500 211.380 4.300 ;
        RECT 212.540 3.500 215.860 4.300 ;
        RECT 217.020 3.500 220.340 4.300 ;
        RECT 221.500 3.500 224.820 4.300 ;
        RECT 225.980 3.500 229.300 4.300 ;
        RECT 230.460 3.500 233.780 4.300 ;
        RECT 234.940 3.500 238.260 4.300 ;
        RECT 239.420 3.500 242.740 4.300 ;
        RECT 243.900 3.500 247.220 4.300 ;
        RECT 248.380 3.500 251.700 4.300 ;
        RECT 252.860 3.500 256.180 4.300 ;
        RECT 257.340 3.500 260.660 4.300 ;
        RECT 261.820 3.500 265.140 4.300 ;
        RECT 266.300 3.500 269.620 4.300 ;
        RECT 270.780 3.500 274.100 4.300 ;
        RECT 275.260 3.500 278.580 4.300 ;
        RECT 279.740 3.500 283.060 4.300 ;
        RECT 284.220 3.500 287.540 4.300 ;
        RECT 288.700 3.500 292.020 4.300 ;
        RECT 293.180 3.500 296.500 4.300 ;
        RECT 297.660 3.500 300.980 4.300 ;
        RECT 302.140 3.500 305.460 4.300 ;
        RECT 306.620 3.500 309.940 4.300 ;
        RECT 311.100 3.500 314.420 4.300 ;
        RECT 315.580 3.500 318.900 4.300 ;
        RECT 320.060 3.500 323.380 4.300 ;
        RECT 324.540 3.500 327.860 4.300 ;
        RECT 329.020 3.500 332.340 4.300 ;
        RECT 333.500 3.500 336.820 4.300 ;
        RECT 337.980 3.500 341.300 4.300 ;
        RECT 342.460 3.500 345.780 4.300 ;
        RECT 346.940 3.500 350.260 4.300 ;
        RECT 351.420 3.500 354.740 4.300 ;
        RECT 355.900 3.500 359.220 4.300 ;
        RECT 360.380 3.500 363.700 4.300 ;
        RECT 364.860 3.500 368.180 4.300 ;
        RECT 369.340 3.500 372.660 4.300 ;
        RECT 373.820 3.500 377.140 4.300 ;
        RECT 378.300 3.500 381.620 4.300 ;
        RECT 382.780 3.500 386.100 4.300 ;
        RECT 387.260 3.500 390.580 4.300 ;
        RECT 391.740 3.500 395.060 4.300 ;
        RECT 396.220 3.500 399.540 4.300 ;
        RECT 400.700 3.500 404.020 4.300 ;
        RECT 405.180 3.500 408.500 4.300 ;
        RECT 409.660 3.500 412.980 4.300 ;
        RECT 414.140 3.500 417.460 4.300 ;
        RECT 418.620 3.500 421.940 4.300 ;
        RECT 423.100 3.500 426.420 4.300 ;
        RECT 427.580 3.500 430.900 4.300 ;
        RECT 432.060 3.500 435.380 4.300 ;
        RECT 436.540 3.500 439.860 4.300 ;
        RECT 441.020 3.500 444.340 4.300 ;
        RECT 445.500 3.500 448.820 4.300 ;
        RECT 449.980 3.500 453.300 4.300 ;
        RECT 454.460 3.500 457.780 4.300 ;
        RECT 458.940 3.500 462.260 4.300 ;
        RECT 463.420 3.500 466.740 4.300 ;
        RECT 467.900 3.500 471.220 4.300 ;
        RECT 472.380 3.500 475.700 4.300 ;
        RECT 476.860 3.500 480.180 4.300 ;
        RECT 481.340 3.500 484.660 4.300 ;
        RECT 485.820 3.500 489.140 4.300 ;
        RECT 490.300 3.500 493.620 4.300 ;
        RECT 494.780 3.500 498.100 4.300 ;
        RECT 499.260 3.500 502.580 4.300 ;
        RECT 503.740 3.500 507.060 4.300 ;
        RECT 508.220 3.500 511.540 4.300 ;
        RECT 512.700 3.500 516.020 4.300 ;
        RECT 517.180 3.500 520.500 4.300 ;
        RECT 521.660 3.500 524.980 4.300 ;
        RECT 526.140 3.500 529.460 4.300 ;
        RECT 530.620 3.500 533.940 4.300 ;
        RECT 535.100 3.500 538.420 4.300 ;
        RECT 539.580 3.500 542.900 4.300 ;
        RECT 544.060 3.500 547.380 4.300 ;
        RECT 548.540 3.500 551.860 4.300 ;
        RECT 553.020 3.500 556.340 4.300 ;
        RECT 557.500 3.500 560.820 4.300 ;
        RECT 561.980 3.500 565.300 4.300 ;
        RECT 566.460 3.500 569.780 4.300 ;
        RECT 570.940 3.500 574.260 4.300 ;
        RECT 575.420 3.500 578.740 4.300 ;
        RECT 579.900 3.500 583.220 4.300 ;
        RECT 584.380 3.500 587.700 4.300 ;
        RECT 588.860 3.500 592.180 4.300 ;
        RECT 593.340 3.500 596.660 4.300 ;
      LAYER Metal3 ;
        RECT 1.210 560.860 597.430 587.860 ;
        RECT 4.300 559.740 597.430 560.860 ;
        RECT 4.300 559.700 595.700 559.740 ;
        RECT 1.210 558.580 595.700 559.700 ;
        RECT 1.210 555.260 597.430 558.580 ;
        RECT 4.300 554.100 595.700 555.260 ;
        RECT 1.210 550.780 597.430 554.100 ;
        RECT 1.210 549.660 595.700 550.780 ;
        RECT 4.300 549.620 595.700 549.660 ;
        RECT 4.300 548.500 597.430 549.620 ;
        RECT 1.210 546.300 597.430 548.500 ;
        RECT 1.210 545.140 595.700 546.300 ;
        RECT 1.210 544.060 597.430 545.140 ;
        RECT 4.300 542.900 597.430 544.060 ;
        RECT 1.210 541.820 597.430 542.900 ;
        RECT 1.210 540.660 595.700 541.820 ;
        RECT 1.210 538.460 597.430 540.660 ;
        RECT 4.300 537.340 597.430 538.460 ;
        RECT 4.300 537.300 595.700 537.340 ;
        RECT 1.210 536.180 595.700 537.300 ;
        RECT 1.210 532.860 597.430 536.180 ;
        RECT 4.300 531.700 595.700 532.860 ;
        RECT 1.210 528.380 597.430 531.700 ;
        RECT 1.210 527.260 595.700 528.380 ;
        RECT 4.300 527.220 595.700 527.260 ;
        RECT 4.300 526.100 597.430 527.220 ;
        RECT 1.210 523.900 597.430 526.100 ;
        RECT 1.210 522.740 595.700 523.900 ;
        RECT 1.210 521.660 597.430 522.740 ;
        RECT 4.300 520.500 597.430 521.660 ;
        RECT 1.210 519.420 597.430 520.500 ;
        RECT 1.210 518.260 595.700 519.420 ;
        RECT 1.210 516.060 597.430 518.260 ;
        RECT 4.300 514.940 597.430 516.060 ;
        RECT 4.300 514.900 595.700 514.940 ;
        RECT 1.210 513.780 595.700 514.900 ;
        RECT 1.210 510.460 597.430 513.780 ;
        RECT 4.300 509.300 595.700 510.460 ;
        RECT 1.210 505.980 597.430 509.300 ;
        RECT 1.210 504.860 595.700 505.980 ;
        RECT 4.300 504.820 595.700 504.860 ;
        RECT 4.300 503.700 597.430 504.820 ;
        RECT 1.210 501.500 597.430 503.700 ;
        RECT 1.210 500.340 595.700 501.500 ;
        RECT 1.210 499.260 597.430 500.340 ;
        RECT 4.300 498.100 597.430 499.260 ;
        RECT 1.210 497.020 597.430 498.100 ;
        RECT 1.210 495.860 595.700 497.020 ;
        RECT 1.210 493.660 597.430 495.860 ;
        RECT 4.300 492.540 597.430 493.660 ;
        RECT 4.300 492.500 595.700 492.540 ;
        RECT 1.210 491.380 595.700 492.500 ;
        RECT 1.210 488.060 597.430 491.380 ;
        RECT 4.300 486.900 595.700 488.060 ;
        RECT 1.210 483.580 597.430 486.900 ;
        RECT 1.210 482.460 595.700 483.580 ;
        RECT 4.300 482.420 595.700 482.460 ;
        RECT 4.300 481.300 597.430 482.420 ;
        RECT 1.210 479.100 597.430 481.300 ;
        RECT 1.210 477.940 595.700 479.100 ;
        RECT 1.210 476.860 597.430 477.940 ;
        RECT 4.300 475.700 597.430 476.860 ;
        RECT 1.210 474.620 597.430 475.700 ;
        RECT 1.210 473.460 595.700 474.620 ;
        RECT 1.210 471.260 597.430 473.460 ;
        RECT 4.300 470.140 597.430 471.260 ;
        RECT 4.300 470.100 595.700 470.140 ;
        RECT 1.210 468.980 595.700 470.100 ;
        RECT 1.210 465.660 597.430 468.980 ;
        RECT 4.300 464.500 595.700 465.660 ;
        RECT 1.210 461.180 597.430 464.500 ;
        RECT 1.210 460.060 595.700 461.180 ;
        RECT 4.300 460.020 595.700 460.060 ;
        RECT 4.300 458.900 597.430 460.020 ;
        RECT 1.210 456.700 597.430 458.900 ;
        RECT 1.210 455.540 595.700 456.700 ;
        RECT 1.210 454.460 597.430 455.540 ;
        RECT 4.300 453.300 597.430 454.460 ;
        RECT 1.210 452.220 597.430 453.300 ;
        RECT 1.210 451.060 595.700 452.220 ;
        RECT 1.210 448.860 597.430 451.060 ;
        RECT 4.300 447.740 597.430 448.860 ;
        RECT 4.300 447.700 595.700 447.740 ;
        RECT 1.210 446.580 595.700 447.700 ;
        RECT 1.210 443.260 597.430 446.580 ;
        RECT 4.300 442.100 595.700 443.260 ;
        RECT 1.210 438.780 597.430 442.100 ;
        RECT 1.210 437.660 595.700 438.780 ;
        RECT 4.300 437.620 595.700 437.660 ;
        RECT 4.300 436.500 597.430 437.620 ;
        RECT 1.210 434.300 597.430 436.500 ;
        RECT 1.210 433.140 595.700 434.300 ;
        RECT 1.210 432.060 597.430 433.140 ;
        RECT 4.300 430.900 597.430 432.060 ;
        RECT 1.210 429.820 597.430 430.900 ;
        RECT 1.210 428.660 595.700 429.820 ;
        RECT 1.210 426.460 597.430 428.660 ;
        RECT 4.300 425.340 597.430 426.460 ;
        RECT 4.300 425.300 595.700 425.340 ;
        RECT 1.210 424.180 595.700 425.300 ;
        RECT 1.210 420.860 597.430 424.180 ;
        RECT 4.300 419.700 595.700 420.860 ;
        RECT 1.210 416.380 597.430 419.700 ;
        RECT 1.210 415.260 595.700 416.380 ;
        RECT 4.300 415.220 595.700 415.260 ;
        RECT 4.300 414.100 597.430 415.220 ;
        RECT 1.210 411.900 597.430 414.100 ;
        RECT 1.210 410.740 595.700 411.900 ;
        RECT 1.210 409.660 597.430 410.740 ;
        RECT 4.300 408.500 597.430 409.660 ;
        RECT 1.210 407.420 597.430 408.500 ;
        RECT 1.210 406.260 595.700 407.420 ;
        RECT 1.210 404.060 597.430 406.260 ;
        RECT 4.300 402.940 597.430 404.060 ;
        RECT 4.300 402.900 595.700 402.940 ;
        RECT 1.210 401.780 595.700 402.900 ;
        RECT 1.210 398.460 597.430 401.780 ;
        RECT 4.300 397.300 595.700 398.460 ;
        RECT 1.210 393.980 597.430 397.300 ;
        RECT 1.210 392.860 595.700 393.980 ;
        RECT 4.300 392.820 595.700 392.860 ;
        RECT 4.300 391.700 597.430 392.820 ;
        RECT 1.210 389.500 597.430 391.700 ;
        RECT 1.210 388.340 595.700 389.500 ;
        RECT 1.210 387.260 597.430 388.340 ;
        RECT 4.300 386.100 597.430 387.260 ;
        RECT 1.210 385.020 597.430 386.100 ;
        RECT 1.210 383.860 595.700 385.020 ;
        RECT 1.210 381.660 597.430 383.860 ;
        RECT 4.300 380.540 597.430 381.660 ;
        RECT 4.300 380.500 595.700 380.540 ;
        RECT 1.210 379.380 595.700 380.500 ;
        RECT 1.210 376.060 597.430 379.380 ;
        RECT 4.300 374.900 595.700 376.060 ;
        RECT 1.210 371.580 597.430 374.900 ;
        RECT 1.210 370.460 595.700 371.580 ;
        RECT 4.300 370.420 595.700 370.460 ;
        RECT 4.300 369.300 597.430 370.420 ;
        RECT 1.210 367.100 597.430 369.300 ;
        RECT 1.210 365.940 595.700 367.100 ;
        RECT 1.210 364.860 597.430 365.940 ;
        RECT 4.300 363.700 597.430 364.860 ;
        RECT 1.210 362.620 597.430 363.700 ;
        RECT 1.210 361.460 595.700 362.620 ;
        RECT 1.210 359.260 597.430 361.460 ;
        RECT 4.300 358.140 597.430 359.260 ;
        RECT 4.300 358.100 595.700 358.140 ;
        RECT 1.210 356.980 595.700 358.100 ;
        RECT 1.210 353.660 597.430 356.980 ;
        RECT 4.300 352.500 595.700 353.660 ;
        RECT 1.210 349.180 597.430 352.500 ;
        RECT 1.210 348.060 595.700 349.180 ;
        RECT 4.300 348.020 595.700 348.060 ;
        RECT 4.300 346.900 597.430 348.020 ;
        RECT 1.210 344.700 597.430 346.900 ;
        RECT 1.210 343.540 595.700 344.700 ;
        RECT 1.210 342.460 597.430 343.540 ;
        RECT 4.300 341.300 597.430 342.460 ;
        RECT 1.210 340.220 597.430 341.300 ;
        RECT 1.210 339.060 595.700 340.220 ;
        RECT 1.210 336.860 597.430 339.060 ;
        RECT 4.300 335.740 597.430 336.860 ;
        RECT 4.300 335.700 595.700 335.740 ;
        RECT 1.210 334.580 595.700 335.700 ;
        RECT 1.210 331.260 597.430 334.580 ;
        RECT 4.300 330.100 595.700 331.260 ;
        RECT 1.210 326.780 597.430 330.100 ;
        RECT 1.210 325.660 595.700 326.780 ;
        RECT 4.300 325.620 595.700 325.660 ;
        RECT 4.300 324.500 597.430 325.620 ;
        RECT 1.210 322.300 597.430 324.500 ;
        RECT 1.210 321.140 595.700 322.300 ;
        RECT 1.210 320.060 597.430 321.140 ;
        RECT 4.300 318.900 597.430 320.060 ;
        RECT 1.210 317.820 597.430 318.900 ;
        RECT 1.210 316.660 595.700 317.820 ;
        RECT 1.210 314.460 597.430 316.660 ;
        RECT 4.300 313.340 597.430 314.460 ;
        RECT 4.300 313.300 595.700 313.340 ;
        RECT 1.210 312.180 595.700 313.300 ;
        RECT 1.210 308.860 597.430 312.180 ;
        RECT 4.300 307.700 595.700 308.860 ;
        RECT 1.210 304.380 597.430 307.700 ;
        RECT 1.210 303.260 595.700 304.380 ;
        RECT 4.300 303.220 595.700 303.260 ;
        RECT 4.300 302.100 597.430 303.220 ;
        RECT 1.210 299.900 597.430 302.100 ;
        RECT 1.210 298.740 595.700 299.900 ;
        RECT 1.210 297.660 597.430 298.740 ;
        RECT 4.300 296.500 597.430 297.660 ;
        RECT 1.210 295.420 597.430 296.500 ;
        RECT 1.210 294.260 595.700 295.420 ;
        RECT 1.210 292.060 597.430 294.260 ;
        RECT 4.300 290.940 597.430 292.060 ;
        RECT 4.300 290.900 595.700 290.940 ;
        RECT 1.210 289.780 595.700 290.900 ;
        RECT 1.210 286.460 597.430 289.780 ;
        RECT 4.300 285.300 595.700 286.460 ;
        RECT 1.210 281.980 597.430 285.300 ;
        RECT 1.210 280.860 595.700 281.980 ;
        RECT 4.300 280.820 595.700 280.860 ;
        RECT 4.300 279.700 597.430 280.820 ;
        RECT 1.210 277.500 597.430 279.700 ;
        RECT 1.210 276.340 595.700 277.500 ;
        RECT 1.210 275.260 597.430 276.340 ;
        RECT 4.300 274.100 597.430 275.260 ;
        RECT 1.210 273.020 597.430 274.100 ;
        RECT 1.210 271.860 595.700 273.020 ;
        RECT 1.210 269.660 597.430 271.860 ;
        RECT 4.300 268.540 597.430 269.660 ;
        RECT 4.300 268.500 595.700 268.540 ;
        RECT 1.210 267.380 595.700 268.500 ;
        RECT 1.210 264.060 597.430 267.380 ;
        RECT 4.300 262.900 595.700 264.060 ;
        RECT 1.210 259.580 597.430 262.900 ;
        RECT 1.210 258.460 595.700 259.580 ;
        RECT 4.300 258.420 595.700 258.460 ;
        RECT 4.300 257.300 597.430 258.420 ;
        RECT 1.210 255.100 597.430 257.300 ;
        RECT 1.210 253.940 595.700 255.100 ;
        RECT 1.210 252.860 597.430 253.940 ;
        RECT 4.300 251.700 597.430 252.860 ;
        RECT 1.210 250.620 597.430 251.700 ;
        RECT 1.210 249.460 595.700 250.620 ;
        RECT 1.210 247.260 597.430 249.460 ;
        RECT 4.300 246.140 597.430 247.260 ;
        RECT 4.300 246.100 595.700 246.140 ;
        RECT 1.210 244.980 595.700 246.100 ;
        RECT 1.210 241.660 597.430 244.980 ;
        RECT 4.300 240.500 595.700 241.660 ;
        RECT 1.210 237.180 597.430 240.500 ;
        RECT 1.210 236.060 595.700 237.180 ;
        RECT 4.300 236.020 595.700 236.060 ;
        RECT 4.300 234.900 597.430 236.020 ;
        RECT 1.210 232.700 597.430 234.900 ;
        RECT 1.210 231.540 595.700 232.700 ;
        RECT 1.210 230.460 597.430 231.540 ;
        RECT 4.300 229.300 597.430 230.460 ;
        RECT 1.210 228.220 597.430 229.300 ;
        RECT 1.210 227.060 595.700 228.220 ;
        RECT 1.210 224.860 597.430 227.060 ;
        RECT 4.300 223.740 597.430 224.860 ;
        RECT 4.300 223.700 595.700 223.740 ;
        RECT 1.210 222.580 595.700 223.700 ;
        RECT 1.210 219.260 597.430 222.580 ;
        RECT 4.300 218.100 595.700 219.260 ;
        RECT 1.210 214.780 597.430 218.100 ;
        RECT 1.210 213.660 595.700 214.780 ;
        RECT 4.300 213.620 595.700 213.660 ;
        RECT 4.300 212.500 597.430 213.620 ;
        RECT 1.210 210.300 597.430 212.500 ;
        RECT 1.210 209.140 595.700 210.300 ;
        RECT 1.210 208.060 597.430 209.140 ;
        RECT 4.300 206.900 597.430 208.060 ;
        RECT 1.210 205.820 597.430 206.900 ;
        RECT 1.210 204.660 595.700 205.820 ;
        RECT 1.210 202.460 597.430 204.660 ;
        RECT 4.300 201.340 597.430 202.460 ;
        RECT 4.300 201.300 595.700 201.340 ;
        RECT 1.210 200.180 595.700 201.300 ;
        RECT 1.210 196.860 597.430 200.180 ;
        RECT 4.300 195.700 595.700 196.860 ;
        RECT 1.210 192.380 597.430 195.700 ;
        RECT 1.210 191.260 595.700 192.380 ;
        RECT 4.300 191.220 595.700 191.260 ;
        RECT 4.300 190.100 597.430 191.220 ;
        RECT 1.210 187.900 597.430 190.100 ;
        RECT 1.210 186.740 595.700 187.900 ;
        RECT 1.210 185.660 597.430 186.740 ;
        RECT 4.300 184.500 597.430 185.660 ;
        RECT 1.210 183.420 597.430 184.500 ;
        RECT 1.210 182.260 595.700 183.420 ;
        RECT 1.210 180.060 597.430 182.260 ;
        RECT 4.300 178.940 597.430 180.060 ;
        RECT 4.300 178.900 595.700 178.940 ;
        RECT 1.210 177.780 595.700 178.900 ;
        RECT 1.210 174.460 597.430 177.780 ;
        RECT 4.300 173.300 595.700 174.460 ;
        RECT 1.210 169.980 597.430 173.300 ;
        RECT 1.210 168.860 595.700 169.980 ;
        RECT 4.300 168.820 595.700 168.860 ;
        RECT 4.300 167.700 597.430 168.820 ;
        RECT 1.210 165.500 597.430 167.700 ;
        RECT 1.210 164.340 595.700 165.500 ;
        RECT 1.210 163.260 597.430 164.340 ;
        RECT 4.300 162.100 597.430 163.260 ;
        RECT 1.210 161.020 597.430 162.100 ;
        RECT 1.210 159.860 595.700 161.020 ;
        RECT 1.210 157.660 597.430 159.860 ;
        RECT 4.300 156.540 597.430 157.660 ;
        RECT 4.300 156.500 595.700 156.540 ;
        RECT 1.210 155.380 595.700 156.500 ;
        RECT 1.210 152.060 597.430 155.380 ;
        RECT 4.300 150.900 595.700 152.060 ;
        RECT 1.210 147.580 597.430 150.900 ;
        RECT 1.210 146.460 595.700 147.580 ;
        RECT 4.300 146.420 595.700 146.460 ;
        RECT 4.300 145.300 597.430 146.420 ;
        RECT 1.210 143.100 597.430 145.300 ;
        RECT 1.210 141.940 595.700 143.100 ;
        RECT 1.210 140.860 597.430 141.940 ;
        RECT 4.300 139.700 597.430 140.860 ;
        RECT 1.210 138.620 597.430 139.700 ;
        RECT 1.210 137.460 595.700 138.620 ;
        RECT 1.210 135.260 597.430 137.460 ;
        RECT 4.300 134.140 597.430 135.260 ;
        RECT 4.300 134.100 595.700 134.140 ;
        RECT 1.210 132.980 595.700 134.100 ;
        RECT 1.210 129.660 597.430 132.980 ;
        RECT 4.300 128.500 595.700 129.660 ;
        RECT 1.210 125.180 597.430 128.500 ;
        RECT 1.210 124.060 595.700 125.180 ;
        RECT 4.300 124.020 595.700 124.060 ;
        RECT 4.300 122.900 597.430 124.020 ;
        RECT 1.210 120.700 597.430 122.900 ;
        RECT 1.210 119.540 595.700 120.700 ;
        RECT 1.210 118.460 597.430 119.540 ;
        RECT 4.300 117.300 597.430 118.460 ;
        RECT 1.210 116.220 597.430 117.300 ;
        RECT 1.210 115.060 595.700 116.220 ;
        RECT 1.210 112.860 597.430 115.060 ;
        RECT 4.300 111.740 597.430 112.860 ;
        RECT 4.300 111.700 595.700 111.740 ;
        RECT 1.210 110.580 595.700 111.700 ;
        RECT 1.210 107.260 597.430 110.580 ;
        RECT 4.300 106.100 595.700 107.260 ;
        RECT 1.210 102.780 597.430 106.100 ;
        RECT 1.210 101.660 595.700 102.780 ;
        RECT 4.300 101.620 595.700 101.660 ;
        RECT 4.300 100.500 597.430 101.620 ;
        RECT 1.210 98.300 597.430 100.500 ;
        RECT 1.210 97.140 595.700 98.300 ;
        RECT 1.210 96.060 597.430 97.140 ;
        RECT 4.300 94.900 597.430 96.060 ;
        RECT 1.210 93.820 597.430 94.900 ;
        RECT 1.210 92.660 595.700 93.820 ;
        RECT 1.210 90.460 597.430 92.660 ;
        RECT 4.300 89.340 597.430 90.460 ;
        RECT 4.300 89.300 595.700 89.340 ;
        RECT 1.210 88.180 595.700 89.300 ;
        RECT 1.210 84.860 597.430 88.180 ;
        RECT 4.300 83.700 595.700 84.860 ;
        RECT 1.210 80.380 597.430 83.700 ;
        RECT 1.210 79.260 595.700 80.380 ;
        RECT 4.300 79.220 595.700 79.260 ;
        RECT 4.300 78.100 597.430 79.220 ;
        RECT 1.210 75.900 597.430 78.100 ;
        RECT 1.210 74.740 595.700 75.900 ;
        RECT 1.210 73.660 597.430 74.740 ;
        RECT 4.300 72.500 597.430 73.660 ;
        RECT 1.210 71.420 597.430 72.500 ;
        RECT 1.210 70.260 595.700 71.420 ;
        RECT 1.210 68.060 597.430 70.260 ;
        RECT 4.300 66.940 597.430 68.060 ;
        RECT 4.300 66.900 595.700 66.940 ;
        RECT 1.210 65.780 595.700 66.900 ;
        RECT 1.210 62.460 597.430 65.780 ;
        RECT 4.300 61.300 595.700 62.460 ;
        RECT 1.210 57.980 597.430 61.300 ;
        RECT 1.210 56.860 595.700 57.980 ;
        RECT 4.300 56.820 595.700 56.860 ;
        RECT 4.300 55.700 597.430 56.820 ;
        RECT 1.210 53.500 597.430 55.700 ;
        RECT 1.210 52.340 595.700 53.500 ;
        RECT 1.210 51.260 597.430 52.340 ;
        RECT 4.300 50.100 597.430 51.260 ;
        RECT 1.210 49.020 597.430 50.100 ;
        RECT 1.210 47.860 595.700 49.020 ;
        RECT 1.210 45.660 597.430 47.860 ;
        RECT 4.300 44.540 597.430 45.660 ;
        RECT 4.300 44.500 595.700 44.540 ;
        RECT 1.210 43.380 595.700 44.500 ;
        RECT 1.210 40.060 597.430 43.380 ;
        RECT 4.300 38.900 595.700 40.060 ;
        RECT 1.210 13.580 597.430 38.900 ;
      LAYER Metal4 ;
        RECT 10.220 15.080 21.940 577.830 ;
        RECT 24.140 15.080 98.740 577.830 ;
        RECT 100.940 15.080 175.540 577.830 ;
        RECT 177.740 15.080 252.340 577.830 ;
        RECT 254.540 15.080 329.140 577.830 ;
        RECT 331.340 15.080 405.940 577.830 ;
        RECT 408.140 15.080 482.740 577.830 ;
        RECT 484.940 15.080 559.540 577.830 ;
        RECT 561.740 15.080 589.540 577.830 ;
        RECT 10.220 14.090 589.540 15.080 ;
  END
END multiplexer
END LIBRARY

