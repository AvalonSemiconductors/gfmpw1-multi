magic
tech gf180mcuD
magscale 1 5
timestamp 1753964060
<< nwell >>
rect 629 11153 12363 11411
rect 629 10369 12363 10799
rect 629 9585 12363 10015
rect 629 8801 12363 9231
rect 629 8017 12363 8447
rect 629 7233 12363 7663
rect 629 6449 12363 6879
rect 629 5665 12363 6095
rect 629 4881 12363 5311
rect 629 4097 12363 4527
rect 629 3313 12363 3743
rect 629 2529 12363 2959
rect 629 1745 12363 2175
<< pwell >>
rect 629 10799 12363 11153
rect 629 10015 12363 10369
rect 629 9231 12363 9585
rect 629 8447 12363 8801
rect 629 7663 12363 8017
rect 629 6879 12363 7233
rect 629 6095 12363 6449
rect 629 5311 12363 5665
rect 629 4527 12363 4881
rect 629 3743 12363 4097
rect 629 2959 12363 3313
rect 629 2175 12363 2529
rect 629 1525 12363 1745
<< obsm1 >>
rect 672 1538 12400 11465
<< metal2 >>
rect 2128 12600 2184 13000
rect 6384 12600 6440 13000
rect 10640 12600 10696 13000
<< obsm2 >>
rect 798 12570 2098 12600
rect 2214 12570 6354 12600
rect 6470 12570 10610 12600
rect 10726 12570 12530 12600
rect 798 905 12530 12570
<< metal3 >>
rect 12600 11984 13000 12040
rect 12600 10976 13000 11032
rect 12600 9968 13000 10024
rect 12600 8960 13000 9016
rect 12600 7952 13000 8008
rect 12600 6944 13000 7000
rect 12600 5936 13000 5992
rect 12600 4928 13000 4984
rect 12600 3920 13000 3976
rect 12600 2912 13000 2968
rect 12600 1904 13000 1960
rect 12600 896 13000 952
<< obsm3 >>
rect 793 11954 12570 12026
rect 793 11062 12600 11954
rect 793 10946 12570 11062
rect 793 10054 12600 10946
rect 793 9938 12570 10054
rect 793 9046 12600 9938
rect 793 8930 12570 9046
rect 793 8038 12600 8930
rect 793 7922 12570 8038
rect 793 7030 12600 7922
rect 793 6914 12570 7030
rect 793 6022 12600 6914
rect 793 5906 12570 6022
rect 793 5014 12600 5906
rect 793 4898 12570 5014
rect 793 4006 12600 4898
rect 793 3890 12570 4006
rect 793 2998 12600 3890
rect 793 2882 12570 2998
rect 793 1990 12600 2882
rect 793 1874 12570 1990
rect 793 982 12600 1874
rect 793 910 12570 982
<< metal4 >>
rect 2048 1538 2208 11398
rect 3504 1538 3664 11398
rect 4960 1538 5120 11398
rect 6416 1538 6576 11398
rect 7872 1538 8032 11398
rect 9328 1538 9488 11398
rect 10784 1538 10944 11398
rect 12240 1538 12400 11398
<< obsm4 >>
rect 3374 5217 3474 10183
rect 3694 5217 4930 10183
rect 5150 5217 6386 10183
rect 6606 5217 7842 10183
rect 8062 5217 9298 10183
rect 9518 5217 10754 10183
rect 10974 5217 11354 10183
<< labels >>
rlabel metal3 s 12600 896 13000 952 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 12600 10976 13000 11032 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 12600 11984 13000 12040 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 12600 1904 13000 1960 6 custom_settings[1]
port 4 nsew signal input
rlabel metal3 s 12600 2912 13000 2968 6 custom_settings[2]
port 5 nsew signal input
rlabel metal3 s 12600 3920 13000 3976 6 custom_settings[3]
port 6 nsew signal input
rlabel metal3 s 12600 4928 13000 4984 6 custom_settings[4]
port 7 nsew signal input
rlabel metal3 s 12600 5936 13000 5992 6 custom_settings[5]
port 8 nsew signal input
rlabel metal3 s 12600 6944 13000 7000 6 custom_settings[6]
port 9 nsew signal input
rlabel metal3 s 12600 7952 13000 8008 6 custom_settings[7]
port 10 nsew signal input
rlabel metal3 s 12600 8960 13000 9016 6 custom_settings[8]
port 11 nsew signal input
rlabel metal3 s 12600 9968 13000 10024 6 custom_settings[9]
port 12 nsew signal input
rlabel metal2 s 10640 12600 10696 13000 6 io_out
port 13 nsew signal output
rlabel metal2 s 6384 12600 6440 13000 6 rst_n
port 14 nsew signal input
rlabel metal4 s 2048 1538 2208 11398 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 4960 1538 5120 11398 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 7872 1538 8032 11398 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 10784 1538 10944 11398 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 3504 1538 3664 11398 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 6416 1538 6576 11398 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 9328 1538 9488 11398 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 12240 1538 12400 11398 6 vss
port 16 nsew ground bidirectional
rlabel metal2 s 2128 12600 2184 13000 6 wb_clk_i
port 17 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 13000 13000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 572530
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/hellorld/runs/25_07_31_14_13/results/signoff/hellorld.magic.gds
string GDS_START 157828
<< end >>

