magic
tech gf180mcuD
magscale 1 10
timestamp 1700061068
<< nwell >>
rect 1258 41145 44662 41984
rect 1258 41120 32557 41145
rect 1258 40391 27629 40416
rect 1258 39577 44662 40391
rect 1258 39552 29981 39577
rect 1258 38823 27965 38848
rect 1258 38009 44662 38823
rect 1258 37984 33798 38009
rect 1258 36443 44662 37280
rect 1258 36441 17264 36443
rect 1258 36416 9192 36441
rect 1258 35687 21021 35712
rect 1258 34873 44662 35687
rect 1258 34848 9373 34873
rect 1258 34119 14259 34144
rect 1258 34117 19168 34119
rect 1258 33305 44662 34117
rect 1258 33280 8477 33305
rect 1258 32551 7960 32576
rect 1258 32549 12784 32551
rect 1258 31739 44662 32549
rect 1258 31737 25104 31739
rect 1258 31712 8029 31737
rect 1258 30981 12672 31008
rect 1258 30171 44662 30981
rect 1258 30169 25216 30171
rect 1258 30146 15457 30169
rect 1258 30144 14144 30146
rect 1258 29415 7960 29440
rect 1258 28603 44662 29415
rect 1258 28601 26896 28603
rect 1258 28576 8365 28601
rect 1258 27847 13392 27872
rect 1258 27035 44662 27847
rect 1258 27033 26000 27035
rect 1258 27010 17921 27033
rect 1258 27008 16608 27010
rect 1258 26302 10560 26304
rect 1258 26279 11873 26302
rect 1258 25465 44662 26279
rect 1258 25440 9696 25465
rect 1258 24711 10704 24736
rect 1258 24709 20176 24711
rect 1258 23897 44662 24709
rect 1258 23872 15632 23897
rect 1258 23166 11232 23168
rect 1258 23143 12545 23166
rect 1258 22329 44662 23143
rect 1258 22306 8625 22329
rect 1258 22304 7312 22306
rect 1258 21598 4288 21600
rect 1258 21575 5601 21598
rect 1258 20761 44662 21575
rect 1258 20736 8800 20761
rect 1258 20030 2496 20032
rect 1258 20007 3809 20030
rect 1258 20005 37872 20007
rect 1258 19193 44662 20005
rect 1258 19168 16024 19193
rect 1258 18439 1968 18464
rect 1258 17625 44662 18439
rect 1258 17600 6112 17625
rect 1258 16869 6569 16896
rect 1258 16057 44662 16869
rect 1258 16032 25428 16057
rect 1258 15303 10381 15328
rect 1258 14489 44662 15303
rect 1258 14464 9821 14489
rect 1258 13735 11725 13760
rect 1258 13733 37872 13735
rect 1258 12921 44662 13733
rect 1258 12896 15757 12921
rect 1258 12167 14749 12192
rect 1258 11353 44662 12167
rect 1258 11328 18040 11353
rect 1258 10599 20280 10624
rect 1258 9785 44662 10599
rect 1258 9760 10157 9785
rect 1258 9031 11432 9056
rect 1258 8217 44662 9031
rect 1258 8192 16673 8217
rect 1258 7486 11120 7488
rect 1258 7463 12433 7486
rect 1258 6651 44662 7463
rect 1258 6624 10544 6651
rect 1258 5918 13808 5920
rect 1258 5895 15121 5918
rect 1258 5081 44662 5895
rect 1258 5056 11958 5081
rect 1258 4350 12464 4352
rect 1258 4327 13777 4350
rect 1258 3513 44662 4327
rect 1258 3488 14590 3513
<< pwell >>
rect 1258 41984 44662 42422
rect 1258 40416 44662 41120
rect 1258 38848 44662 39552
rect 1258 37280 44662 37984
rect 1258 35712 44662 36416
rect 1258 34144 44662 34848
rect 1258 32576 44662 33280
rect 1258 31008 44662 31712
rect 1258 29440 44662 30144
rect 1258 27872 44662 28576
rect 1258 26304 44662 27008
rect 1258 24736 44662 25440
rect 1258 23168 44662 23872
rect 1258 21600 44662 22304
rect 1258 20032 44662 20736
rect 1258 18464 44662 19168
rect 1258 16896 44662 17600
rect 1258 15328 44662 16032
rect 1258 13760 44662 14464
rect 1258 12192 44662 12896
rect 1258 10624 44662 11328
rect 1258 9056 44662 9760
rect 1258 7488 44662 8192
rect 1258 5920 44662 6624
rect 1258 4352 44662 5056
rect 1258 3050 44662 3488
<< obsm1 >>
rect 1344 3076 44576 42396
<< obsm2 >>
rect 1596 2706 44660 43102
<< metal3 >>
rect 45200 43008 46000 43120
rect 45200 39648 46000 39760
rect 45200 36288 46000 36400
rect 45200 32928 46000 33040
rect 45200 29568 46000 29680
rect 45200 26208 46000 26320
rect 45200 22848 46000 22960
rect 45200 19488 46000 19600
rect 45200 16128 46000 16240
rect 45200 12768 46000 12880
rect 45200 9408 46000 9520
rect 45200 6048 46000 6160
rect 45200 2688 46000 2800
<< obsm3 >>
rect 2034 42948 45140 43092
rect 2034 39820 45332 42948
rect 2034 39588 45140 39820
rect 2034 36460 45332 39588
rect 2034 36228 45140 36460
rect 2034 33100 45332 36228
rect 2034 32868 45140 33100
rect 2034 29740 45332 32868
rect 2034 29508 45140 29740
rect 2034 26380 45332 29508
rect 2034 26148 45140 26380
rect 2034 23020 45332 26148
rect 2034 22788 45140 23020
rect 2034 19660 45332 22788
rect 2034 19428 45140 19660
rect 2034 16300 45332 19428
rect 2034 16068 45140 16300
rect 2034 12940 45332 16068
rect 2034 12708 45140 12940
rect 2034 9580 45332 12708
rect 2034 9348 45140 9580
rect 2034 6220 45332 9348
rect 2034 5988 45140 6220
rect 2034 2860 45332 5988
rect 2034 2716 45140 2860
<< metal4 >>
rect 4448 3076 4768 42396
rect 19808 3076 20128 42396
rect 35168 3076 35488 42396
<< obsm4 >>
rect 18844 6066 19748 42094
rect 20188 6066 35108 42094
rect 35548 6066 36372 42094
<< labels >>
rlabel metal3 s 45200 2688 46000 2800 6 clk
port 1 nsew signal input
rlabel metal3 s 45200 9408 46000 9520 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 45200 12768 46000 12880 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 45200 16128 46000 16240 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 45200 19488 46000 19600 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 45200 22848 46000 22960 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 45200 26208 46000 26320 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 45200 29568 46000 29680 6 io_out[0]
port 8 nsew signal output
rlabel metal3 s 45200 32928 46000 33040 6 io_out[1]
port 9 nsew signal output
rlabel metal3 s 45200 36288 46000 36400 6 io_out[2]
port 10 nsew signal output
rlabel metal3 s 45200 39648 46000 39760 6 io_out[3]
port 11 nsew signal output
rlabel metal3 s 45200 43008 46000 43120 6 io_out[4]
port 12 nsew signal output
rlabel metal3 s 45200 6048 46000 6160 6 rst_n
port 13 nsew signal input
rlabel metal4 s 4448 3076 4768 42396 6 vdd
port 14 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 42396 6 vdd
port 14 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 42396 6 vss
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 46000 46000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1392682
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/tbb1143/runs/23_11_15_16_07/results/signoff/tholin_avalonsemi_tbb1143.magic.gds
string GDS_START 255134
<< end >>

