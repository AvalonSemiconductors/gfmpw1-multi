* NGSPICE file created from multiplexer.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt multiplexer ay8913_do[0] ay8913_do[10] ay8913_do[11] ay8913_do[12] ay8913_do[13]
+ ay8913_do[14] ay8913_do[15] ay8913_do[16] ay8913_do[17] ay8913_do[18] ay8913_do[19]
+ ay8913_do[1] ay8913_do[20] ay8913_do[21] ay8913_do[22] ay8913_do[23] ay8913_do[24]
+ ay8913_do[25] ay8913_do[26] ay8913_do[27] ay8913_do[2] ay8913_do[3] ay8913_do[4]
+ ay8913_do[5] ay8913_do[6] ay8913_do[7] ay8913_do[8] ay8913_do[9] blinker_do[0] blinker_do[1]
+ blinker_do[2] custom_settings[0] custom_settings[10] custom_settings[11] custom_settings[12]
+ custom_settings[13] custom_settings[14] custom_settings[15] custom_settings[16]
+ custom_settings[17] custom_settings[18] custom_settings[19] custom_settings[1] custom_settings[20]
+ custom_settings[21] custom_settings[22] custom_settings[23] custom_settings[24]
+ custom_settings[25] custom_settings[26] custom_settings[27] custom_settings[28]
+ custom_settings[29] custom_settings[2] custom_settings[30] custom_settings[31] custom_settings[3]
+ custom_settings[4] custom_settings[5] custom_settings[6] custom_settings[7] custom_settings[8]
+ custom_settings[9] diceroll_do[0] diceroll_do[1] diceroll_do[2] diceroll_do[3] diceroll_do[4]
+ diceroll_do[5] diceroll_do[6] diceroll_do[7] diceroll_do[8] hellorld_do io_in_0
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16]
+ io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30]
+ io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] mc14500_do[0] mc14500_do[10] mc14500_do[11]
+ mc14500_do[12] mc14500_do[13] mc14500_do[14] mc14500_do[15] mc14500_do[16] mc14500_do[17]
+ mc14500_do[18] mc14500_do[19] mc14500_do[1] mc14500_do[20] mc14500_do[21] mc14500_do[22]
+ mc14500_do[23] mc14500_do[24] mc14500_do[25] mc14500_do[26] mc14500_do[27] mc14500_do[28]
+ mc14500_do[29] mc14500_do[2] mc14500_do[30] mc14500_do[3] mc14500_do[4] mc14500_do[5]
+ mc14500_do[6] mc14500_do[7] mc14500_do[8] mc14500_do[9] mc14500_sram_addr[0] mc14500_sram_addr[1]
+ mc14500_sram_addr[2] mc14500_sram_addr[3] mc14500_sram_addr[4] mc14500_sram_addr[5]
+ mc14500_sram_gwe mc14500_sram_in[0] mc14500_sram_in[1] mc14500_sram_in[2] mc14500_sram_in[3]
+ mc14500_sram_in[4] mc14500_sram_in[5] mc14500_sram_in[6] mc14500_sram_in[7] pdp11_do[0]
+ pdp11_do[10] pdp11_do[11] pdp11_do[12] pdp11_do[13] pdp11_do[14] pdp11_do[15] pdp11_do[16]
+ pdp11_do[17] pdp11_do[18] pdp11_do[19] pdp11_do[1] pdp11_do[20] pdp11_do[21] pdp11_do[22]
+ pdp11_do[23] pdp11_do[24] pdp11_do[25] pdp11_do[26] pdp11_do[27] pdp11_do[28] pdp11_do[29]
+ pdp11_do[2] pdp11_do[30] pdp11_do[31] pdp11_do[32] pdp11_do[3] pdp11_do[4] pdp11_do[5]
+ pdp11_do[6] pdp11_do[7] pdp11_do[8] pdp11_do[9] pdp11_oeb[0] pdp11_oeb[10] pdp11_oeb[11]
+ pdp11_oeb[12] pdp11_oeb[13] pdp11_oeb[14] pdp11_oeb[15] pdp11_oeb[16] pdp11_oeb[17]
+ pdp11_oeb[18] pdp11_oeb[19] pdp11_oeb[1] pdp11_oeb[20] pdp11_oeb[21] pdp11_oeb[22]
+ pdp11_oeb[23] pdp11_oeb[24] pdp11_oeb[25] pdp11_oeb[26] pdp11_oeb[27] pdp11_oeb[28]
+ pdp11_oeb[29] pdp11_oeb[2] pdp11_oeb[30] pdp11_oeb[31] pdp11_oeb[32] pdp11_oeb[3]
+ pdp11_oeb[4] pdp11_oeb[5] pdp11_oeb[6] pdp11_oeb[7] pdp11_oeb[8] pdp11_oeb[9] qcpu_do[0]
+ qcpu_do[10] qcpu_do[11] qcpu_do[12] qcpu_do[13] qcpu_do[14] qcpu_do[15] qcpu_do[16]
+ qcpu_do[17] qcpu_do[18] qcpu_do[19] qcpu_do[1] qcpu_do[20] qcpu_do[21] qcpu_do[22]
+ qcpu_do[23] qcpu_do[24] qcpu_do[25] qcpu_do[26] qcpu_do[27] qcpu_do[28] qcpu_do[29]
+ qcpu_do[2] qcpu_do[30] qcpu_do[31] qcpu_do[32] qcpu_do[3] qcpu_do[4] qcpu_do[5]
+ qcpu_do[6] qcpu_do[7] qcpu_do[8] qcpu_do[9] qcpu_oeb[0] qcpu_oeb[10] qcpu_oeb[11]
+ qcpu_oeb[12] qcpu_oeb[13] qcpu_oeb[14] qcpu_oeb[15] qcpu_oeb[16] qcpu_oeb[17] qcpu_oeb[18]
+ qcpu_oeb[19] qcpu_oeb[1] qcpu_oeb[20] qcpu_oeb[21] qcpu_oeb[22] qcpu_oeb[23] qcpu_oeb[24]
+ qcpu_oeb[25] qcpu_oeb[26] qcpu_oeb[27] qcpu_oeb[28] qcpu_oeb[29] qcpu_oeb[2] qcpu_oeb[30]
+ qcpu_oeb[31] qcpu_oeb[32] qcpu_oeb[3] qcpu_oeb[4] qcpu_oeb[5] qcpu_oeb[6] qcpu_oeb[7]
+ qcpu_oeb[8] qcpu_oeb[9] qcpu_sram_addr[0] qcpu_sram_addr[1] qcpu_sram_addr[2] qcpu_sram_addr[3]
+ qcpu_sram_addr[4] qcpu_sram_addr[5] qcpu_sram_gwe qcpu_sram_in[0] qcpu_sram_in[1]
+ qcpu_sram_in[2] qcpu_sram_in[3] qcpu_sram_in[4] qcpu_sram_in[5] qcpu_sram_in[6]
+ qcpu_sram_in[7] qcpu_sram_out[0] qcpu_sram_out[1] qcpu_sram_out[2] qcpu_sram_out[3]
+ qcpu_sram_out[4] qcpu_sram_out[5] qcpu_sram_out[6] qcpu_sram_out[7] rst_ay8913 rst_blinker
+ rst_diceroll rst_hellorld rst_mc14500 rst_pdp11 rst_qcpu rst_sid rst_sn76489 rst_tbb1143
+ rst_tholin_riscv rst_ue1 sid_do[0] sid_do[10] sid_do[11] sid_do[12] sid_do[13] sid_do[14]
+ sid_do[15] sid_do[16] sid_do[17] sid_do[18] sid_do[19] sid_do[1] sid_do[20] sid_do[2]
+ sid_do[3] sid_do[4] sid_do[5] sid_do[6] sid_do[7] sid_do[8] sid_do[9] sid_oeb sn76489_do[0]
+ sn76489_do[10] sn76489_do[11] sn76489_do[12] sn76489_do[13] sn76489_do[14] sn76489_do[15]
+ sn76489_do[16] sn76489_do[17] sn76489_do[18] sn76489_do[19] sn76489_do[1] sn76489_do[20]
+ sn76489_do[21] sn76489_do[22] sn76489_do[23] sn76489_do[24] sn76489_do[25] sn76489_do[26]
+ sn76489_do[27] sn76489_do[2] sn76489_do[3] sn76489_do[4] sn76489_do[5] sn76489_do[6]
+ sn76489_do[7] sn76489_do[8] sn76489_do[9] tbb1143_do[0] tbb1143_do[1] tbb1143_do[2]
+ tbb1143_do[3] tbb1143_do[4] tholin_riscv_do[0] tholin_riscv_do[10] tholin_riscv_do[11]
+ tholin_riscv_do[12] tholin_riscv_do[13] tholin_riscv_do[14] tholin_riscv_do[15]
+ tholin_riscv_do[16] tholin_riscv_do[17] tholin_riscv_do[18] tholin_riscv_do[19]
+ tholin_riscv_do[1] tholin_riscv_do[20] tholin_riscv_do[21] tholin_riscv_do[22] tholin_riscv_do[23]
+ tholin_riscv_do[24] tholin_riscv_do[25] tholin_riscv_do[26] tholin_riscv_do[27]
+ tholin_riscv_do[28] tholin_riscv_do[29] tholin_riscv_do[2] tholin_riscv_do[30] tholin_riscv_do[31]
+ tholin_riscv_do[32] tholin_riscv_do[3] tholin_riscv_do[4] tholin_riscv_do[5] tholin_riscv_do[6]
+ tholin_riscv_do[7] tholin_riscv_do[8] tholin_riscv_do[9] tholin_riscv_oeb[0] tholin_riscv_oeb[10]
+ tholin_riscv_oeb[11] tholin_riscv_oeb[12] tholin_riscv_oeb[13] tholin_riscv_oeb[14]
+ tholin_riscv_oeb[15] tholin_riscv_oeb[16] tholin_riscv_oeb[17] tholin_riscv_oeb[18]
+ tholin_riscv_oeb[19] tholin_riscv_oeb[1] tholin_riscv_oeb[20] tholin_riscv_oeb[21]
+ tholin_riscv_oeb[22] tholin_riscv_oeb[23] tholin_riscv_oeb[24] tholin_riscv_oeb[25]
+ tholin_riscv_oeb[26] tholin_riscv_oeb[27] tholin_riscv_oeb[28] tholin_riscv_oeb[29]
+ tholin_riscv_oeb[2] tholin_riscv_oeb[30] tholin_riscv_oeb[31] tholin_riscv_oeb[32]
+ tholin_riscv_oeb[3] tholin_riscv_oeb[4] tholin_riscv_oeb[5] tholin_riscv_oeb[6]
+ tholin_riscv_oeb[7] tholin_riscv_oeb[8] tholin_riscv_oeb[9] ue1_do[0] ue1_do[1]
+ ue1_do[2] ue1_do[3] ue1_do[4] ue1_do[5] ue1_do[6] ue1_do[7] ue1_do[8] ue1_do[9]
+ ue1_oeb vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_stb_i wbs_we_i irq[2] irq[1] irq[0]
XFILLER_0_94_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3155_ _1582_ _1616_ _1619_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5968__A1 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3086_ _1459_ _1570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5512__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input108_I pdp11_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5196__A2 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ _2177_ _2170_ _2178_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5727_ _1187_ _1200_ net469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_60_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ net189 _1144_ _1149_ net123 net325 _1146_ _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input73_I mc14500_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5589_ _0662_ _1090_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_115_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4609_ _2625_ _2626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_92_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5120__A2 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3131__A1 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5111__A2 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_143_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_125_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3869__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4474__B _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4960_ dffram.data\[42\]\[7\] _2906_ _2910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4622__A1 net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ dffram.data\[51\]\[5\] _2126_ _2128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ wb_counter\[22\] _2855_ _2860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3842_ dffram.data\[52\]\[1\] _2077_ _2079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6630_ _0550_ clknet_leaf_117_wb_clk_i wb_counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6561_ _0481_ clknet_leaf_133_wb_clk_i design_select\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3773_ _1838_ _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5512_ dffram.data\[32\]\[6\] dffram.data\[34\]\[6\] dffram.data\[36\]\[6\] dffram.data\[38\]\[6\]
+ _0758_ _0760_ _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4925__A2 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6492_ _0412_ clknet_leaf_81_wb_clk_i dffram.data\[45\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5443_ dffram.data\[32\]\[4\] dffram.data\[34\]\[4\] dffram.data\[36\]\[4\] dffram.data\[38\]\[4\]
+ _0758_ _0760_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5525__S _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _0721_ _0870_ _0881_ _0755_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xoutput434 net434 custom_settings[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput423 net423 custom_settings[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput467 net467 io_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput478 net478 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_35_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput456 net456 io_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4325_ _2355_ _2394_ _2397_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput445 net445 custom_settings[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput489 net489 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4256_ dffram.data\[16\]\[4\] _2353_ _2354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5260__S _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3207_ dffram.data\[62\]\[5\] _1653_ _1656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4187_ _2301_ _2309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3138_ _1558_ _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input225_I qcpu_sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmultiplexer_569 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3069_ _1501_ _1550_ _1555_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3019__I _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5435__S _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output444_I net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5234__I _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_47_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_166_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3343__A1 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4110_ _2225_ _2253_ _2257_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5090_ dffram.data\[9\]\[5\] _2992_ _2994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4041_ _2167_ _2206_ _2211_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_56_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ net227 _1428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4943_ _2898_ _2900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6613_ _0533_ clknet_leaf_128_wb_clk_i wb_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4874_ _2411_ _2846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3825_ _2035_ _2062_ _2067_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__I _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _0464_ clknet_leaf_122_wb_clk_i net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3756_ dffram.data\[23\]\[4\] _2021_ _2022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3582__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _0395_ clknet_leaf_83_wb_clk_i dffram.data\[46\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_65_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5426_ _0929_ _0932_ _0846_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3687_ _1965_ _1977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input175_I qcpu_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _0757_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input342_I tholin_riscv_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5288_ _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4308_ _2359_ _2381_ _2386_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input36_I diceroll_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4239_ _1921_ _2265_ _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_74_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5229__I _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_83_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output561_I net561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_92_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _1905_ _1923_ _1926_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5553__A2 _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__I _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _2427_ _2555_ _2608_ _2609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3541_ _1872_ _1879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3472_ _1829_ _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6260_ _0180_ clknet_leaf_30_wb_clk_i dffram.data\[57\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6191_ _0111_ clknet_leaf_102_wb_clk_i dffram.data\[31\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5142_ _0648_ _0657_ net523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_62_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5073_ dffram.data\[39\]\[7\] _2979_ _2983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4024_ _2169_ _2199_ _2201_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4218__I _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1387_ _1414_ _1415_ net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA_clkbuf_4_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4926_ _2850_ _2886_ _2887_ _2846_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4857_ _2821_ _2831_ _2832_ _2829_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_43_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input292_I tholin_riscv_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3808_ _2037_ _2055_ _2057_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_60_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4788_ _2760_ _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _0447_ clknet_leaf_136_wb_clk_i dffram.data\[17\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3739_ dffram.data\[54\]\[7\] _2006_ _2010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6458_ _0378_ clknet_leaf_60_wb_clk_i dffram.data\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5409_ dffram.data\[49\]\[3\] dffram.data\[51\]\[3\] dffram.data\[53\]\[3\] dffram.data\[55\]\[3\]
+ _0816_ _0817_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6389_ _0309_ clknet_leaf_138_wb_clk_i dffram.data\[19\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_89_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4807__A1 net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3794__A1 _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3546__A1 _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3877__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _1214_ _1220_ _1228_ net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5691_ _1145_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4711_ _2692_ _2713_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4642_ _2615_ _2655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_135_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _0962_ _0981_ _2568_ _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3524_ dffram.data\[26\]\[5\] _1867_ _1869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6312_ _0232_ clknet_leaf_1_wb_clk_i dffram.data\[55\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3455_ dffram.data\[5\]\[1\] _1818_ _1820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6243_ _0163_ clknet_leaf_36_wb_clk_i dffram.data\[58\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3386_ dffram.data\[28\]\[1\] _1772_ _1775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6174_ _0094_ clknet_leaf_5_wb_clk_i dffram.data\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5125_ design_select\[4\] design_select\[1\] _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA_input138_I pdp11_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5056_ _2971_ _2973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ _2175_ _2186_ _2190_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input305_I tholin_riscv_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5958_ net274 _1278_ _1370_ net59 net307 _1357_ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_75_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4909_ _2796_ _2872_ _2874_ _2875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5889_ _1237_ _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3528__A1 dffram.data\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3027__I _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput312 tholin_riscv_do[29] net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput301 tholin_riscv_do[19] net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput345 tholin_riscv_oeb[29] net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput334 tholin_riscv_oeb[19] net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput323 tholin_riscv_do[9] net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output524_I net524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold41 net581 net618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold30 _2438_ net607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput356 tholin_riscv_oeb[9] net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput367 ue1_oeb net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold52 wbs_adr_i[17] net634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold74 net668 net651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput378 wbs_adr_i[7] net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput389 net609 net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold96 wbs_dat_i[9] net674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold85 wbs_adr_i[19] net663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5300__S1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6006__C _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_85_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3519__A1 _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__I _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_5 _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4321__I _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3240_ _1676_ _1678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5580__C _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__B2 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A1 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5152__I _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3171_ dffram.data\[63\]\[3\] _1626_ _1630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _1274_ _1238_ _1275_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5743_ _1087_ _1207_ _1211_ _1212_ net473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_137_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5528__S _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5674_ _1113_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5327__I _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _1523_ _2640_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4183__A1 _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4556_ _2566_ wb_counter\[2\] _2576_ _2578_ _2559_ _2579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_130_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3507_ _1856_ _1846_ _1857_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _2131_ _1858_ _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6226_ _0146_ clknet_leaf_42_wb_clk_i dffram.data\[60\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3438_ dffram.data\[60\]\[3\] _1805_ _1809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input255_I sid_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5683__B2 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A1 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _0077_ clknet_leaf_88_wb_clk_i dffram.data\[33\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3369_ _1756_ _1763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _0629_ wb_override_act _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6088_ _0008_ clknet_leaf_78_wb_clk_i dffram.data\[35\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5986__A2 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5039_ _2942_ _2959_ _2962_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5530__S1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3749__A1 _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output474_I net474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5237__I _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput120 pdp11_do[8] net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_132_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_132_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_133_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput142 pdp11_oeb[28] net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput131 pdp11_oeb[18] net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput153 pdp11_oeb[8] net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput175 qcpu_do[28] net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput186 qcpu_do[8] net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput164 qcpu_do[18] net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5977__A2 _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput197 qcpu_oeb[18] net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3988__A1 _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__S _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _2461_ net631 _2457_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_10_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _0777_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3912__A1 _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _1521_ _2411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_169_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4272_ dffram.data\[18\]\[1\] _2363_ _2365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3223_ _1645_ _1664_ _1667_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6011_ dffram.data\[36\]\[0\] _1446_ _1447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3154_ dffram.data\[0\]\[5\] _1617_ _1619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4935__B _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3085_ _1568_ _1564_ _1569_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A1 _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3987_ dffram.data\[50\]\[7\] _2171_ _2178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5726_ net208 _1197_ _1183_ net142 net344 _1198_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ _1123_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4156__A1 _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input66_I mc14500_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5588_ _0655_ _0661_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4608_ _2624_ _2625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_92_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4539_ _2545_ _2560_ _2563_ _2564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4896__I _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5656__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _0129_ clknet_leaf_68_wb_clk_i dffram.data\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5120__A3 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4136__I _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__B _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5895__A1 net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5647__A1 net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5430__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4622__A2 _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_103_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5258__S0 _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3910_ _2104_ _2125_ _2127_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _2858_ _2859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5586__B _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3841_ _2026_ _2076_ _2078_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3772_ _2031_ _2028_ _2032_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4386__A1 net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _0480_ clknet_leaf_116_wb_clk_i net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_144_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5511_ dffram.data\[40\]\[6\] dffram.data\[42\]\[6\] dffram.data\[44\]\[6\] dffram.data\[46\]\[6\]
+ _0807_ _0808_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_113_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _0411_ clknet_leaf_81_wb_clk_i dffram.data\[45\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A1 _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5442_ dffram.data\[40\]\[4\] dffram.data\[42\]\[4\] dffram.data\[44\]\[4\] dffram.data\[46\]\[4\]
+ _0865_ _0866_ _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__5886__B2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5373_ _0876_ _0880_ _0749_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput435 net435 custom_settings[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput424 net424 custom_settings[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput468 net468 io_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput446 net446 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_35_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput457 net457 io_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4324_ dffram.data\[17\]\[5\] _2395_ _2397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput479 net479 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5489__I1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4255_ _2341_ _2353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3206_ _1581_ _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4186_ _2301_ _2308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3137_ _1588_ _1602_ _1607_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input120_I pdp11_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input218_I qcpu_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5810__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3068_ dffram.data\[43\]\[7\] _1551_ _1555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5810__B2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3795__I _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ net202 _1174_ _1178_ net136 net338 _1175_ _1189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_94_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6689_ _0609_ clknet_leaf_92_wb_clk_i dffram.data\[39\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5877__A1 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__B2 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__S0 _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output437_I net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5488__S0 _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5361__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4040_ dffram.data\[4\]\[3\] _2207_ _2211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4485__B _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1426_ _0829_ _1427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _2898_ _2899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6612_ _0532_ clknet_leaf_131_wb_clk_i wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4873_ _2841_ _2843_ _2845_ _2829_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_166_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3824_ dffram.data\[22\]\[3\] _2063_ _2067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3031__A1 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5536__S _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ _0463_ clknet_leaf_124_wb_clk_i net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3755_ _2013_ _2021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6474_ _0394_ clknet_leaf_83_wb_clk_i dffram.data\[46\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3686_ _1965_ _1976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5859__A1 net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5425_ _0930_ _0931_ _0893_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5335__I _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ _0861_ _0862_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input168_I qcpu_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _0681_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4307_ dffram.data\[44\]\[7\] _2382_ _2386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input335_I tholin_riscv_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _1444_ _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input29_I blinker_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ dffram.data\[15\]\[6\] _2292_ _2297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3022__A1 _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3089__A1 _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3013__A1 _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3540_ _1842_ _1873_ _1878_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5356__S _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4761__A1 _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3471_ _1443_ _1829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5210_ _0715_ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _0110_ clknet_leaf_102_wb_clk_i dffram.data\[31\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5141_ _0653_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4994__I _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _2954_ _2978_ _2982_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4023_ dffram.data\[49\]\[4\] _2200_ _2201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5974_ net63 _1218_ _1116_ net109 net311 _1118_ _1415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_87_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3252__A1 _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ net403 _2776_ _2887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ net387 _2824_ _2832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3807_ dffram.data\[13\]\[4\] _2056_ _2057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input285_I sn76489_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4787_ _2762_ _2774_ _2775_ _2769_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6526_ _0446_ clknet_leaf_136_wb_clk_i dffram.data\[17\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3738_ _1981_ _2005_ _2009_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6457_ _0377_ clknet_leaf_62_wb_clk_i dffram.data\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5065__I _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3669_ _1423_ _0961_ _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_140_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5701__B1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6388_ _0308_ clknet_leaf_59_wb_clk_i dffram.data\[19\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5408_ _0910_ _0913_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4504__A1 dffram.data\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0677_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_89_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4991__A1 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold37_I wbs_dat_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__B1 _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _1162_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_139_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4054__I _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4710_ net547 _2697_ _2698_ _2712_ _2713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _2653_ wb_counter\[12\] _2654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4572_ wb_counter\[4\] _2593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3523_ _1845_ _1866_ _1868_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6311_ _0231_ clknet_leaf_2_wb_clk_i dffram.data\[55\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3454_ _1769_ _1817_ _1819_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6242_ _0162_ clknet_leaf_42_wb_clk_i dffram.data\[58\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3385_ _1567_ _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6173_ _0093_ clknet_leaf_5_wb_clk_i dffram.data\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ design_select\[3\] _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5055_ _2971_ _2972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4229__I _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ dffram.data\[29\]\[6\] _2187_ _2190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input200_I qcpu_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5957_ net171 _1249_ _1334_ net105 _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3225__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4908_ _2721_ _2859_ _2873_ _2874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_36_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input96_I pdp11_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _1115_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4839_ _2646_ wb_counter\[12\] _2809_ _2818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_71_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6509_ _0429_ clknet_leaf_104_wb_clk_i dffram.data\[18\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput302 tholin_riscv_do[1] net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold7_I wbs_dat_i[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput335 tholin_riscv_oeb[1] net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput324 tholin_riscv_oeb[0] net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput313 tholin_riscv_do[2] net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold20 net626 net597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold31 wbs_dat_i[11] net611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput346 tholin_riscv_oeb[2] net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput357 ue1_do[0] net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_output517_I net517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold64 net614 net641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 net617 net630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput368 wb_rst_i net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold42 _2442_ net619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput379 net655 net379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold75 net667 net652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold86 wbs_dat_i[5] net664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold97 wbs_dat_i[1] net675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3464__A1 _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3218__I _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_6 _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5677__C1 net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _1571_ _1625_ _1629_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ net251 _1215_ _1255_ net116 _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5742_ net147 _1156_ _1106_ net349 _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_57_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4955__A1 _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ _1160_ _1161_ net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4624_ net564 _2623_ _2626_ _2639_ _2640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_167_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _1140_ _2556_ _2577_ _2578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3506_ dffram.data\[58\]\[7\] _1847_ _1857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3128__I _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4486_ _1444_ _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input150_I pdp11_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3437_ _1776_ _1804_ _1808_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6225_ _0145_ clknet_leaf_43_wb_clk_i dffram.data\[60\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5132__A1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _0076_ clknet_leaf_77_wb_clk_i dffram.data\[33\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3368_ _1712_ _1757_ _1762_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input248_I sid_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5107_ wb_rst_override _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6087_ _0007_ clknet_leaf_91_wb_clk_i dffram.data\[36\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3299_ dffram.data\[32\]\[4\] _1716_ _1717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input11_I ay8913_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5038_ dffram.data\[38\]\[1\] _2960_ _2962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output467_I net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__S _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 pdp11_do[29] net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput143 pdp11_oeb[29] net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput132 pdp11_oeb[19] net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput154 pdp11_oeb[9] net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput121 pdp11_do[9] net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_158_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput176 qcpu_do[29] net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput165 qcpu_do[19] net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput187 qcpu_do[9] net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__3437__A1 _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput198 qcpu_oeb[19] net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_167_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4340_ net380 _2409_ _2410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_169_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4271_ _2340_ _2362_ _2364_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3222_ dffram.data\[33\]\[1\] _1665_ _1667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6010_ _1435_ _1446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input3_I ay8913_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3153_ _1577_ _1616_ _1618_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3084_ dffram.data\[7\]\[1\] _1565_ _1569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3428__A1 _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3986_ _2114_ _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _1187_ _1199_ net468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_31_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _0670_ _1142_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_128_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input198_I qcpu_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4607_ net372 _2540_ _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input365_I ue1_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ net257 _1086_ _1088_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_103_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4538_ wb_override_act _2562_ _2563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input59_I mc14500_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ net372 _2507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_106_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6208_ _0128_ clknet_leaf_6_wb_clk_i dffram.data\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3667__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5801__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6139_ _0059_ clknet_leaf_33_wb_clk_i dffram.data\[63\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4417__I _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__S _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3991__I _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5647__A2 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3830__A1 dffram.data\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5586__C _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__S1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3840_ dffram.data\[52\]\[0\] _2077_ _2078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3771_ dffram.data\[53\]\[1\] _2029_ _2032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5510_ _1012_ _1013_ _0811_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6490_ _0410_ clknet_leaf_82_wb_clk_i dffram.data\[45\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5441_ _0945_ _0946_ _0863_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5372_ _0877_ _0878_ _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput425 net425 custom_settings[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput414 net414 custom_settings[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput469 net469 io_oeb[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput436 net436 custom_settings[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput447 net447 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput458 net458 io_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4323_ _2351_ _2394_ _2396_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5638__A2 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4254_ _2341_ _2352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5621__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ _2288_ _2302_ _2307_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3205_ _1651_ _1652_ _1654_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3136_ dffram.data\[8\]\[7\] _1603_ _1607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _1494_ _1550_ _1554_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input113_I pdp11_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5777__B _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3141__I _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4074__A1 _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3821__A1 _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5708_ _1187_ _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3969_ _2097_ _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_94_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6688_ _0608_ clknet_leaf_92_wb_clk_i dffram.data\[39\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5639_ _1123_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5877__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__S1 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__S0 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__I _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__S1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3051__I _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3812__A1 _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_120_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__I _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5990_ _0827_ _1426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _2300_ _1885_ _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ net390 _2844_ _2845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3823_ _2033_ _2062_ _2066_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _0531_ clknet_leaf_131_wb_clk_i wb_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_31_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6542_ _0462_ clknet_leaf_122_wb_clk_i net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3754_ _2013_ _2020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ _0393_ clknet_leaf_82_wb_clk_i dffram.data\[46\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3685_ _1844_ _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5424_ dffram.data\[16\]\[3\] dffram.data\[18\]\[3\] dffram.data\[20\]\[3\] dffram.data\[22\]\[3\]
+ _0841_ _0842_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4520__I _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5355_ _0810_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ _0794_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4306_ _2357_ _2381_ _2385_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4237_ _2298_ _2334_ _2339_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input328_I tholin_riscv_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input230_I qcpu_sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4168_ _2111_ _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3119_ _1595_ _1597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4047__A1 _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ _2235_ _2246_ _2250_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3046__I _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__B _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__A1 dffram.data\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_79_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5786__A1 net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__B2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A1 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ _1788_ _1823_ _1828_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__S _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5140_ _0655_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ dffram.data\[39\]\[6\] _2979_ _2982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5171__I _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ _2192_ _2200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ net175 _1413_ _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_149_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4924_ wb_counter\[30\] _2885_ _2886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ wb_counter\[16\] _2830_ _2831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3806_ _2048_ _2056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4786_ net405 _2764_ _2775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_60_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6525_ _0445_ clknet_leaf_136_wb_clk_i dffram.data\[17\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ dffram.data\[54\]\[6\] _2006_ _2009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input180_I qcpu_do[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input278_I sn76489_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5388__S0 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3668_ _1829_ _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6456_ _0376_ clknet_leaf_106_wb_clk_i dffram.data\[47\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5701__B2 net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _0307_ clknet_leaf_59_wb_clk_i dffram.data\[19\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5407_ _0813_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3599_ _1917_ _1912_ _1918_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5338_ _0837_ _0845_ _0846_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input41_I hellorld_do vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5269_ dffram.data\[1\]\[0\] dffram.data\[3\]\[0\] dffram.data\[5\]\[0\] dffram.data\[7\]\[0\]
+ _0776_ _0778_ _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__S0 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4440__A1 net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output497_I net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_22_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5940__A1 net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__S0 _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__B1 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3504__I _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A1 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5759__B2 net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _2608_ _2653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5166__I _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _2541_ _2592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6310_ _0230_ clknet_leaf_2_wb_clk_i dffram.data\[55\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3522_ dffram.data\[26\]\[4\] _1867_ _1868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3453_ dffram.data\[5\]\[0\] _1818_ _1819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _0161_ clknet_leaf_42_wb_clk_i dffram.data\[58\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _0092_ clknet_leaf_35_wb_clk_i dffram.data\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3384_ _1769_ _1771_ _1773_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3170__A1 _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ design_select\[2\] _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_97_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _1703_ _1562_ _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4005_ _2173_ _2186_ _2189_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3473__A2 _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__A1 net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5956_ net17 _1400_ _1401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4422__A1 net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ net241 _1247_ _1233_ net48 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ wb_counter\[25\] wb_counter\[26\] _2873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_168_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4838_ _2802_ _2816_ _2817_ _2814_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input89_I pdp11_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5922__B2 net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__I _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4769_ _2760_ _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6508_ _0428_ clknet_leaf_61_wb_clk_i dffram.data\[18\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _0359_ clknet_leaf_9_wb_clk_i dffram.data\[48\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput303 tholin_riscv_do[20] net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput336 tholin_riscv_oeb[20] net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput325 tholin_riscv_oeb[10] net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput314 tholin_riscv_do[30] net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3324__I _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold32 net666 net609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold10 wbs_dat_i[22] net590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold21 _2474_ net598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput358 ue1_do[1] net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput347 tholin_riscv_oeb[30] net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5533__S0 _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold54 _2462_ net631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 wbs_dat_i[21] net626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold65 net634 net642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput369 net654 net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold87 wbs_dat_i[6] net665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold76 net675 net653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_168_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_7 _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A2 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_94_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_23_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5524__S0 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5810_ net68 _1254_ _1252_ net35 _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_123_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ net213 _1210_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ net192 _1144_ _1149_ net126 net328 _1146_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3409__I _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4623_ _2636_ _2638_ _2639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4554_ _2547_ _2577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3505_ _1855_ _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6224_ _0144_ clknet_leaf_96_wb_clk_i dffram.data\[34\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4485_ _2517_ _2518_ _2501_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3436_ dffram.data\[60\]\[2\] _1805_ _1808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3143__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5132__A2 net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _0075_ clknet_leaf_77_wb_clk_i dffram.data\[33\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3367_ dffram.data\[2\]\[3\] _1758_ _1762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input143_I pdp11_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6086_ _0006_ clknet_leaf_92_wb_clk_i dffram.data\[36\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5515__S0 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5037_ _2937_ _2959_ _2961_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3298_ _1704_ _1716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input310_I tholin_riscv_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__B1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__A1 net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5939_ _1386_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_119_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput100 pdp11_do[1] net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput111 pdp11_do[2] net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput144 pdp11_oeb[2] net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput133 pdp11_oeb[1] net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput122 pdp11_oeb[0] net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4882__A1 net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput155 qcpu_do[0] net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput177 qcpu_do[2] net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput166 qcpu_do[1] net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4594__B _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__B1 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput199 qcpu_oeb[1] net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput188 qcpu_oeb[0] net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4634__A1 net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_141_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_141_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold97_I wbs_dat_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4937__A2 _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3229__I _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5114__A2 _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4270_ dffram.data\[18\]\[0\] _2363_ _2364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3221_ _1637_ _1664_ _1666_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3125__A1 _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__S _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3152_ dffram.data\[0\]\[4\] _1617_ _1618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3083_ _1567_ _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4625__A1 _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5425__I0 _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ _2175_ _2170_ _2176_ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ net207 _1197_ _1193_ net141 net343 _1198_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_128_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _1142_ _1147_ net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _2582_ _2623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5586_ _0638_ _1087_ _0641_ _0650_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3364__A1 _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input260_I sn76489_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4537_ _2561_ _2562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input358_I ue1_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4468_ _0620_ _2505_ _2506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3419_ _1790_ _1797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6207_ _0127_ clknet_leaf_16_wb_clk_i dffram.data\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ _0058_ clknet_leaf_31_wb_clk_i dffram.data\[63\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4399_ net420 _2447_ _2454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6069_ _1496_ _1440_ _1497_ _1437_ _1498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4616__A1 net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_153_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A1 _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A2 net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3355__A1 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3107__A1 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__A1 net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__I _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5032__A1 _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3770_ _1835_ _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5440_ dffram.data\[33\]\[4\] dffram.data\[35\]\[4\] dffram.data\[37\]\[4\] dffram.data\[39\]\[4\]
+ _0804_ _0805_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _0746_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput426 net426 custom_settings[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput415 net415 custom_settings[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput437 net437 custom_settings[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput448 net448 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4322_ dffram.data\[17\]\[4\] _2395_ _2396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput459 net459 io_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4253_ _1478_ _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3204_ dffram.data\[62\]\[4\] _1653_ _1654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4184_ dffram.data\[46\]\[3\] _2303_ _2307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3135_ _1585_ _1602_ _1606_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3066_ dffram.data\[43\]\[6\] _1551_ _1554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input106_I pdp11_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5023__A1 _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ _2163_ _2160_ _2164_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5707_ _0672_ _1186_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_128_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3585__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3899_ dffram.data\[51\]\[0\] _2120_ _2121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6687_ _0607_ clknet_leaf_92_wb_clk_i dffram.data\[39\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5638_ _1120_ _1134_ net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_116_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input71_I mc14500_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5569_ _1057_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__S1 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4837__A1 net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__C1 net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__B _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_14_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4828__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4940_ _2897_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5005__A1 _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _2780_ _2844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3822_ dffram.data\[22\]\[2\] _2063_ _2066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6610_ _0530_ clknet_leaf_134_wb_clk_i wb_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _0461_ clknet_leaf_124_wb_clk_i net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3753_ _1973_ _2014_ _2019_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3684_ _1973_ _1966_ _1974_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6472_ _0392_ clknet_leaf_56_wb_clk_i dffram.data\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5713__C1 net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ dffram.data\[24\]\[3\] dffram.data\[26\]\[3\] dffram.data\[28\]\[3\] dffram.data\[30\]\[3\]
+ _0889_ _0890_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__3319__A1 _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ dffram.data\[33\]\[2\] dffram.data\[35\]\[2\] dffram.data\[37\]\[2\] dffram.data\[39\]\[2\]
+ _0799_ _0800_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ dffram.data\[44\]\[6\] _2382_ _2385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_34_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _0676_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ dffram.data\[45\]\[7\] _2335_ _2339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4167_ _2294_ _2291_ _2295_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3118_ _1595_ _1596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input223_I qcpu_sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4098_ dffram.data\[14\]\[6\] _2247_ _2250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3049_ _1507_ _1542_ _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3558__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_142_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_52_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_148_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output442_I net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3730__A1 _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_70_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5070_ _2952_ _2978_ _2981_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4021_ _2192_ _2199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4068__I _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _1365_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5777__A2 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3700__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4923_ wb_counter\[28\] wb_counter\[29\] _2879_ _2885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_87_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _2664_ _2671_ _2822_ _2830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_166_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3805_ _2048_ _2055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4785_ wb_counter\[3\] _2773_ _2774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6524_ _0444_ clknet_leaf_93_wb_clk_i dffram.data\[17\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ _1979_ _2005_ _2008_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5388__S1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3667_ _1919_ _1956_ _1961_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6455_ _0375_ clknet_leaf_107_wb_clk_i dffram.data\[47\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input173_I qcpu_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6386_ _0306_ clknet_leaf_58_wb_clk_i dffram.data\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5406_ _0911_ _0912_ _0811_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3598_ dffram.data\[25\]\[6\] _1913_ _1918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5337_ _0813_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input340_I tholin_riscv_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5268_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input34_I diceroll_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4219_ _2327_ _2329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5199_ _0694_ _0699_ _0708_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_104_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__S1 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5379__S1 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__S _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3703__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3520__I _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4195__A1 _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ net559 _2583_ _2591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4351__I _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3521_ _1859_ _1867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3452_ _1816_ _1818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _0160_ clknet_leaf_15_wb_clk_i dffram.data\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3383_ dffram.data\[28\]\[0\] _1772_ _1773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6171_ _0091_ clknet_leaf_34_wb_clk_i dffram.data\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5182__I _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _0632_ _0641_ net528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5053_ _2956_ _2965_ _2970_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4004_ dffram.data\[29\]\[5\] _2187_ _2189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3430__I _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5955_ _1225_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_9_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5886_ net160 _1262_ _1326_ net6 _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_118_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ wb_counter\[25\] _2868_ wb_counter\[26\] _2872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4837_ net383 _2804_ _2817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input290_I tbb1143_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__A2 _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4768_ _2759_ _2760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _0427_ clknet_leaf_61_wb_clk_i dffram.data\[18\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4699_ _2692_ _2703_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3719_ _1983_ _1992_ _1997_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6438_ _0358_ clknet_leaf_146_wb_clk_i dffram.data\[48\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__I _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6369_ _0289_ clknet_leaf_55_wb_clk_i dffram.data\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput326 tholin_riscv_oeb[11] net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput315 tholin_riscv_do[31] net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput304 tholin_riscv_do[21] net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold11 net611 net588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold22 wbs_dat_i[24] net602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput359 ue1_do[2] net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput348 tholin_riscv_oeb[31] net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput337 tholin_riscv_oeb[21] net337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5533__S1 _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold55 net671 net632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold44 net663 net621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold33 _2464_ net610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4110__A1 _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold66 net640 net643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 wbs_adr_i[16] net654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold88 wbs_dat_i[18] net666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_86_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5461__I1 dffram.data\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__I _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5374__B1 _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3924__A1 _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_8 _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5677__A1 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__B2 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5524__S1 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4101__A1 _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3250__I _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5740_ _1121_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_130_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5671_ _1159_ _1092_ _1160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_84_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ net445 _2616_ _2637_ _2638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4553_ _0882_ _0907_ _2568_ _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3504_ _1499_ _1855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4484_ net408 _2510_ _2518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3435_ _1774_ _1804_ _1807_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6223_ _0143_ clknet_leaf_94_wb_clk_i dffram.data\[34\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5132__A3 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6154_ _0074_ clknet_leaf_77_wb_clk_i dffram.data\[33\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3366_ _1710_ _1757_ _1761_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_55_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4340__A1 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5105_ _0620_ _0626_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_100_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _0005_ clknet_leaf_91_wb_clk_i dffram.data\[36\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3297_ _1704_ _1715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input136_I pdp11_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ dffram.data\[38\]\[0\] _2960_ _2961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5515__S1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__B2 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A1 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input303_I tholin_riscv_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5938_ _1237_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5869_ _1139_ _1326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5087__I _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3906__A1 _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput101 pdp11_do[20] net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput112 pdp11_do[30] net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput134 pdp11_oeb[20] net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput123 pdp11_oeb[10] net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput145 pdp11_oeb[30] net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output522_I net522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput156 qcpu_do[10] net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput167 qcpu_do[20] net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput178 qcpu_do[30] net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5831__A1 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput189 qcpu_oeb[10] net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4634__A2 _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__B2 net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3070__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__I1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5898__A1 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_110_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5442__S0 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4570__A1 net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_169_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_120_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3220_ dffram.data\[33\]\[0\] _1665_ _1666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _1609_ _1617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3082_ _1451_ _1567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ dffram.data\[50\]\[6\] _2171_ _2176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5723_ _1126_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5654_ net220 _1144_ _1135_ net154 net356 _1146_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__5189__I0 _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_99_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4605_ _2613_ _2542_ _2620_ _2622_ _1522_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_143_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5585_ _0622_ _0625_ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4536_ _2507_ _2561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _2504_ _2505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3418_ _1778_ _1791_ _1796_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4313__A1 _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input253_I sid_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _0126_ clknet_leaf_11_wb_clk_i dffram.data\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4398_ _2452_ net583 _2446_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6137_ _0057_ clknet_leaf_31_wb_clk_i dffram.data\[63\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3349_ _1714_ _1748_ _1750_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ net409 _1204_ _1497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_29_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _1478_ _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5592__A3 _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5424__S0 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output472_I net472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__A1 net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4304__A1 _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5804__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__B2 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3043__A1 _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5370_ dffram.data\[48\]\[2\] dffram.data\[50\]\[2\] dffram.data\[52\]\[2\] dffram.data\[54\]\[2\]
+ _0742_ _0744_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput416 net416 custom_settings[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput438 net438 custom_settings[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput427 net427 custom_settings[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4321_ _2387_ _2395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput449 net449 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_129_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _2349_ _2342_ _2350_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3203_ _1641_ _1653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4183_ _2286_ _2302_ _2306_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3134_ dffram.data\[8\]\[6\] _1603_ _1606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3065_ _1487_ _1550_ _1553_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3967_ dffram.data\[50\]\[1\] _2161_ _2164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_132_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1091_ _1185_ _1186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__A1 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3898_ _2118_ _2120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6686_ _0606_ clknet_leaf_92_wb_clk_i dffram.data\[39\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ net216 _1131_ _1124_ net150 net352 _1133_ _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input64_I mc14500_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ dffram.data\[0\]\[7\] dffram.data\[2\]\[7\] dffram.data\[4\]\[7\] dffram.data\[6\]\[7\]
+ _1058_ _1059_ _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_44_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4519_ _2541_ _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5499_ dffram.data\[9\]\[5\] dffram.data\[11\]\[5\] dffram.data\[13\]\[5\] dffram.data\[15\]\[5\]
+ _0776_ _0778_ _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3273__A1 _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__A1 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5970__C2 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5275__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ wb_counter\[19\] _2842_ _2843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3821_ _2031_ _2062_ _2065_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5005__A2 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__S _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ _0460_ clknet_leaf_123_wb_clk_i net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5961__B1 _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ dffram.data\[23\]\[3\] _2015_ _2019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3683_ dffram.data\[55\]\[3\] _1967_ _1974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _0391_ clknet_leaf_14_wb_clk_i dffram.data\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5422_ _0927_ _0928_ _0836_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ dffram.data\[41\]\[2\] dffram.data\[43\]\[2\] dffram.data\[45\]\[2\] dffram.data\[47\]\[2\]
+ _0859_ _0860_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _2355_ _2381_ _2384_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5284_ _0756_ _0793_ net512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_26_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4235_ _2296_ _2334_ _2338_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4166_ dffram.data\[15\]\[5\] _2292_ _2295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3117_ _1591_ _1594_ _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input216_I qcpu_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A2 _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4097_ _2233_ _2246_ _2249_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3048_ _1541_ _1542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3007__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4999_ _2534_ _2931_ _2934_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__A1 _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5952__B1 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6669_ _0589_ clknet_leaf_66_wb_clk_i dffram.data\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output435_I net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3246__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5640__C1 net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A1 net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_88_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_17_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4349__I net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4020_ _2167_ _2193_ _2198_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3485__A1 _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1386_ _1410_ _1411_ _1412_ net501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__3237__A1 _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4922_ _2850_ _2883_ _2884_ _2871_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_142_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _2821_ _2827_ _2828_ _2829_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5934__B1 _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _2035_ _2049_ _2054_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4784_ wb_counter\[0\] _2567_ wb_counter\[2\] _2773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _0443_ clknet_leaf_61_wb_clk_i dffram.data\[17\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3735_ dffram.data\[54\]\[5\] _2006_ _2008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _0374_ clknet_leaf_115_wb_clk_i dffram.data\[47\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__C1 net336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ dffram.data\[32\]\[3\] dffram.data\[34\]\[3\] dffram.data\[36\]\[3\] dffram.data\[38\]\[3\]
+ _0807_ _0808_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3666_ dffram.data\[24\]\[7\] _1957_ _1961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6385_ _0305_ clknet_leaf_58_wb_clk_i dffram.data\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3597_ _1852_ _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5336_ _0840_ _0843_ _0844_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input166_I qcpu_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__I _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _0725_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input333_I tholin_riscv_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4218_ _2327_ _2328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input27_I ay8913_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5198_ _0707_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_3_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4149_ dffram.data\[15\]\[0\] _2282_ _2283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4976__A1 _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_124_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_115_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5456__A2 _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__C1 net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_135_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3520_ _1859_ _1866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3451_ _1816_ _1817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3382_ _1770_ _1772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ _0090_ clknet_leaf_35_wb_clk_i dffram.data\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _0637_ _0638_ _0640_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_23_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3458__A1 _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ dffram.data\[38\]\[7\] _2966_ _2970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4003_ _2169_ _2186_ _2188_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3711__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _1396_ _1397_ _1398_ _1399_ net497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_75_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ net365 _1111_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3630__A1 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _2864_ _2869_ _2870_ _2871_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_146_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ wb_counter\[12\] _2815_ _2816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6506_ _0426_ clknet_leaf_61_wb_clk_i dffram.data\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5574__S _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input283_I sn76489_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _2507_ net371 _2401_ _2503_ _2759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_160_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4698_ net545 _2697_ _2698_ _2702_ _2703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3718_ dffram.data\[12\]\[7\] _1993_ _1997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _1949_ _1951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6437_ _0357_ clknet_leaf_146_wb_clk_i dffram.data\[48\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6368_ _0288_ clknet_leaf_8_wb_clk_i dffram.data\[52\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5319_ _0743_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput327 tholin_riscv_oeb[12] net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput316 tholin_riscv_do[32] net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput305 tholin_riscv_do[22] net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6299_ _0219_ clknet_leaf_66_wb_clk_i dffram.data\[24\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold12 _2445_ net589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold23 net674 net600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput349 tholin_riscv_oeb[32] net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput338 tholin_riscv_oeb[22] net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3449__A1 _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold34 wbs_dat_i[23] net614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold45 _2795_ net622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold56 _2496_ net633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold67 net608 net644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold89 wbs_dat_i[3] net667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold78 wbs_cyc_i net655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_168_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_119_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4949__A1 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_9 _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5126__A1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_128_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3531__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__A1 _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3612__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5670_ _0640_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4621_ _2631_ _2637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ net555 _2542_ _2575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3503_ _1853_ _1846_ _1854_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5193__I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4483_ _0639_ _2512_ _2517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3434_ dffram.data\[60\]\[1\] _1805_ _1807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6222_ _0142_ clknet_leaf_97_wb_clk_i dffram.data\[34\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ _0073_ clknet_leaf_77_wb_clk_i dffram.data\[33\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3365_ dffram.data\[2\]\[2\] _1758_ _1761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _0622_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6084_ _0004_ clknet_leaf_91_wb_clk_i dffram.data\[36\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3296_ _1576_ _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5035_ _2958_ _2960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3441__I _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input129_I pdp11_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3851__A1 _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5937_ _1381_ _1385_ net494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_76_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input94_I pdp11_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5868_ _1261_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5799_ net67 _1264_ _1181_ net317 _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_91_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _2776_ _2802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_151_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_112_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3616__I _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 pdp11_do[21] net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 pdp11_do[31] net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput135 pdp11_oeb[21] net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput124 pdp11_oeb[11] net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput146 pdp11_oeb[31] net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output515_I net515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput168 qcpu_do[21] net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput157 qcpu_do[11] net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput179 qcpu_do[31] net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4095__A1 _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__S _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__I _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5442__S1 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_169_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3150_ _1609_ _1616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3081_ _1557_ _1564_ _1566_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__I _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_145_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3261__I _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3833__A1 _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1162_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_128_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3983_ _2111_ _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4092__I _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5653_ _1145_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5584_ _0635_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4010__A1 _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4604_ _2621_ wb_counter\[7\] _2592_ _2559_ _2622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4535_ _2548_ _2549_ _2554_ _2558_ _2559_ _2560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_29_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _2502_ _2401_ _2503_ _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3417_ dffram.data\[34\]\[3\] _1792_ _1796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5361__I1 _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6205_ _0125_ clknet_leaf_11_wb_clk_i dffram.data\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4397_ net385 _2444_ _2453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input246_I sid_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ dffram.data\[30\]\[4\] _1749_ _1750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6136_ _0056_ clknet_leaf_6_wb_clk_i dffram.data\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_163_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6066__A2 _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _1659_ _1696_ _1701_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6067_ net88 _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_29_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A1 _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input413_I wbs_we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _2946_ _2939_ _2947_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3824__A1 dffram.data\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5424__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output465_I net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3346__I _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5188__S0 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_129_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4177__I _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_164_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5360__S0 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3815__A1 _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4640__I _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput417 net417 custom_settings[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput428 net428 custom_settings[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4320_ _2387_ _2394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput439 net439 custom_settings[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4251_ dffram.data\[16\]\[3\] _2343_ _2350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3202_ _1641_ _1652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input1_I ay8913_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4182_ dffram.data\[46\]\[2\] _2303_ _2306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3133_ _1582_ _1602_ _1605_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3064_ dffram.data\[43\]\[5\] _1551_ _1553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3282__A2 _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3966_ _2094_ _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__A1 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5705_ _1159_ _0654_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6685_ _0605_ clknet_leaf_74_wb_clk_i dffram.data\[39\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_34_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5636_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5646__I net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input196_I qcpu_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _2118_ _2119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4550__I _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5567_ _0844_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input363_I ue1_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5498_ _0999_ _1002_ _0814_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4518_ net533 _2542_ _2543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input57_I mc14500_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _2488_ net636 _2491_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6039__A2 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6119_ _0039_ clknet_leaf_18_wb_clk_i dffram.data\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__S0 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3025__A2 _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__A1 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__B2 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__I _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5291__I _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__B2 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A1 net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ dffram.data\[22\]\[1\] _2063_ _2065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _1971_ _2014_ _2018_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5961__A1 net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3682_ _1841_ _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6470_ _0390_ clknet_leaf_13_wb_clk_i dffram.data\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__B2 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5713__A1 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ dffram.data\[25\]\[3\] dffram.data\[27\]\[3\] dffram.data\[29\]\[3\] dffram.data\[31\]\[3\]
+ _0832_ _0834_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _0796_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_26_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ dffram.data\[44\]\[5\] _2382_ _2384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5283_ _0771_ _0774_ _0790_ _0792_ _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_103_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ dffram.data\[45\]\[6\] _2335_ _2338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5572__S0 _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4165_ _2108_ _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3116_ _1593_ _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4096_ dffram.data\[14\]\[5\] _2247_ _2249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input111_I pdp11_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3047_ _1540_ _0720_ _1541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4452__A1 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input209_I qcpu_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4204__A1 _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_82_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4998_ dffram.data\[40\]\[5\] _2932_ _2934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5952__A1 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3949_ _2101_ _2146_ _2151_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5376__I _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _0588_ clknet_leaf_66_wb_clk_i dffram.data\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5619_ _1109_ _1112_ _1119_ net475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__5704__A1 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6599_ _0519_ clknet_leaf_119_wb_clk_i net550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_148_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3191__A1 _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6000__I _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__S0 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output428_I net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4443__A1 net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3182__A1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4682__A1 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ net277 _1322_ _1206_ net62 net310 _1366_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__5482__I0 _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4921_ net401 _2776_ _2884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_47_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4852_ _2768_ _2829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3803_ dffram.data\[13\]\[3\] _2050_ _2054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5934__B2 net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__A1 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _2762_ _2771_ _2772_ _2769_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_160_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _0442_ clknet_leaf_93_wb_clk_i dffram.data\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ _1975_ _2005_ _2007_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3665_ _1917_ _1956_ _1960_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6453_ _0373_ clknet_leaf_113_wb_clk_i dffram.data\[47\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ dffram.data\[40\]\[3\] dffram.data\[42\]\[3\] dffram.data\[44\]\[3\] dffram.data\[46\]\[3\]
+ _0865_ _0866_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6384_ _0304_ clknet_leaf_4_wb_clk_i dffram.data\[51\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3596_ _1915_ _1912_ _1916_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5335_ _0691_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5266_ _0677_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5545__S0 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input159_I qcpu_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4217_ _2047_ _1542_ _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input326_I tholin_riscv_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5197_ _0706_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4148_ _2280_ _2282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_67_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4425__A1 net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4079_ dffram.data\[48\]\[7\] _2231_ _2238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5925__A1 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5861__B1 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__C2 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A1 net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_104_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _1526_ _1559_ _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3155__A1 _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3381_ _1770_ _1771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ _0639_ _0623_ _0624_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_62_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__S0 _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5051_ _2954_ _2965_ _2969_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4002_ dffram.data\[29\]\[4\] _2187_ _2188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4655__A1 net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5953_ net273 _1278_ _1370_ net58 net306 _1357_ _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_1_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ _1285_ _1333_ _1335_ _1339_ net487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_75_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _2411_ _2871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5907__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5907__B2 net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4835_ _2646_ _2809_ _2815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4766_ _2754_ _2402_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6505_ _0425_ clknet_leaf_61_wb_clk_i dffram.data\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_99_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4591__B1 _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3717_ _1981_ _1992_ _1996_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _2699_ _2700_ _2701_ _2702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5135__A2 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3648_ _1949_ _1950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _0356_ clknet_leaf_53_wb_clk_i dffram.data\[48\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input276_I sn76489_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3579_ _1899_ _1902_ _1904_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3174__I _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6367_ _0287_ clknet_leaf_1_wb_clk_i dffram.data\[52\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5318_ _0826_ _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4894__A1 net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput306 tholin_riscv_do[23] net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput317 tholin_riscv_do[3] net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6298_ _0218_ clknet_leaf_69_wb_clk_i dffram.data\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5518__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold13 wbs_dat_i[16] net593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput339 tholin_riscv_oeb[23] net339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput328 tholin_riscv_oeb[13] net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5249_ _0681_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold35 net590 net612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold46 wbs_adr_i[18] net623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold24 _2440_ net601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold68 net602 net645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold57 wbs_dat_i[31] net637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold79 _1524_ net656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_98_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output495_I net495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_156_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5374__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__B1 _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5126__A2 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3137__A1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold28_I wbs_dat_i[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3860__A2 _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5062__A1 _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _2621_ wb_counter\[9\] _2636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3376__A1 _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_72_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _2565_ _2573_ _2574_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ dffram.data\[58\]\[6\] _1847_ _1854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4482_ _0660_ _2505_ _2516_ _2514_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3433_ _1769_ _1804_ _1806_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6221_ _0141_ clknet_leaf_97_wb_clk_i dffram.data\[34\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6152_ _0072_ clknet_leaf_17_wb_clk_i dffram.data\[62\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5103_ _0623_ _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3364_ _1708_ _1757_ _1760_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_55_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _1712_ _1705_ _1713_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6083_ _0003_ clknet_leaf_74_wb_clk_i dffram.data\[36\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3722__I _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5034_ _2958_ _2959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3300__A1 _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5053__A1 _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5936_ net13 _1362_ _1363_ _1384_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5867_ _1319_ _1324_ net485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_63_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5798_ _1217_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input87_I mc14500_sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _2799_ _2801_ _2605_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _2734_ _2745_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6419_ _0339_ clknet_leaf_32_wb_clk_i dffram.data\[49\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4867__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput114 pdp11_do[32] net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput136 pdp11_oeb[22] net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput103 pdp11_do[22] net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput125 pdp11_oeb[12] net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4619__A1 _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput147 pdp11_oeb[32] net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput158 qcpu_do[12] net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput169 qcpu_do[22] net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output508_I net508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__I _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3079__I _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3358__A1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3542__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__I _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__B1 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3080_ dffram.data\[7\]\[0\] _1565_ _1566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3982_ _2173_ _2170_ _2174_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5721_ _1187_ _1196_ net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_85_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5652_ _1125_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3349__A1 _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5583_ _1085_ net519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4603_ _2608_ _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4534_ _2502_ _2559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_57_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4849__A1 _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4465_ wb_feedback_delay _1524_ _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3416_ _1776_ _1791_ _1795_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6204_ _0124_ clknet_leaf_37_wb_clk_i dffram.data\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4396_ net419 _2447_ _2452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3452__I _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3347_ _1741_ _1749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6135_ _0055_ clknet_leaf_6_wb_clk_i dffram.data\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input141_I pdp11_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input239_I sid_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ _1472_ _1494_ _1495_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ dffram.data\[3\]\[3\] _2940_ _2947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3278_ dffram.data\[6\]\[7\] _1697_ _1701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A1 _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3588__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5919_ _1217_ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_119_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3627__I _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3760__A1 dffram.data\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5188__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output458_I net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__S1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A2 _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3579__A1 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold95_I wbs_dat_i[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3751__A1 _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput429 net429 custom_settings[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput418 net418 custom_settings[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4250_ _1469_ _2349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_35_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4181_ _2284_ _2302_ _2305_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3503__A1 _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3201_ _1576_ _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_52_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__I _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3132_ dffram.data\[8\]\[5\] _1603_ _1605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3063_ _1479_ _1550_ _1552_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3965_ _2158_ _2160_ _2162_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5704_ _0670_ _0672_ _1182_ _1184_ net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6684_ _0604_ clknet_leaf_75_wb_clk_i dffram.data\[39\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3896_ _1507_ _2117_ _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5635_ _1125_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5716__C1 net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input189_I qcpu_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ dffram.data\[8\]\[7\] dffram.data\[10\]\[7\] dffram.data\[12\]\[7\] dffram.data\[14\]\[7\]
+ _1058_ _1059_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__5662__I _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5497_ _1000_ _1001_ _0893_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4517_ _2541_ _2542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input356_I tholin_riscv_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4448_ _2468_ _2491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4278__I _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_146_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4379_ net411 _2432_ _2440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6118_ _0038_ clknet_leaf_17_wb_clk_i dffram.data\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5342__S1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ dffram.data\[36\]\[4\] _1480_ _1481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_107_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_87_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5270__I1 _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__I2 dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_129_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_129_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold10_I wbs_dat_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4461__A2 _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5747__I _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3750_ dffram.data\[23\]\[2\] _2015_ _2018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5961__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3681_ _1971_ _1966_ _1972_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5420_ dffram.data\[17\]\[3\] dffram.data\[19\]\[3\] dffram.data\[21\]\[3\] dffram.data\[23\]\[3\]
+ _0884_ _0885_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5351_ _0794_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3724__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5282_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4302_ _2351_ _2381_ _2383_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4233_ _2294_ _2334_ _2337_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5572__S1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _2290_ _2291_ _2293_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3115_ _1592_ _1432_ _1593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4095_ _2229_ _2246_ _2248_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3046_ _0844_ _1540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input104_I pdp11_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4997_ _2530_ _2931_ _2933_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__I _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5952__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3948_ dffram.data\[59\]\[3\] _2147_ _2151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6667_ _0587_ clknet_leaf_67_wb_clk_i dffram.data\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3879_ _2090_ _2105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5618_ net199 _1114_ _1116_ net133 net335 _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _0518_ clknet_leaf_118_wb_clk_i net549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5549_ dffram.data\[49\]\[7\] dffram.data\[51\]\[7\] dffram.data\[53\]\[7\] dffram.data\[55\]\[7\]
+ _0975_ _0976_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3715__A1 _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5563__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4140__A1 _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5640__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__B2 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5995__C net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_30_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_26_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ wb_counter\[29\] _2882_ _2883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ net386 _2824_ _2828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3802_ _2033_ _2049_ _2053_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4782_ net402 _2764_ _2772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3945__A1 _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _0441_ clknet_leaf_94_wb_clk_i dffram.data\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_60_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ dffram.data\[54\]\[4\] _2006_ _2007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _0372_ clknet_leaf_82_wb_clk_i dffram.data\[47\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3664_ dffram.data\[24\]\[6\] _1957_ _1960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5698__B2 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5698__A1 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5403_ _0908_ _0909_ _0863_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6383_ _0303_ clknet_leaf_4_wb_clk_i dffram.data\[51\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3595_ dffram.data\[25\]\[5\] _1913_ _1916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4370__A1 net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5334_ dffram.data\[16\]\[1\] dffram.data\[18\]\[1\] dffram.data\[20\]\[1\] dffram.data\[22\]\[1\]
+ _0841_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5265_ dffram.data\[9\]\[0\] dffram.data\[11\]\[0\] dffram.data\[13\]\[0\] dffram.data\[15\]\[0\]
+ _0696_ _0697_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_103_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5545__S1 _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4216_ _2298_ _2321_ _2326_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5196_ _0702_ _0705_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4122__A1 _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5170__I0 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__A1 net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__B2 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4147_ _2280_ _2281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input221_I qcpu_sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input319_I tholin_riscv_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4078_ _2114_ _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_168_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3029_ _1445_ _1528_ _1530_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_84_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A1 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5481__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3936__A1 _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4361__A1 net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output440_I net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__B2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3370__I _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__S _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5916__A2 _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_144_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_144_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3380_ _1434_ _1726_ _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_21_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5050_ dffram.data\[38\]\[6\] _2966_ _2969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5527__S1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6077__B _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4001_ _2179_ _2187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_141_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ net170 _1249_ _1334_ net104 _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_149_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ net397 _2866_ _2870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ net364 _1098_ _1338_ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_146_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5907__A2 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4834_ _2802_ _2812_ _2813_ _2814_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_28_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3918__A1 _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4765_ _2754_ _2758_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6504_ _0424_ clknet_leaf_106_wb_clk_i dffram.data\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3716_ dffram.data\[12\]\[6\] _1993_ _1996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ net426 _2665_ _2672_ _2701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6435_ _0355_ clknet_leaf_52_wb_clk_i dffram.data\[48\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _1921_ _1858_ _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input171_I qcpu_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3578_ dffram.data\[25\]\[0\] _1903_ _1904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input269_I sn76489_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _0286_ clknet_leaf_1_wb_clk_i dffram.data\[52\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5317_ _0722_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput307 tholin_riscv_do[24] net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput318 tholin_riscv_do[4] net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6297_ _0217_ clknet_leaf_65_wb_clk_i dffram.data\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5518__S1 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold14 net599 net591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_41_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput329 tholin_riscv_oeb[14] net329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input32_I diceroll_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5248_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold47 net661 net624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold25 wbs_dat_i[19] net605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold36 _2476_ net613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold58 net673 net635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 net665 net646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5179_ _0688_ _0673_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_168_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output488_I net488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4334__A1 net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_5_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5834__A1 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__B2 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4550_ _2419_ _2574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3501_ _1852_ _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4481_ net407 _2504_ _2516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6220_ _0140_ clknet_leaf_69_wb_clk_i dffram.data\[34\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3432_ dffram.data\[60\]\[0\] _1805_ _1806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5373__I0 _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__B1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4325__A1 _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_41_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3363_ dffram.data\[2\]\[1\] _1758_ _1760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6151_ _0071_ clknet_leaf_19_wb_clk_i dffram.data\[62\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5102_ design_select\[2\] _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5825__A1 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6082_ _0002_ clknet_leaf_76_wb_clk_i dffram.data\[36\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3294_ dffram.data\[32\]\[3\] _1706_ _1713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__B2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5033_ _1703_ _1740_ _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_36_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5935_ _1382_ _1383_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5866_ _1257_ _1320_ _1321_ _1323_ _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ net410 _2800_ _2801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5665__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5797_ net279 _1260_ _1262_ net181 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_91_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4748_ net553 _2739_ _2740_ _2744_ _2745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4679_ _2608_ _2686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_112_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6418_ _0338_ clknet_leaf_29_wb_clk_i dffram.data\[49\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_112_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6349_ _0269_ clknet_leaf_141_wb_clk_i dffram.data\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6069__A1 _1496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput104 pdp11_do[23] net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput126 pdp11_oeb[13] net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput115 pdp11_do[3] net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 pdp11_oeb[23] net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput148 pdp11_oeb[3] net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput159 qcpu_do[13] net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_99_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3055__A1 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__S0 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3358__A2 _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4555__A1 _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold40_I wbs_dat_i[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3530__A2 _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5807__B2 net318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5807__A1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_59_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3981_ dffram.data\[50\]\[5\] _2171_ _2174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5720_ net206 _1190_ _1193_ net140 net342 _1191_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_85_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4794__A1 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5651_ _1121_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5582_ _1065_ _1084_ _1085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ net443 _2616_ net519 _2617_ _2619_ _2620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_143_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4533_ _2400_ _2556_ _2557_ _2558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_68_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_57_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6203_ _0123_ clknet_leaf_38_wb_clk_i dffram.data\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4464_ net372 _2502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3415_ dffram.data\[34\]\[2\] _1792_ _1795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4395_ _2450_ net595 _2446_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3346_ _1741_ _1748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6134_ _0054_ clknet_leaf_5_wb_clk_i dffram.data\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6065_ dffram.data\[36\]\[6\] _1480_ _1495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input134_I pdp11_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5016_ _1469_ _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3277_ _1657_ _1696_ _1700_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_77_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input301_I tholin_riscv_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5918_ _1361_ _1369_ net491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_64_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__S0 _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5849_ net28 _1266_ _1252_ net40 _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__I _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3908__I _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_86_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_168_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output520_I net520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4776__A1 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold88_I wbs_dat_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3200__A1 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput419 net419 custom_settings[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3553__I _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3200_ _1649_ _1642_ _1650_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4180_ dffram.data\[46\]\[1\] _2303_ _2305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3131_ _1577_ _1602_ _1604_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3267__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3062_ dffram.data\[43\]\[4\] _1551_ _1552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3964_ dffram.data\[50\]\[0\] _2161_ _2162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ net201 _1103_ _1183_ net135 _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6683_ _0603_ clknet_leaf_74_wb_clk_i dffram.data\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3895_ _1963_ _2117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5634_ _1121_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_147_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__A1 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1066_ _1067_ _0693_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4516_ _2540_ _2541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ dffram.data\[16\]\[5\] dffram.data\[18\]\[5\] dffram.data\[20\]\[5\] dffram.data\[22\]\[5\]
+ _0795_ _0797_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_111_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4447_ net399 _2489_ _2490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input349_I tholin_riscv_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5334__I3 dffram.data\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input251_I sid_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6117_ _0037_ clknet_leaf_17_wb_clk_i dffram.data\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4378_ net445 _2436_ _2439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _1718_ _1734_ _1737_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1435_ _1480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3258__A1 _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_165_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3638__I _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output470_I net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4930__A1 net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4469__I net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4997__A1 _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ dffram.data\[55\]\[2\] _1967_ _1972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5564__I3 dffram.data\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5350_ _0825_ _0858_ net513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_3_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4921__A1 net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3283__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _0772_ _0719_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4301_ dffram.data\[44\]\[4\] _2382_ _2383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ dffram.data\[45\]\[5\] _2335_ _2337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4163_ dffram.data\[15\]\[4\] _2292_ _2293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3114_ _1426_ _1503_ _1592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4094_ dffram.data\[14\]\[4\] _2247_ _2248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3045_ _1501_ _1534_ _1539_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4996_ dffram.data\[40\]\[4\] _2932_ _2933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3412__A1 _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3947_ _2098_ _2146_ _2150_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_82_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input299_I tholin_riscv_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6666_ _0586_ clknet_leaf_67_wb_clk_i dffram.data\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3878_ _2103_ _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5617_ _1117_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_104_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6597_ _0517_ clknet_leaf_119_wb_clk_i net548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5548_ _1042_ _1045_ _1050_ _0719_ _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_42_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input62_I mc14500_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4289__I _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5479_ _0982_ _0983_ _0863_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3651__A1 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5928__B1 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5251__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A1 net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_131_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3890__A1 _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3642__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _2671_ _2826_ _2827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4662__I _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3801_ dffram.data\[13\]\[2\] _2050_ _2053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6520_ _0440_ clknet_leaf_107_wb_clk_i dffram.data\[44\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4781_ wb_counter\[2\] _2770_ _2771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3732_ _1998_ _2006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5147__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _0371_ clknet_leaf_81_wb_clk_i dffram.data\[47\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3663_ _1915_ _1956_ _1959_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5402_ dffram.data\[33\]\[3\] dffram.data\[35\]\[3\] dffram.data\[37\]\[3\] dffram.data\[39\]\[3\]
+ _0799_ _0800_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6382_ _0302_ clknet_leaf_3_wb_clk_i dffram.data\[51\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5333_ _0796_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3594_ _1849_ _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _0773_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_143_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4215_ dffram.data\[1\]\[7\] _2322_ _2326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5195_ _0703_ _0686_ _0704_ _0700_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5870__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4146_ _1724_ _1935_ _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input214_I qcpu_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4077_ _2235_ _2230_ _2236_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ dffram.data\[37\]\[0\] _1529_ _1530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3188__I _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ dffram.data\[41\]\[6\] _2919_ _2922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5481__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5138__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6649_ _0569_ clknet_leaf_110_wb_clk_i dffram.data\[42\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output433_I net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3872__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3624__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__I _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_113_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4000_ _2179_ _2186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3863__A1 dffram.data\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5951_ net16 _1362_ _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ wb_counter\[25\] _2868_ _2869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_38_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5882_ _1274_ _1336_ _1337_ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_118_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _2768_ _2814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_161_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3918__A2 _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ net557 _2739_ _2740_ _2757_ _2758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6503_ _0423_ clknet_leaf_106_wb_clk_i dffram.data\[16\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3715_ _1979_ _1992_ _1995_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6434_ _0354_ clknet_leaf_53_wb_clk_i dffram.data\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4695_ wb_counter\[20\] _2700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3646_ _1919_ _1943_ _1948_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3577_ _1901_ _1903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6365_ _0285_ clknet_leaf_8_wb_clk_i dffram.data\[52\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _0721_ _0815_ _0824_ _0755_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_87_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6296_ _0216_ clknet_leaf_140_wb_clk_i dffram.data\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input164_I qcpu_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput308 tholin_riscv_do[25] net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5247_ _0676_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input331_I tholin_riscv_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput319 tholin_riscv_do[5] net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_110_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3471__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold26 net587 net603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold37 wbs_dat_i[17] net617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold15 _2472_ net592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input25_I ay8913_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ net77 _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold59 _2490_ net636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold48 _2498_ net625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4129_ dffram.data\[20\]\[1\] _2268_ _2270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6020__A2 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4334__A2 net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4477__I _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3381__I _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3845__A1 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_106_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _1492_ _1852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4480_ _0642_ _2505_ _2515_ _2514_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3431_ _1803_ _1805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3362_ _1702_ _1757_ _1759_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ _0070_ clknet_leaf_20_wb_clk_i dffram.data\[62\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6078__A2 _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5101_ design_select\[3\] _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3293_ _1573_ _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6081_ _0001_ clknet_leaf_76_wb_clk_i dffram.data\[36\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4089__A1 _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5825__A2 _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_81_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5032_ _2956_ _2949_ _2957_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ net167 _1365_ _1132_ net303 _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_EDGE_ROW_124_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5865_ net260 _1322_ _1254_ net45 _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4816_ net622 _2800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ _1261_ _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_133_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_79_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input281_I sn76489_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _2742_ _2743_ _2744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4678_ _2670_ _2685_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_112_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3629_ dffram.data\[11\]\[0\] _1938_ _1939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6417_ _0337_ clknet_leaf_28_wb_clk_i dffram.data\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _0268_ clknet_leaf_50_wb_clk_i dffram.data\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput105 pdp11_do[24] net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput127 pdp11_oeb[14] net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput116 pdp11_do[4] net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6279_ _0199_ clknet_leaf_103_wb_clk_i dffram.data\[25\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput138 pdp11_oeb[24] net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput149 pdp11_oeb[4] net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__I _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5427__S1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5752__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3818__A1 dffram.data\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__S0 _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__I _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A1 _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4243__A1 _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3980_ _2108_ _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5766__I _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _1142_ _1143_ net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_116_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _2618_ _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5581_ _0772_ _1074_ _1083_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4532_ _2547_ _2557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4463_ _2499_ net628 _2501_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3414_ _1774_ _1791_ _1794_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6202_ _0122_ clknet_leaf_38_wb_clk_i dffram.data\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4394_ net384 _2444_ _2451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5006__I _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3345_ _1712_ _1742_ _1747_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6133_ _0053_ clknet_leaf_6_wb_clk_i dffram.data\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5354__S0 _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6064_ _1493_ _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3276_ dffram.data\[6\]\[6\] _1697_ _1700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5015_ _2944_ _2939_ _2945_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input127_I pdp11_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4482__A1 _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_132_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5917_ net9 _1362_ _1363_ _1368_ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_152_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5982__A1 net315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5409__S1 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input92_I pdp11_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5848_ net360 _1110_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5779_ _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_141_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_168_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5345__S0 _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output513_I net513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_150_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4473__A1 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_142_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4225__A1 _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_91_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3130_ dffram.data\[8\]\[4\] _1603_ _1604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3061_ _1543_ _1551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4216__A1 _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _2159_ _2161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4767__A2 net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _1177_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6682_ _0602_ clknet_leaf_74_wb_clk_i dffram.data\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3894_ _2115_ _2105_ _2116_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__B2 net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A1 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _1120_ _1130_ net478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5564_ dffram.data\[1\]\[7\] dffram.data\[3\]\[7\] dffram.data\[5\]\[7\] dffram.data\[7\]\[7\]
+ _0696_ _0697_ _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4515_ _2508_ _2503_ _2540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3744__I _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5495_ dffram.data\[24\]\[5\] dffram.data\[26\]\[5\] dffram.data\[28\]\[5\] dffram.data\[30\]\[5\]
+ _0889_ _0890_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5575__S0 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4446_ _2430_ _2489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4377_ _2437_ net607 _2435_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6116_ _0036_ clknet_leaf_43_wb_clk_i dffram.data\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input244_I sid_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3328_ dffram.data\[31\]\[5\] _1735_ _1737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3259_ _1608_ _1640_ _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6047_ _1478_ _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4455__A1 net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_87_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3919__I _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3194__A1 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output463_I net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__S0 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5494__I0 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_138_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_138_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3564__I _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0780_ _0789_ _0708_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4300_ _2374_ _2382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5557__S0 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _2290_ _2334_ _2336_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__S0 _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ _2280_ _2292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3113_ _1590_ _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4437__A1 net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4093_ _2239_ _2247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3044_ dffram.data\[37\]\[7\] _1535_ _1539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5937__A1 _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4995_ _2924_ _2932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3946_ dffram.data\[59\]\[2\] _2147_ _2150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input194_I qcpu_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6665_ _0585_ clknet_leaf_111_wb_clk_i dffram.data\[40\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3877_ _1477_ _2103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _1104_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3176__A1 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6596_ _0516_ clknet_leaf_119_wb_clk_i net547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3474__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ _1047_ _1049_ _0813_ _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input361_I ue1_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5478_ dffram.data\[33\]\[5\] dffram.data\[35\]\[5\] dffram.data\[37\]\[5\] dffram.data\[39\]\[5\]
+ _0804_ _0805_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_148_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input55_I mc14500_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _2475_ net613 _2469_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_126_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4428__A1 net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5928__B2 net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5928__A1 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3649__I _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4943__I _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3800_ _2031_ _2049_ _2052_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4780_ _2549_ _2567_ _2770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3731_ _1998_ _2005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_32_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__A2 _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6450_ _0370_ clknet_leaf_93_wb_clk_i dffram.data\[47\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ dffram.data\[24\]\[5\] _1957_ _1959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ dffram.data\[41\]\[3\] dffram.data\[43\]\[3\] dffram.data\[45\]\[3\] dffram.data\[47\]\[3\]
+ _0859_ _0860_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6381_ _0301_ clknet_leaf_4_wb_clk_i dffram.data\[51\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3593_ _1911_ _1912_ _1914_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _0831_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5263_ _0772_ _0753_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4214_ _2296_ _2321_ _2325_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5194_ net373 _0686_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_167_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4145_ _2088_ _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_3_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__A1 _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ dffram.data\[48\]\[6\] _2231_ _2236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3027_ _1527_ _1529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input207_I qcpu_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _2534_ _2918_ _2921_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3929_ _2132_ _2139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6648_ _0568_ clknet_leaf_110_wb_clk_i dffram.data\[42\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3149__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6579_ _0499_ clknet_leaf_130_wb_clk_i net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4649__A1 net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5846__B1 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3321__A1 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output426_I net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5074__A1 _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5594__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A2 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3560__A1 _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5950_ _1274_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_88_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4901_ _2721_ _2859_ _2868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ net47 _1217_ _1105_ net295 _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4832_ net382 _2804_ _2813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _2755_ _2756_ _2757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4694_ _2618_ _2699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3714_ dffram.data\[12\]\[5\] _1993_ _1995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _0422_ clknet_leaf_106_wb_clk_i dffram.data\[16\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6433_ _0353_ clknet_leaf_52_wb_clk_i dffram.data\[48\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3645_ dffram.data\[11\]\[7\] _1944_ _1948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4879__A1 net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3576_ _1901_ _1902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6364_ _0284_ clknet_leaf_29_wb_clk_i dffram.data\[52\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5315_ _0820_ _0823_ _0749_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_77_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6295_ _0215_ clknet_leaf_140_wb_clk_i dffram.data\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput309 tholin_riscv_do[26] net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5246_ _0709_ _0721_ _0750_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA_input157_I qcpu_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3303__A1 _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold38 net593 net615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold27 _2456_ net604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold16 wbs_dat_i[13] net596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_input324_I tholin_riscv_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold49 wbs_dat_i[2] net629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5177_ net376 _0686_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4128_ _2218_ _2267_ _2269_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I ay8913_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4059_ dffram.data\[48\]\[1\] _2221_ _2224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4803__A1 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4031__A2 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A3 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__A1 _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5770__A2 _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _1803_ _1804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3361_ dffram.data\[2\]\[0\] _1758_ _1759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5100_ net578 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6080_ _0000_ clknet_leaf_74_wb_clk_i dffram.data\[36\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3292_ _1710_ _1705_ _1711_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ dffram.data\[3\]\[7\] _2950_ _2957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__A2 _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ net55 _1315_ _1096_ net101 _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_24_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5864_ _1221_ _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_146_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _2794_ _2798_ _2799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5795_ _1101_ _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5210__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3772__A1 _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4746_ net434 _2688_ _2726_ _2743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ net541 _2676_ _2677_ _2684_ _2685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3628_ _1936_ _1938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6416_ _0336_ clknet_leaf_140_wb_clk_i dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input274_I sn76489_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6347_ _0267_ clknet_leaf_50_wb_clk_i dffram.data\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3482__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3524__A1 dffram.data\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3559_ dffram.data\[10\]\[2\] _1888_ _1891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput106 pdp11_do[25] net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput117 pdp11_do[5] net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6278_ _0198_ clknet_leaf_139_wb_clk_i dffram.data\[25\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput139 pdp11_oeb[25] net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput128 pdp11_oeb[15] net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_157_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5403__S _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5229_ _0738_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_93_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__A1 _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5985__C1 net316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output493_I net493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3763__A1 _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3515__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4488__I _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__S1 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__C1 net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _2546_ _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_96_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5580_ _1042_ _1077_ _1082_ _0753_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _2555_ _2556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4462_ _2468_ _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3413_ dffram.data\[34\]\[1\] _1792_ _1794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6201_ _0121_ clknet_leaf_38_wb_clk_i dffram.data\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4393_ net418 _2447_ _2450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6132_ _0052_ clknet_leaf_35_wb_clk_i dffram.data\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3344_ dffram.data\[30\]\[3\] _1743_ _1747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3275_ _1655_ _1696_ _1699_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6063_ _1492_ _1493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5014_ dffram.data\[3\]\[2\] _2940_ _2945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5354__S1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5916_ _1364_ _1367_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_153_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3993__A1 _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5847_ net187 _1210_ _1097_ net121 _1307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_119_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ _0668_ _0669_ _1168_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA_input85_I mc14500_sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4810__B _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4729_ net550 _2719_ _2720_ _2728_ _2729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4170__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3940__I _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5345__S1 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output506_I net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5958__C1 net307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3736__A1 _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4011__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3060_ _1543_ _1550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _1159_ _0654_ _1181_ net337 _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3962_ _2159_ _2160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6681_ _0601_ clknet_leaf_95_wb_clk_i dffram.data\[38\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3297__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3893_ dffram.data\[21\]\[7\] _2106_ _2116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5632_ net215 _1122_ _1124_ net149 net351 _1127_ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_147_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ dffram.data\[9\]\[7\] dffram.data\[11\]\[7\] dffram.data\[13\]\[7\] dffram.data\[15\]\[7\]
+ _0696_ _0697_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4514_ _2538_ _2531_ _2539_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5494_ _0997_ _0998_ _0765_ _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5575__S1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4445_ net433 _2481_ _2488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ net410 _2432_ _2438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6115_ _0035_ clknet_leaf_44_wb_clk_i dffram.data\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3327_ _1714_ _1734_ _1736_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input237_I sid_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ _1659_ _1683_ _1688_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6046_ _1477_ _1478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3189_ _1641_ _1643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4391__A1 net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__B _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5566__S1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output456_I net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5891__A1 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3670__I _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5946__A2 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold93_I wbs_dat_i[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3957__A1 _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5254__S0 _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3709__A1 _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3185__A2 _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4382__A1 net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5557__S1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__A1 _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ dffram.data\[45\]\[4\] _2335_ _2336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5882__A1 _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _2280_ _2291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5309__S1 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3112_ _1540_ _0791_ _1590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4092_ _2239_ _2246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3043_ _1494_ _1534_ _1538_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__S _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _2924_ _2931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3945_ _2095_ _2146_ _2149_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5493__S0 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6664_ _0584_ clknet_leaf_112_wb_clk_i dffram.data\[40\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _1115_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3876_ _2101_ _2091_ _2102_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6595_ _0515_ clknet_leaf_119_wb_clk_i net546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3755__I _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5546_ _0836_ _1048_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input187_I qcpu_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5477_ dffram.data\[41\]\[5\] dffram.data\[43\]\[5\] dffram.data\[45\]\[5\] dffram.data\[47\]\[5\]
+ _0859_ _0860_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input354_I tholin_riscv_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4428_ net394 _2466_ _2476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5873__B2 net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A1 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input48_I mc14500_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4359_ _2421_ _2423_ _2424_ _2420_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3490__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6029_ _1436_ _1461_ _1462_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3939__A1 _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5484__S0 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4364__A1 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4116__A1 _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__I0 net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _1973_ _1999_ _2004_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _1911_ _1956_ _1958_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_75_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6380_ _0300_ clknet_leaf_26_wb_clk_i dffram.data\[51\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5400_ _0882_ _0907_ net514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3592_ dffram.data\[25\]\[4\] _1913_ _1914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5331_ dffram.data\[24\]\[1\] dffram.data\[26\]\[1\] dffram.data\[28\]\[1\] dffram.data\[30\]\[1\]
+ _0838_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_2_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__A1 net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _0710_ _0714_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_103_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4213_ dffram.data\[1\]\[6\] _2322_ _2325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5193_ net74 _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_143_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4144_ _2237_ _2273_ _2278_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4075_ _2111_ _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_121_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3026_ _1527_ _1528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_84_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input102_I pdp11_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5466__S0 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4977_ dffram.data\[41\]\[5\] _2919_ _2921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3928_ _2101_ _2133_ _2138_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5218__S0 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3859_ _2088_ _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_62_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6647_ _0567_ clknet_leaf_113_wb_clk_i dffram.data\[42\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _0498_ clknet_leaf_130_wb_clk_i net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5529_ _1029_ _1032_ _0814_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5846__A1 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput560 net560 wbs_dat_o[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5846__B2 net323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output419_I net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3085__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_139_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3395__I _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_122_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5880_ net240 _1269_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4900_ _2864_ _2865_ _2867_ _2854_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_38_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _2646_ _2809_ _2812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6014__A1 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5785__I _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4576__A1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ net438 _2629_ _2632_ _2756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4693_ _2625_ _2698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3713_ _1975_ _1992_ _1994_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6501_ _0421_ clknet_leaf_105_wb_clk_i dffram.data\[16\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3644_ _1917_ _1943_ _1947_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6432_ _0352_ clknet_leaf_7_wb_clk_i dffram.data\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _0283_ clknet_leaf_29_wb_clk_i dffram.data\[52\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3575_ _1900_ _1726_ _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_77_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5314_ _0821_ _0822_ _0747_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_77_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6294_ _0214_ clknet_leaf_13_wb_clk_i dffram.data\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_110_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4500__A1 _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold17 net596 net594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold28 wbs_dat_i[26] net608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold39 _2460_ net616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5176_ _0673_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4127_ dffram.data\[20\]\[0\] _2268_ _2269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input317_I tholin_riscv_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4058_ _2094_ _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3067__A1 _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _1508_ _1516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5439__S0 _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__A1 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_156_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4567__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_134_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__I _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5819__B2 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3360_ _1756_ _1758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3291_ dffram.data\[32\]\[2\] _1706_ _1711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _1500_ _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_55_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3049__A1 _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ net248 _1282_ _1260_ net270 net289 _0664_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5863_ net238 _1215_ _1255_ net91 _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5794_ _1259_ _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_1_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4814_ _2796_ _2797_ _2798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_161_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3221__A1 _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5210__A2 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4745_ _2686_ _2741_ _2742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4676_ _2682_ _2683_ _2684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3627_ _1936_ _1937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6415_ _0335_ clknet_leaf_140_wb_clk_i dffram.data\[29\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3558_ _1836_ _1887_ _1890_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6346_ _0266_ clknet_leaf_49_wb_clk_i dffram.data\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input267_I sn76489_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__A1 net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput107 pdp11_do[26] net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput118 pdp11_do[6] net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3489_ _1842_ _1832_ _1843_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6277_ _0197_ clknet_leaf_139_wb_clk_i dffram.data\[25\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput129 pdp11_oeb[16] net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input30_I blinker_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _0722_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5159_ _0666_ _0670_ net522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_99_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5985__B1 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__C2 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3460__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output486_I net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_140_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3673__I _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3279__A1 _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold19_I wbs_dat_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_10_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__I _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4951__A1 _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ net370 _2555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__I _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4461_ net404 _2431_ _2500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3412_ _1769_ _1791_ _1793_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6200_ _0120_ clknet_leaf_100_wb_clk_i dffram.data\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5900__B1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6131_ _0051_ clknet_leaf_37_wb_clk_i dffram.data\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4392_ _2448_ net580 _2446_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3343_ _1710_ _1742_ _1746_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5504__S _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_37_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3274_ dffram.data\[6\]\[5\] _1697_ _1699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6062_ net234 _1473_ _1491_ _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5013_ _1460_ _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_109_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ net163 _1365_ _1366_ net299 _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5846_ net285 _1223_ _1234_ net323 _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_119_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_153_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _0622_ _0656_ _0653_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_17_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4728_ _2725_ _2727_ _2728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3493__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input78_I mc14500_sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4659_ _2418_ _2669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_168_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6329_ _0249_ clknet_leaf_54_wb_clk_i dffram.data\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_129_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5213__I _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__A1 _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3433__A1 _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A1 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_29_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_82_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3961_ _1885_ _2117_ _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3424__A1 _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5700_ _1105_ _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__A4 _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _0600_ clknet_leaf_95_wb_clk_i dffram.data\[38\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3892_ _2114_ _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_2_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5793__I _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1120_ _1129_ net477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_6_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__A1 net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5562_ _0715_ _1051_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_54_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_91_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4513_ dffram.data\[27\]\[7\] _2532_ _2539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5493_ dffram.data\[25\]\[5\] dffram.data\[27\]\[5\] dffram.data\[29\]\[5\] dffram.data\[31\]\[5\]
+ _0838_ _0839_ _0998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4444_ _2486_ _2487_ _2480_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4375_ net444 _2436_ _2437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6114_ _0034_ clknet_leaf_43_wb_clk_i dffram.data\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3326_ dffram.data\[31\]\[4\] _1735_ _1736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5637__C1 net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ net232 _1473_ _1476_ _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA_input132_I pdp11_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3257_ dffram.data\[61\]\[7\] _1684_ _1688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3188_ _1641_ _1642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3663__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_124_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3415__A1 dffram.data\[34\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5917__B _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ net357 _1236_ _1291_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_107_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3951__I _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output449_I net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5628__C1 net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold86_I wbs_dat_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5254__S1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_147_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_147_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4022__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3861__I _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _2103_ _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3111_ _1588_ _1578_ _1589_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4091_ _2227_ _2240_ _2245_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5788__I _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput290 tbb1143_do[4] net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3042_ dffram.data\[37\]\[6\] _1535_ _1538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4692__I _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4993_ _2528_ _2925_ _2930_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3944_ dffram.data\[59\]\[1\] _2147_ _2149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5493__S1 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3875_ dffram.data\[21\]\[3\] _2092_ _2102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_82_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _0583_ clknet_leaf_113_wb_clk_i dffram.data\[40\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5614_ _1094_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6594_ _0514_ clknet_leaf_119_wb_clk_i net545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5545_ dffram.data\[32\]\[7\] dffram.data\[34\]\[7\] dffram.data\[36\]\[7\] dffram.data\[38\]\[7\]
+ _0883_ _0828_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5476_ _0962_ _0981_ net516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_2_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4427_ net428 _2470_ _2475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input347_I tholin_riscv_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4358_ net406 _2406_ _2424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_161_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4289_ _2374_ _2375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3309_ _1722_ _1715_ _1723_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6028_ dffram.data\[36\]\[2\] _1446_ _1462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3636__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6050__A2 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5484__S1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__B _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4777__I _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__I1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3660_ dffram.data\[24\]\[4\] _1957_ _1958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3591_ _1901_ _1913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5330_ _0833_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5261_ _0766_ _0770_ _0708_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5855__A2 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4212_ _2294_ _2321_ _2324_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3591__I _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_44_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5192_ net221 _0701_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_43_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4143_ dffram.data\[20\]\[7\] _2274_ _2278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4074_ _2233_ _2230_ _2234_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _1425_ _1526_ _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3618__A1 _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__S1 _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4976_ _2530_ _2918_ _2920_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3927_ dffram.data\[19\]\[3\] _2134_ _2138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3766__I _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5218__S1 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input297_I tholin_riscv_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3858_ _1443_ _2088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6646_ _0566_ clknet_leaf_113_wb_clk_i dffram.data\[42\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3789_ _2043_ _2038_ _2044_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6577_ _0497_ clknet_leaf_130_wb_clk_i net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _1030_ _1031_ _0802_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I mc14500_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ dffram.data\[25\]\[4\] dffram.data\[27\]\[4\] dffram.data\[29\]\[4\] dffram.data\[31\]\[4\]
+ _0838_ _0839_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_2_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput561 net561 wbs_dat_o[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput550 net550 wbs_dat_o[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3857__A1 _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__B _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5422__S _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_15_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold49_I wbs_dat_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4300__I _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__S0 _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4273__A1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__I _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4830_ _2754_ _2811_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5773__A1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _2548_ wb_counter\[31\] _2755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ _0420_ clknet_leaf_93_wb_clk_i dffram.data\[16\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4692_ _2544_ _2697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3712_ dffram.data\[12\]\[4\] _1993_ _1994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3643_ dffram.data\[11\]\[6\] _1944_ _1947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6431_ _0351_ clknet_leaf_7_wb_clk_i dffram.data\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6362_ _0282_ clknet_leaf_28_wb_clk_i dffram.data\[52\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5313_ dffram.data\[48\]\[1\] dffram.data\[50\]\[1\] dffram.data\[52\]\[1\] dffram.data\[54\]\[1\]
+ _0742_ _0744_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_87_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3574_ _1661_ _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_114_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6293_ _0213_ clknet_leaf_13_wb_clk_i dffram.data\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5384__S0 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5244_ _0715_ _0753_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5175_ dffram.data\[33\]\[0\] dffram.data\[35\]\[0\] dffram.data\[37\]\[0\] dffram.data\[39\]\[0\]
+ _0678_ _0683_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xhold18 _2451_ net595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold29 net669 net606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4126_ _2266_ _2268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5300__I1 dffram.data\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ _2218_ _2220_ _2222_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input212_I qcpu_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3008_ _1508_ _1515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__S1 _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4016__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_130_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4959_ _2536_ _2905_ _2909_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3496__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6629_ _0549_ clknet_leaf_126_wb_clk_i wb_counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5216__I _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output529_I net529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output431_I net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__A1 _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_59_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3290_ _1570_ _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5366__S0 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__A1 _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4246__A1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5931_ _1376_ _1380_ net493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5796__I _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ net362 _1098_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _1221_ _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4813_ _2793_ _2628_ _2790_ _2797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4744_ wb_counter\[28\] _2741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4675_ net422 _2655_ _2660_ _2683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3626_ _1507_ _1935_ _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6414_ _0334_ clknet_leaf_139_wb_clk_i dffram.data\[29\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3557_ dffram.data\[10\]\[1\] _1888_ _1890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6345_ _0265_ clknet_leaf_49_wb_clk_i dffram.data\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6276_ _0196_ clknet_leaf_64_wb_clk_i dffram.data\[25\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input162_I qcpu_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput108 pdp11_do[27] net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3488_ dffram.data\[58\]\[3\] _1833_ _1843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5227_ _0728_ _0732_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput119 pdp11_do[7] net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_102_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input23_I ay8913_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5158_ _0656_ _0667_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4109_ dffram.data\[47\]\[2\] _2254_ _2257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5089_ _2948_ _2991_ _2993_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4237__A1 _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__B2 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5985__A1 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__A1 net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output479_I net479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_120_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4476__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5976__A1 net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A1 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__B2 net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4460_ net438 _2492_ _2499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5900__A1 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3411_ dffram.data\[34\]\[0\] _1792_ _1793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ net383 _2444_ _2449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5900__B2 net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3342_ dffram.data\[30\]\[2\] _1743_ _1746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6130_ _0050_ clknet_leaf_36_wb_clk_i dffram.data\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3273_ _1651_ _1696_ _1698_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6061_ _1489_ _1464_ _1490_ _1437_ _1491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5012_ _2942_ _2939_ _2943_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_109_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__S _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__I _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5511__S0 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5914_ _1125_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5845_ _1285_ _1300_ _1301_ _1305_ net482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _1231_ _1235_ _1243_ net508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_134_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ net431 _2688_ _2726_ _2727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input377_I wbs_adr_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _2645_ _2668_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput90 pdp11_do[10] net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3609_ dffram.data\[56\]\[1\] _1924_ _1926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _2546_ _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_168_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6328_ _0248_ clknet_leaf_0_wb_clk_i dffram.data\[54\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6259_ _0179_ clknet_leaf_29_wb_clk_i dffram.data\[57\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4458__A1 net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5958__B2 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5958__A1 net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__S0 _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4630__A1 _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3197__A1 _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold31_I wbs_dat_i[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3121__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__A1 _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ _2088_ _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_69_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3891_ _1499_ _2114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5630_ net214 _1122_ _1124_ net148 net350 _1127_ _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_5_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ _1042_ _1054_ _1063_ _0753_ _1064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_81_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4512_ _1500_ _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5492_ dffram.data\[17\]\[5\] dffram.data\[19\]\[5\] dffram.data\[21\]\[5\] dffram.data\[23\]\[5\]
+ _0884_ _0885_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__A1 net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4443_ net398 _2478_ _2487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ _2422_ _2436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6113_ _0033_ clknet_leaf_43_wb_clk_i dffram.data\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3325_ _1727_ _1735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_146_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3256_ _1657_ _1683_ _1687_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6044_ _1474_ _1464_ _1475_ _1457_ _1476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_42_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_163_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3187_ _1638_ _1640_ _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input125_I pdp11_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input90_I pdp11_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ _1214_ _1289_ _1290_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_107_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5759_ net258 _1223_ _1103_ net155 _1227_ _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__S _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3009__I _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3351__A1 _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold1_I wbs_dat_i[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output511_I net511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3103__A1 _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__A1 net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6055__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__A2 _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5134__I _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ dffram.data\[7\]\[7\] _1579_ _1589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4090_ dffram.data\[14\]\[3\] _2241_ _2245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5095__A1 _2956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3041_ _1487_ _1534_ _1537_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4973__I _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput280 sn76489_do[4] net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput291 tholin_riscv_do[0] net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4992_ dffram.data\[40\]\[3\] _2926_ _2930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3943_ _2089_ _2146_ _2148_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3874_ _2100_ _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_82_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _0582_ clknet_leaf_113_wb_clk_i dffram.data\[40\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5613_ _1113_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _0513_ clknet_leaf_118_wb_clk_i net543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ _0802_ _1046_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5475_ _0963_ _0970_ _0979_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_148_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4426_ _2473_ net598 _2469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_165_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3333__A1 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input242_I sid_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5044__I _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4357_ _2422_ _2423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_126_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4288_ _2074_ _1542_ _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3308_ dffram.data\[32\]\[7\] _1716_ _1723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3239_ _1676_ _1677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6027_ _1460_ _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5561__A2 _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3962__I _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3572__A1 _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output559_I net559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output461_I net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__I _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3202__I _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4033__I _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5001__A1 _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3590_ _1901_ _1912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5260_ _0767_ _0768_ _0769_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4211_ dffram.data\[1\]\[5\] _2322_ _2324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_143_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5068__A1 _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _2235_ _2273_ _2277_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073_ dffram.data\[48\]\[5\] _2231_ _2234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3024_ _1525_ _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_121_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4208__I _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4975_ dffram.data\[41\]\[4\] _2919_ _2920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3926_ _2098_ _2133_ _2137_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input192_I qcpu_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6645_ _0565_ clknet_leaf_84_wb_clk_i dffram.data\[42\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _2045_ _2082_ _2087_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_119_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ dffram.data\[53\]\[6\] _2039_ _2044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6576_ _0496_ clknet_leaf_130_wb_clk_i net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5527_ dffram.data\[16\]\[6\] dffram.data\[18\]\[6\] dffram.data\[20\]\[6\] dffram.data\[22\]\[6\]
+ _0795_ _0797_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4878__I _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input53_I mc14500_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3306__A1 _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput562 net562 wbs_dat_o[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput540 net540 wbs_dat_o[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput551 net551 wbs_dat_o[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5458_ dffram.data\[17\]\[4\] dffram.data\[19\]\[4\] dffram.data\[21\]\[4\] dffram.data\[23\]\[4\]
+ _0884_ _0885_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_121_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ _0781_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4409_ net388 _2455_ _2462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_139_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__S1 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5412__I _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4760_ _2434_ _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4691_ _2692_ _2696_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3711_ _1985_ _1993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3642_ _1915_ _1943_ _1946_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6430_ _0350_ clknet_leaf_5_wb_clk_i dffram.data\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_131_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_131_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_157_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3536__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6361_ _0281_ clknet_leaf_29_wb_clk_i dffram.data\[52\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ dffram.data\[56\]\[1\] dffram.data\[58\]\[1\] dffram.data\[60\]\[1\] dffram.data\[62\]\[1\]
+ _0739_ _0740_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3573_ _1829_ _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_114_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6292_ _0212_ clknet_leaf_48_wb_clk_i dffram.data\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5243_ _0751_ _0716_ _0717_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_41_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ dffram.data\[41\]\[0\] dffram.data\[43\]\[0\] dffram.data\[45\]\[0\] dffram.data\[47\]\[0\]
+ _0678_ _0683_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xhold19 wbs_dat_i[20] net599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4125_ _2266_ _2267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_166_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5322__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4056_ dffram.data\[48\]\[0\] _2221_ _2222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3007_ _1470_ _1509_ _1514_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input205_I qcpu_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ dffram.data\[42\]\[6\] _2906_ _2909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3775__A1 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3909_ dffram.data\[51\]\[4\] _2126_ _2127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5992__I net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _2704_ _2709_ _2715_ _2847_ _2858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_117_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6628_ _0548_ clknet_leaf_127_wb_clk_i wb_counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3527__A1 _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6559_ _0479_ clknet_leaf_106_wb_clk_i net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_7_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output424_I net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5232__I _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6063__I _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3687__I _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4311__I _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5407__I _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_94_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4191__A1 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__S1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5930_ net11 _1362_ _1363_ _1379_ _1380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5294__I1 _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5994__A2 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5861_ net157 _1154_ _1312_ net3 net293 _1181_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_5_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5792_ _1246_ _1248_ _1251_ _1258_ net509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_111_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ net622 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4743_ _2624_ _2740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3757__A1 _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6413_ _0333_ clknet_leaf_139_wb_clk_i dffram.data\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4674_ _2653_ wb_counter\[17\] _2682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3625_ _1590_ _1935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5317__I _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3556_ _1830_ _1887_ _1889_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6344_ _0264_ clknet_leaf_3_wb_clk_i dffram.data\[53\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _0195_ clknet_leaf_65_wb_clk_i dffram.data\[25\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput109 pdp11_do[28] net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3487_ _1841_ _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5226_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_input155_I qcpu_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4377__B _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input322_I tholin_riscv_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0666_ _0669_ net530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4108_ _2223_ _2253_ _2256_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5088_ dffram.data\[9\]\[4\] _2992_ _2993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input16_I ay8913_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4039_ _2165_ _2206_ _2210_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5985__A2 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5936__B _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4173__A1 _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5338__S _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5137__I _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3410_ _1790_ _1792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4164__A1 _2290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ net417 _2447_ _2448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3341_ _1708_ _1742_ _1745_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3880__I _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I ay8913_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3272_ dffram.data\[6\]\[4\] _1697_ _1698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6060_ net408 _1465_ _1490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5011_ dffram.data\[3\]\[1\] _2940_ _2943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5600__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5511__S1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _1113_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5844_ net359 _1236_ _1304_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_17_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5775_ net357 _1236_ _1239_ _1242_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_146_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4726_ _2631_ _2726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ net538 _2651_ _2652_ _2667_ _2668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput91 pdp11_do[11] net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3608_ _1899_ _1923_ _1925_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input272_I sn76489_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput80 mc14500_sram_gwe net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3902__A1 _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4588_ _1026_ _1041_ _2552_ _2607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6327_ _0247_ clknet_leaf_9_wb_clk_i dffram.data\[54\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3539_ dffram.data\[57\]\[3\] _1874_ _1878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6258_ _0178_ clknet_leaf_30_wb_clk_i dffram.data\[57\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6189_ _0109_ clknet_leaf_102_wb_clk_i dffram.data\[31\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5209_ net225 _0647_ _0718_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_93_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A2 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5502__S1 _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4126__I _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output491_I net491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4394__A1 net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4146__A1 _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5497__I1 _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5257__S0 _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3890_ _2112_ _2105_ _2113_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5421__I1 dffram.data\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5560_ _1056_ _1061_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_38_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5491_ _0944_ _0988_ _0995_ _0961_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_4511_ _2536_ _2531_ _2537_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4442_ net432 _2481_ _2486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5885__A1 net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4373_ _2429_ _2433_ _2435_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _0032_ clknet_leaf_112_wb_clk_i dffram.data\[43\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3324_ _1727_ _1734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5637__A1 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5637__B2 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3255_ dffram.data\[61\]\[6\] _1684_ _1687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6043_ net406 _1465_ _1475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_163_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3186_ _1639_ _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_124_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input118_I pdp11_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__S0 _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ net184 _1261_ _1232_ net70 _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5758_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A1 net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input83_I mc14500_sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ _2699_ _2709_ _2711_ _2712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5689_ _1172_ _1173_ net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4128__A1 _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__S0 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5628__B2 net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A1 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__S _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output504_I net504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A1 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6071__I _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__A1 net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4119__A1 dffram.data\[47\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5316__B1 _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3040_ dffram.data\[37\]\[5\] _1535_ _1537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput281 sn76489_do[5] net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput270 sn76489_do[20] net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput292 tholin_riscv_do[10] net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_69_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6044__A1 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4991_ _2526_ _2925_ _2929_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3942_ dffram.data\[59\]\[0\] _2147_ _2148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3873_ _1468_ _2100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6661_ _0581_ clknet_leaf_85_wb_clk_i dffram.data\[40\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5612_ _1100_ _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6592_ _0512_ clknet_leaf_119_wb_clk_i net542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4358__A1 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ dffram.data\[40\]\[7\] dffram.data\[42\]\[7\] dffram.data\[44\]\[7\] dffram.data\[46\]\[7\]
+ _0883_ _0828_ _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _0791_ _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5402__S0 _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ net393 _2466_ _2474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4356_ _2405_ _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3307_ _1587_ _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_126_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5261__S _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4287_ _2359_ _2368_ _2373_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input235_I qcpu_sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _1459_ _1460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3238_ _1526_ _1623_ _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3169_ dffram.data\[63\]\[2\] _1626_ _1629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4404__I _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__B2 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__A1 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output454_I net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold91_I wbs_dat_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__B1 _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4210_ _2290_ _2321_ _2323_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4984__I _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _0643_ _0645_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_43_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_143_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ dffram.data\[20\]\[6\] _2274_ _2277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ _2108_ _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ _1427_ _1505_ _1525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _2911_ _2919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4579__A1 net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3925_ dffram.data\[19\]\[2\] _2134_ _2137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_158_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6644_ _0564_ clknet_leaf_83_wb_clk_i dffram.data\[42\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ dffram.data\[52\]\[7\] _2083_ _2087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3003__A1 _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__S _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3787_ _1852_ _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6575_ _0495_ clknet_leaf_130_wb_clk_i net544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5526_ dffram.data\[24\]\[6\] dffram.data\[26\]\[6\] dffram.data\[28\]\[6\] dffram.data\[30\]\[6\]
+ _0841_ _0842_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input185_I qcpu_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4751__A1 net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _0773_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input352_I tholin_riscv_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput530 net530 rst_tholin_riscv vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5055__I _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4408_ net422 _2458_ _2461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput563 net563 wbs_dat_o[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput541 net541 wbs_dat_o[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput552 net552 wbs_dat_o[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input46_I mc14500_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5388_ dffram.data\[9\]\[2\] dffram.data\[11\]\[2\] dffram.data\[13\]\[2\] dffram.data\[15\]\[2\]
+ _0848_ _0849_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4339_ _2408_ _2409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6009_ _1444_ _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5767__B1 _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3242__A1 _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_42_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3481__A1 _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3233__A1 _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3710_ _1985_ _1992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ net543 _2676_ _2677_ _2695_ _2696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3641_ dffram.data\[11\]\[5\] _1944_ _1946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3883__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3572_ _1856_ _1893_ _1898_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6360_ _0280_ clknet_leaf_142_wb_clk_i dffram.data\[22\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _0818_ _0819_ _0736_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_114_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6291_ _0211_ clknet_leaf_48_wb_clk_i dffram.data\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_100_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5242_ net225 _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4928__B _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5173_ _0682_ _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4124_ _2074_ _2265_ _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput1 ay8913_do[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4219__I _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4055_ _2219_ _2221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3006_ dffram.data\[35\]\[3\] _1510_ _1514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input100_I pdp11_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4957_ _2534_ _2905_ _2908_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4972__A1 _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3908_ _2118_ _2126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4888_ _2841_ _2856_ _2857_ _2854_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_35_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3839_ _2075_ _2077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6627_ _0547_ clknet_leaf_127_wb_clk_i wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6558_ _0478_ clknet_leaf_115_wb_clk_i net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_15_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6489_ _0409_ clknet_leaf_81_wb_clk_i dffram.data\[45\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5509_ dffram.data\[33\]\[6\] dffram.data\[35\]\[6\] dffram.data\[37\]\[6\] dffram.data\[39\]\[6\]
+ _0804_ _0805_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_125_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output417_I net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__B _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__I _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3454__A1 _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5860_ _1313_ _1318_ net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4811_ _2502_ _2618_ _2508_ _2403_ _2795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_158_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _1253_ _1256_ _1257_ _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_115_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4742_ _2544_ _2739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4673_ _2670_ _2681_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_151_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6412_ _0332_ clknet_leaf_63_wb_clk_i dffram.data\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3509__A2 _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3624_ _1919_ _1929_ _1934_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4502__I _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5903__B1 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3118__I _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3555_ dffram.data\[10\]\[0\] _1888_ _1889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6343_ _0263_ clknet_leaf_3_wb_clk_i dffram.data\[53\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _0194_ clknet_leaf_65_wb_clk_i dffram.data\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3486_ _1468_ _1841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input148_I pdp11_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__A2 _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__I _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _0651_ _0667_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4107_ dffram.data\[47\]\[1\] _2254_ _2256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5087_ _2984_ _2992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input315_I tholin_riscv_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4038_ dffram.data\[4\]\[2\] _2207_ _2210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3445__A1 _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5989_ _1424_ _1425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_23_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4945__A1 _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_25_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_160_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__S _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__C1 net325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_54_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3684__A1 _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3340_ dffram.data\[30\]\[1\] _1743_ _1745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_111_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__C1 net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5010_ _1452_ _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3271_ _1689_ _1697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3675__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__A3 _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ net51 _1315_ _1267_ net97 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _1257_ _1302_ _1303_ _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__S _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5774_ _1240_ _1241_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4725_ _2686_ wb_counter\[25\] _2725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _2627_ _2664_ _2666_ _2667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3607_ dffram.data\[56\]\[0\] _1924_ _1925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput70 mc14500_do[6] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput81 mc14500_sram_in[0] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4587_ net561 _2583_ _2606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput92 pdp11_do[12] net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3538_ _1839_ _1873_ _1877_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input265_I sn76489_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6326_ _0246_ clknet_leaf_0_wb_clk_i dffram.data\[54\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _0177_ clknet_leaf_39_wb_clk_i dffram.data\[57\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3469_ dffram.data\[5\]\[7\] _1824_ _1828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_129_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6188_ _0108_ clknet_leaf_72_wb_clk_i dffram.data\[31\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5208_ _0716_ _0717_ _0647_ _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5139_ _0639_ _0654_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3418__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4091__A1 _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output484_I net484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_42_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3657__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__S1 _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_51_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4909__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5490_ _0991_ _0994_ _0924_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4510_ dffram.data\[27\]\[6\] _2532_ _2537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3891__I _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _2484_ _2485_ _2480_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3896__A1 _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _0031_ clknet_leaf_87_wb_clk_i dffram.data\[43\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_60_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4372_ _2434_ _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3323_ _1712_ _1728_ _1733_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3254_ _1655_ _1683_ _1686_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6042_ net85 _1474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_163_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3185_ _1560_ _1432_ _1639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5496__S1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3820__A1 dffram.data\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5826_ net118 _1155_ _1126_ net320 _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5757_ net1 _1225_ _1096_ net89 _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ net428 _2705_ _2710_ _2711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5688_ net196 _1163_ _1166_ net130 net332 _1164_ _1173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input76_I mc14500_sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4639_ _2625_ _2652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__S1 _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6309_ _0229_ clknet_leaf_1_wb_clk_i dffram.data\[55\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5628__A2 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__S1 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3976__I _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__S _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__S0 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput260 sn76489_do[11] net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput271 sn76489_do[21] net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput293 tholin_riscv_do[11] net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_106_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput282 sn76489_do[6] net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_125_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ dffram.data\[40\]\[2\] _2926_ _2929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3802__A1 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3941_ _2145_ _2147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ _2098_ _2091_ _2099_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6660_ _0580_ clknet_leaf_85_wb_clk_i dffram.data\[40\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_82_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5611_ net367 _1111_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6591_ _0511_ clknet_leaf_119_wb_clk_i net541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5542_ _1043_ _1044_ _0747_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5473_ _0973_ _0978_ _0905_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_148_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5402__S1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ net427 _2470_ _2473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4355_ net440 _2421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5542__S _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3306_ _1720_ _1715_ _1721_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4286_ dffram.data\[18\]\[7\] _2369_ _2373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input130_I pdp11_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3237_ _1659_ _1670_ _1675_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5491__B1 _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ net230 _1438_ _1458_ _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_20_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3168_ _1568_ _1625_ _1628_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input228_I qcpu_sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3099_ _1577_ _1578_ _1580_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3796__I _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _1237_ _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5546__A1 _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__I _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output447_I net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3036__I _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4285__A1 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4037__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__C _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold84_I wbs_dat_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4330__I net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5362__S _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4140_ _2233_ _2273_ _2276_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_143_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5161__I _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _2229_ _2230_ _2232_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_160_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3022_ _1523_ net656 _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_121_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4028__A1 _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _2911_ _2918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3924_ _2095_ _2133_ _2136_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5379__I1 dffram.data\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _0563_ clknet_leaf_86_wb_clk_i dffram.data\[42\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_93_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3855_ _2043_ _2082_ _2086_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4200__A1 _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3786_ _2041_ _2038_ _2042_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _0494_ clknet_leaf_134_wb_clk_i net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5525_ _1027_ _1028_ _0765_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput520 net520 rst_ay8913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__4240__I _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5456_ _0944_ _0951_ _0960_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_48_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input178_I qcpu_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput531 net531 rst_ue1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4407_ _2459_ net616 _2457_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput542 net542 wbs_dat_o[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput553 net553 wbs_dat_o[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input345_I tholin_riscv_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5387_ _0888_ _0894_ _0846_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput564 net564 wbs_dat_o[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4338_ _2405_ _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input39_I diceroll_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4269_ _2361_ _2363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5303__I1 _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4267__A1 _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6008_ _1443_ _1444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5767__B2 net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5767__A1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4415__I _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__S0 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__S0 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__A1 net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3640_ _1911_ _1943_ _1945_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5930__A1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3571_ dffram.data\[10\]\[7\] _1894_ _1898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6290_ _0210_ clknet_leaf_49_wb_clk_i dffram.data\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5310_ dffram.data\[57\]\[1\] dffram.data\[59\]\[1\] dffram.data\[61\]\[1\] dffram.data\[63\]\[1\]
+ _0729_ _0731_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_84_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__S0 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4995__I _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__A1 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ _0701_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5172_ _0681_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4123_ _2011_ _2265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_140_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput2 ay8913_do[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4054_ _2219_ _2220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3005_ _1461_ _1509_ _1513_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5541__S0 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__C _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ dffram.data\[42\]\[5\] _2906_ _2908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4421__A1 net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3907_ _2118_ _2125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4887_ net394 _2844_ _2857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input295_I tholin_riscv_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3838_ _2075_ _2076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6626_ _0546_ clknet_leaf_126_wb_clk_i wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5921__A1 net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6557_ _0477_ clknet_leaf_106_wb_clk_i net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_162_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3769_ _2026_ _2028_ _2030_ _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_89_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5066__I _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5508_ dffram.data\[41\]\[6\] dffram.data\[43\]\[6\] dffram.data\[45\]\[6\] dffram.data\[47\]\[6\]
+ _0799_ _0800_ _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6488_ _0408_ clknet_leaf_56_wb_clk_i dffram.data\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ dffram.data\[41\]\[4\] dffram.data\[43\]\[4\] dffram.data\[45\]\[4\] dffram.data\[47\]\[4\]
+ _0859_ _0860_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3314__I _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__A1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_70_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3215__A2 _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5460__I0 _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4412__A1 net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5912__A1 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__B2 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5979__A1 net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__S0 _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4055__I _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4810_ _2793_ _2790_ _2628_ _2794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5790_ net31 _0627_ _1213_ _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_118_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _2734_ _2738_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4672_ net540 _2676_ _2677_ _2680_ _2681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5903__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_116_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6411_ _0331_ clknet_leaf_63_wb_clk_i dffram.data\[29\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3623_ dffram.data\[56\]\[7\] _1930_ _1934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3554_ _1886_ _1888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6342_ _0262_ clknet_leaf_3_wb_clk_i dffram.data\[53\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5614__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3390__A1 _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3485_ _1839_ _1832_ _1840_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6273_ _0193_ clknet_leaf_62_wb_clk_i dffram.data\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5667__B1 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5224_ _0700_ _0687_ _0689_ _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_110_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5155_ _0666_ _0668_ net525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5419__B1 _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4106_ _2218_ _2253_ _2255_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5086_ _2984_ _2991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4037_ _2163_ _2206_ _2209_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input308_I tholin_riscv_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input210_I qcpu_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5988_ _1423_ _0944_ _1424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4939_ net532 _2846_ _2895_ _2896_ _2897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_133_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _0529_ clknet_leaf_132_wb_clk_i wb_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5122__A2 _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3133__A1 _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output527_I net527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5460__S _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4633__A1 _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4603__I _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__B1 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3219__I _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3372__A1 _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3270_ _1689_ _1696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4872__A1 net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5967__A4 _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5911_ _1213_ _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_88_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5842_ net186 _1261_ _1139_ net27 _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5773_ net12 _1225_ _1096_ net100 _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_115_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__I _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4724_ _2714_ _2724_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3129__I _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4655_ net419 _2665_ _2632_ _2666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 mc14500_do[25] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3606_ _1922_ _1924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput71 mc14500_do[7] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput82 mc14500_sram_in[1] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _2599_ _2604_ _2605_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput93 pdp11_do[13] net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3537_ dffram.data\[57\]\[2\] _1874_ _1877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6325_ _0245_ clknet_leaf_0_wb_clk_i dffram.data\[54\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input160_I qcpu_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input258_I sn76489_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3468_ _1786_ _1823_ _1827_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6256_ _0176_ clknet_leaf_13_wb_clk_i dffram.data\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_129_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6187_ _0107_ clknet_leaf_72_wb_clk_i dffram.data\[31\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5280__S _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3399_ _1581_ _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5207_ net78 _0650_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input21_I ay8913_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _0637_ _0619_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_99_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5258__I3 dffram.data\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ dffram.data\[39\]\[5\] _2979_ _2981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output477_I net477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__B1 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5894__A3 _1342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3354__A1 dffram.data\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__A1 _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3593__A1 _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4440_ net397 _2478_ _2485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3345__A1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ _0030_ clknet_leaf_87_wb_clk_i dffram.data\[43\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _2418_ _2434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3322_ dffram.data\[31\]\[3\] _1729_ _1733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3253_ dffram.data\[61\]\[5\] _1684_ _1686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6041_ _1437_ _1473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_0_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3184_ _1622_ _1638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_163_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5825_ net282 _1287_ _1250_ net25 _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_146_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__I _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5756_ _1224_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5687_ _0626_ _1171_ _1110_ _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_60_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _2630_ _2710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input375_I wbs_adr_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _2582_ _2651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input69_I mc14500_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5730__C1 net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4569_ _2584_ _2590_ _2574_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6308_ _0228_ clknet_leaf_25_wb_clk_i dffram.data\[55\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5089__A1 _2948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6239_ _0159_ clknet_leaf_18_wb_clk_i dffram.data\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4836__A1 wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3575__A1 _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5316__A2 _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3327__A1 _1714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__S1 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput250 sid_do[3] net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput261 sn76489_do[12] net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput272 sn76489_do[22] net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput294 tholin_riscv_do[12] net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_106_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput283 sn76489_do[7] net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_19_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3940_ _2145_ _2146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ dffram.data\[21\]\[2\] _2092_ _2099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5610_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6590_ _0510_ clknet_leaf_120_wb_clk_i net540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5541_ dffram.data\[33\]\[7\] dffram.data\[35\]\[7\] dffram.data\[37\]\[7\] dffram.data\[39\]\[7\]
+ _0724_ _0727_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3566__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _0974_ _0977_ _0903_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4423_ _2471_ net592 _2469_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_165_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4354_ _2416_ _2407_ _2417_ _2420_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3305_ dffram.data\[32\]\[6\] _1716_ _1721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4285_ _2357_ _2368_ _2372_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6024_ _1455_ _1216_ _1456_ _1457_ _1458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3236_ dffram.data\[33\]\[7\] _1671_ _1675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3167_ dffram.data\[63\]\[1\] _1626_ _1628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input123_I pdp11_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ dffram.data\[7\]\[4\] _1579_ _1580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ net280 _1223_ _1210_ net182 _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5739_ _1185_ _1207_ _1208_ _1209_ net472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_31_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3309__A1 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4148__I _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_109_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3548__A1 _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold77_I wbs_adr_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3720__A1 _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_118_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_160_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4070_ dffram.data\[48\]\[4\] _2231_ _2232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_160_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3021_ net412 net379 _1524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3897__I _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4972_ _2528_ _2912_ _2917_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3923_ dffram.data\[19\]\[1\] _2134_ _2136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_158_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_127_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6642_ _0562_ clknet_leaf_84_wb_clk_i dffram.data\[42\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3854_ dffram.data\[52\]\[6\] _2083_ _2086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6573_ _0493_ clknet_leaf_108_wb_clk_i dffram.data\[27\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3785_ dffram.data\[53\]\[5\] _2039_ _2042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4521__I net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5524_ dffram.data\[25\]\[6\] dffram.data\[27\]\[6\] dffram.data\[29\]\[6\] dffram.data\[31\]\[6\]
+ _0838_ _0839_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput510 net510 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5455_ _0754_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_70_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput521 net521 rst_blinker vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ net387 _2455_ _2460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput543 net543 wbs_dat_o[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput554 net554 wbs_dat_o[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput532 net532 wbs_ack_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5386_ _0891_ _0892_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input240_I sid_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__I _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4337_ _2406_ _2407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input338_I tholin_riscv_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4268_ _2361_ _2362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3219_ _1663_ _1665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6007_ net228 _1438_ _1442_ _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4199_ dffram.data\[1\]\[0\] _2316_ _2317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3778__A1 _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4431__I _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5378__S1 _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__S _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5550__S1 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__A1 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3510__I _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4606__I _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3769__A1 _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3570_ _1853_ _1893_ _1897_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4341__I _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5369__S1 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5373__S _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _0737_ _0748_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5171_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _2237_ _2259_ _2264_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_85_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4053_ _1921_ _2117_ _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xinput3 ay8913_do[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3004_ dffram.data\[35\]\[2\] _1510_ _1513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5997__A2 _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__S1 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_135_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3420__I _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _2530_ _2905_ _2907_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3906_ _2101_ _2119_ _2124_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4886_ _2709_ _2855_ _2856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ _2074_ _1964_ _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_7_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _0545_ clknet_leaf_126_wb_clk_i wb_counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input288_I tbb1143_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5921__A2 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input190_I qcpu_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3768_ dffram.data\[53\]\[0\] _2029_ _2030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4185__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6556_ _0476_ clknet_leaf_115_wb_clk_i net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _0996_ _1011_ net517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3932__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_144_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6487_ _0407_ clknet_leaf_56_wb_clk_i dffram.data\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3699_ _1434_ _1935_ _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input51_I mc14500_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ _0720_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_7_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5369_ dffram.data\[56\]\[2\] dffram.data\[58\]\[2\] dffram.data\[60\]\[2\] dffram.data\[62\]\[2\]
+ _0739_ _0740_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_153_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3999__A1 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4161__I _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_162_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5912__A2 _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__I1 _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5523__S1 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3240__I _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4740_ net552 _2719_ _2720_ _2737_ _2738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5167__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4671_ _2678_ _2679_ _2680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _0330_ clknet_leaf_64_wb_clk_i dffram.data\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4167__A1 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3622_ _1917_ _1929_ _1933_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5903__A2 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3914__A1 _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _0261_ clknet_leaf_3_wb_clk_i dffram.data\[53\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3553_ _1886_ _1887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3484_ dffram.data\[58\]\[2\] _1833_ _1840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _0192_ clknet_leaf_10_wb_clk_i dffram.data\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5667__A1 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5667__B2 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ net224 _0700_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5154_ _0620_ _0622_ _0667_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_138_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4105_ dffram.data\[47\]\[0\] _2254_ _2255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5085_ _2946_ _2985_ _2990_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4036_ dffram.data\[4\]\[1\] _2207_ _2209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3150__I _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input203_I qcpu_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _1057_ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4938_ _2508_ net660 _2553_ _2896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input99_I pdp11_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5077__I _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4869_ wb_counter\[18\] _2834_ _2842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _0528_ clknet_leaf_131_wb_clk_i wb_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _0459_ clknet_leaf_123_wb_clk_i net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_140_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5658__B2 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5658__A1 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3325__I _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output422_I net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3060__I _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__S0 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4397__A1 net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__B2 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5649__A1 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5649__B2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_119_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5113__A3 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5450__I _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5910_ _1266_ _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_152_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5841_ net284 _1259_ _1126_ net322 _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5772_ net269 _1222_ _1170_ net32 _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ net549 _2719_ _2720_ _2723_ _2724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5432__S0 _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _2614_ _2665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5625__I _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput61 mc14500_do[26] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput50 mc14500_do[16] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3605_ _1922_ _1923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput72 mc14500_do[8] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4585_ _2419_ _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput94 pdp11_do[14] net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3536_ _1836_ _1873_ _1876_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6324_ _0244_ clknet_leaf_19_wb_clk_i dffram.data\[54\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput83 mc14500_sram_in[2] net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_168_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _0175_ clknet_leaf_14_wb_clk_i dffram.data\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input153_I pdp11_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3467_ dffram.data\[5\]\[6\] _1824_ _1827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3115__A2 _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ net377 _0712_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_129_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6186_ _0106_ clknet_leaf_62_wb_clk_i dffram.data\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3398_ _1780_ _1781_ _1783_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5137_ _0649_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_165_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input320_I tholin_riscv_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _2948_ _2978_ _2980_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5499__S0 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input14_I ay8913_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A1 _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ dffram.data\[49\]\[3\] _2194_ _2198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A1 net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5879__A1 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5423__S0 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput410 net606 net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4854__A2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_4_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5406__I1 _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4614__I _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5414__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4370_ net409 _2432_ _2433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3321_ _1710_ _1728_ _1732_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6040_ _1435_ _1472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3252_ _1651_ _1683_ _1685_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input6_I ay8913_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _1556_ _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_163_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_87_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_141_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_16_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _1259_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_119_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5755_ _1138_ _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3033__A1 _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5686_ _1170_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ wb_counter\[22\] _2709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_45_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5405__S0 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__I _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4637_ _2645_ _2650_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input368_I wb_rst_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input270_I sn76489_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4568_ _2545_ _2588_ _2589_ _2590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_25_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3519_ _1842_ _1860_ _1865_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4499_ dffram.data\[27\]\[3\] _2522_ _2529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6307_ _0227_ clknet_leaf_25_wb_clk_i dffram.data\[55\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _0158_ clknet_leaf_17_wb_clk_i dffram.data\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6169_ _0089_ clknet_leaf_34_wb_clk_i dffram.data\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold22_I wbs_dat_i[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput240 sid_do[13] net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput251 sid_do[4] net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput262 sn76489_do[13] net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput295 tholin_riscv_do[13] net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_106_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput284 sn76489_do[8] net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput273 sn76489_do[23] net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_19_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_86_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3263__A1 _1637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4344__I net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3870_ _2097_ _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_85_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3015__A1 _1494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ dffram.data\[41\]\[7\] dffram.data\[43\]\[7\] dffram.data\[45\]\[7\] dffram.data\[47\]\[7\]
+ _0724_ _0727_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ dffram.data\[0\]\[4\] dffram.data\[2\]\[4\] dffram.data\[4\]\[4\] dffram.data\[6\]\[4\]
+ _0975_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_48_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_134_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4422_ net392 _2466_ _2472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_165_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4353_ _2419_ _2420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3304_ _1584_ _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4284_ dffram.data\[18\]\[6\] _2369_ _2372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3235_ _1657_ _1670_ _1674_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6023_ _1100_ _1457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_126_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5491__A2 _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _1557_ _1625_ _1627_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3097_ _1563_ _1579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input116_I pdp11_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3254__A1 _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4254__I _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5807_ net23 _1250_ _1234_ net318 _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_3999_ _2167_ _2180_ _2185_ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ net212 _1154_ _1156_ net146 _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input81_I mc14500_sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ _1087_ _1153_ _1157_ _1158_ net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_5_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output502_I net502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A1 _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_81_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__I _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4339__I _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3020_ _1522_ _1523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5630__C1 net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ dffram.data\[41\]\[3\] _2913_ _2917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3922_ _2089_ _2133_ _2135_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_158_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6641_ _0561_ clknet_leaf_136_wb_clk_i wb_sram_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ _2041_ _2082_ _2085_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _0492_ clknet_leaf_107_wb_clk_i dffram.data\[27\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3784_ _1849_ _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_136_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ dffram.data\[17\]\[6\] dffram.data\[19\]\[6\] dffram.data\[21\]\[6\] dffram.data\[23\]\[6\]
+ _0832_ _0834_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput500 net500 io_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput511 net511 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _0954_ _0959_ _0924_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput522 net522 rst_diceroll vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5385_ _0810_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4405_ net421 _2458_ _2459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput533 net533 wbs_dat_o[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput544 net544 wbs_dat_o[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_121_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput555 net555 wbs_dat_o[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4336_ _2405_ _2406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4267_ _1885_ _2265_ _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4198_ _2314_ _2316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3218_ _1663_ _1664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_2_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6006_ _1439_ _1216_ _1441_ _1101_ _1442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_2_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input233_I qcpu_sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3149_ _1574_ _1610_ _1615_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3227__A1 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A1 net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5924__B1 _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__C1 net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output452_I net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3466__A1 _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__A1 _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5915__B1 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5170_ net223 _0679_ _0646_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4121_ dffram.data\[47\]\[7\] _2260_ _2264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4069__I _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _2088_ _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput4 ay8913_do[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3003_ _1453_ _1509_ _1512_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3701__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4957__A1 _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ dffram.data\[42\]\[4\] _2906_ _2907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ dffram.data\[51\]\[3\] _2120_ _2124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4885_ _2704_ _2847_ _2855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3836_ _1433_ _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _0544_ clknet_leaf_125_wb_clk_i wb_counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3767_ _2027_ _2029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6555_ _0475_ clknet_leaf_115_wb_clk_i net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _0963_ _1003_ _1010_ _0980_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA_input183_I qcpu_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _0406_ clknet_leaf_56_wb_clk_i dffram.data\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3698_ _1983_ _1976_ _1984_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input350_I tholin_riscv_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5437_ _0926_ _0943_ net515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_7_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I mc14500_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _0871_ _0874_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4319_ _2349_ _2388_ _2393_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5299_ _0759_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_96_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4707__I _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6184__CLK clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3620__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3439__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3521__I _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A1 net532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4352__I _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ net421 _2655_ _2660_ _2679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3621_ dffram.data\[56\]\[6\] _1930_ _1933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6340_ _0260_ clknet_leaf_27_wb_clk_i dffram.data\[53\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3552_ _1591_ _1885_ _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5116__A1 _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3483_ _1838_ _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6271_ _0191_ clknet_leaf_10_wb_clk_i dffram.data\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ dffram.data\[57\]\[0\] dffram.data\[59\]\[0\] dffram.data\[61\]\[0\] dffram.data\[63\]\[0\]
+ _0729_ _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3678__A1 _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _0661_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4104_ _2252_ _2254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5419__A2 _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5084_ dffram.data\[9\]\[3\] _2986_ _2990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3431__I _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ _2158_ _2206_ _2208_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5986_ _1396_ _1246_ _1422_ net506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_149_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3602__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4937_ net660 _2553_ wb_sram_we _2895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_157_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _2761_ _2841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3819_ _2026_ _2062_ _2064_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _0527_ clknet_leaf_132_wb_clk_i wb_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5294__S _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _2768_ _2786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6538_ _0458_ clknet_leaf_125_wb_clk_i net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_31_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3606__I _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6469_ _0389_ clknet_leaf_14_wb_clk_i dffram.data\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3669__A1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output415_I net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__S1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3841__A1 _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold52_I wbs_adr_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_111_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4085__A1 _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3832__A1 dffram.data\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ net255 _1282_ _1171_ net39 _1301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_158_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5771_ _1237_ _1238_ _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_146_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5178__I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__I _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _2619_ _2721_ _2722_ _2723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 diceroll_do[8] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4653_ wb_counter\[14\] _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_25_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput62 mc14500_do[27] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput51 mc14500_do[17] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput73 mc14500_do[9] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5432__S1 _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3604_ _1921_ _1623_ _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4584_ _2592_ _2602_ _2603_ _2604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
Xinput95 pdp11_do[15] net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3535_ dffram.data\[57\]\[1\] _1874_ _1876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6323_ _0243_ clknet_leaf_19_wb_clk_i dffram.data\[54\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput84 mc14500_sram_in[3] net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_168_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3466_ _1784_ _1823_ _1826_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6254_ _0174_ clknet_leaf_12_wb_clk_i dffram.data\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _0710_ _0714_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__5360__I1 dffram.data\[34\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _0105_ clknet_leaf_72_wb_clk_i dffram.data\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3397_ dffram.data\[28\]\[4\] _1782_ _1783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input146_I pdp11_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5136_ _0648_ _0652_ net520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3161__I _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ dffram.data\[39\]\[4\] _2979_ _2980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5499__S1 _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input313_I tholin_riscv_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _2165_ _2193_ _2197_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__A1 _2033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5969_ net174 _1325_ _1299_ net108 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5576__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5879__A2 _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__S1 _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3336__I _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output532_I net532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput400 net638 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput411 net600 net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5199__S _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3814__A1 _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_104_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__A1 _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__S1 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3320_ dffram.data\[31\]\[2\] _1729_ _1732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3251_ dffram.data\[61\]\[4\] _1684_ _1685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3182_ _1588_ _1631_ _1636_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ net253 _1247_ _1171_ net37 _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_130_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5754_ _1222_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_56_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5636__I _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _1090_ _1170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4705_ _2692_ _2708_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__S1 _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ net535 _2623_ _2626_ _2649_ _2650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5730__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5730__B2 net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _0226_ clknet_leaf_28_wb_clk_i dffram.data\[55\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input263_I sn76489_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4567_ _0637_ _2562_ _2589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3518_ dffram.data\[26\]\[3\] _1861_ _1865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4498_ _1469_ _2528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6237_ _0157_ clknet_leaf_17_wb_clk_i dffram.data\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5371__I _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3449_ _1788_ _1810_ _1815_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _0088_ clknet_leaf_24_wb_clk_i dffram.data\[61\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5119_ design_select\[4\] _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6099_ _0019_ clknet_leaf_75_wb_clk_i dffram.data\[37\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5246__B1 _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4049__A1 _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__B2 net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A1 net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__S0 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A1 _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output482_I net482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4450__I _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__S _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4288__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6029__A2 _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput241 sid_do[14] net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput252 sid_do[5] net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput263 sn76489_do[14] net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput230 qcpu_sram_in[2] net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput296 tholin_riscv_do[14] net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_106_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput285 sn76489_do[9] net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput274 sn76489_do[24] net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_19_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4460__A1 net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__I0 _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A1 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__A1 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ _0726_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4360__I net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ net426 _2470_ _2471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5392__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__A2 _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4352_ _2418_ _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_165_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3303_ _1718_ _1715_ _1719_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_103_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4283_ _2355_ _2368_ _2371_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3234_ dffram.data\[33\]\[6\] _1671_ _1674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6022_ net402 _1440_ _1456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3165_ dffram.data\[63\]\[0\] _1626_ _1627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3096_ _1563_ _1578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input109_I pdp11_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4451__A1 net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1246_ _1263_ _1265_ _1271_ net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_119_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3998_ dffram.data\[29\]\[3\] _2181_ _2185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ net348 _1152_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1092_ _1141_ _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I mc14500_sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5703__A1 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__B2 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4619_ _1523_ _2635_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5599_ _1100_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4442__A1 net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5942__A1 net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__I _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5942__B2 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_143_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4355__I net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4970_ _2526_ _2912_ _2916_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5387__S _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3921_ dffram.data\[19\]\[0\] _2134_ _2135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_158_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _0560_ clknet_leaf_133_wb_clk_i wb_rst_override vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3852_ dffram.data\[52\]\[5\] _2083_ _2085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5933__A1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6571_ _0491_ clknet_leaf_108_wb_clk_i dffram.data\[27\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5933__B2 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5186__I _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5522_ _0944_ _1018_ _1025_ _0961_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_3783_ _2037_ _2038_ _2040_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_4_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_136_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput501 net501 io_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_136_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5453_ _0955_ _0958_ _0879_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput523 net523 rst_hellorld vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput512 net512 qcpu_sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5384_ dffram.data\[16\]\[2\] dffram.data\[18\]\[2\] dffram.data\[20\]\[2\] dffram.data\[22\]\[2\]
+ _0841_ _0842_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput534 net534 wbs_dat_o[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4404_ _2422_ _2458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput545 net545 wbs_dat_o[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3172__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4335_ net370 _2401_ _2404_ _2405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput556 net556 wbs_dat_o[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4266_ _2359_ _2352_ _2360_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4197_ _2314_ _2315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3217_ _1425_ _1662_ _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6005_ net380 _1440_ _1441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_2_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3148_ dffram.data\[0\]\[3\] _1611_ _1615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input226_I qcpu_sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _1563_ _1565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4424__A1 net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5924__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5924__B2 net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output445_I net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4663__A1 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5915__B2 net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__A1 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5734__I _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_114_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__S0 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4120_ _2235_ _2259_ _2263_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _2177_ _2212_ _2217_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput5 ay8913_do[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3002_ dffram.data\[35\]\[1\] _1510_ _1512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4953_ _2898_ _2906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _2098_ _2119_ _2123_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6623_ _0543_ clknet_leaf_124_wb_clk_i wb_counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4884_ _2841_ _2852_ _2853_ _2854_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3835_ _2045_ _2068_ _2073_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3766_ _2027_ _2028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6554_ _0474_ clknet_leaf_115_wb_clk_i net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__3393__A1 _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ _0405_ clknet_leaf_14_wb_clk_i dffram.data\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5505_ _1006_ _1009_ _0905_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5436_ _0774_ _0933_ _0942_ _0792_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_3697_ dffram.data\[55\]\[7\] _1977_ _1984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input176_I qcpu_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3145__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input343_I tholin_riscv_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3164__I _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _0734_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_58_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4318_ dffram.data\[17\]\[3\] _2389_ _2393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5298_ _0757_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_22_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input37_I diceroll_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _2347_ _2342_ _2348_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__B1 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5070__A1 _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_61_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3384__A1 _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output562_I net562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__I _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_76_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5490__S _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__S0 _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_85_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3249__I _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3620_ _1915_ _1929_ _1932_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_133_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3551_ _1754_ _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_12_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_94_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5116__A2 _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3127__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3482_ _1459_ _1838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6270_ _0190_ clknet_leaf_10_wb_clk_i dffram.data\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5221_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5152_ _0631_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4103_ _2252_ _2253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5083_ _2944_ _2985_ _2989_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4627__A1 net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4034_ dffram.data\[4\]\[0\] _2207_ _2208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ net180 _1114_ _1343_ net114 net316 _1219_ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4936_ _0629_ _2510_ _2894_ _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4867_ _2754_ _2840_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input293_I tholin_riscv_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3818_ dffram.data\[22\]\[0\] _2063_ _2064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6606_ _0526_ clknet_leaf_114_wb_clk_i net532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3366__A1 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2998__I _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ net407 _2781_ _2785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6537_ _0457_ clknet_leaf_126_wb_clk_i net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_166_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3749_ _1969_ _2014_ _2017_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _0388_ clknet_leaf_46_wb_clk_i dffram.data\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5419_ _0721_ _0915_ _0925_ _0755_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_6399_ _0319_ clknet_leaf_23_wb_clk_i dffram.data\[59\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4718__I _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__I0 _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5043__A1 _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5751__C1 net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3532__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_128_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4363__I net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5770_ net30 _0627_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5424__I3 dffram.data\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__A1 _1915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4721_ net430 _2705_ _2710_ _2722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _2645_ _2663_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput30 blinker_do[1] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ _1593_ _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_47_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput41 hellorld_do net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput63 mc14500_do[28] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput52 mc14500_do[18] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4583_ _0623_ _2561_ _2603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput96 pdp11_do[16] net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3534_ _1830_ _1873_ _1875_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6322_ _0242_ clknet_leaf_19_wb_clk_i dffram.data\[54\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput85 mc14500_sram_in[4] net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput74 mc14500_sram_addr[0] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3465_ dffram.data\[5\]\[5\] _1824_ _1826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6253_ _0173_ clknet_leaf_13_wb_clk_i dffram.data\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_168_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _0711_ _0712_ _0713_ _0701_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_21_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3396_ _1770_ _1782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6184_ _0104_ clknet_4_12_0_wb_clk_i dffram.data\[32\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5135_ _0651_ _0649_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_97_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input139_I pdp11_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _2971_ _2979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4017_ dffram.data\[49\]\[2\] _2194_ _2197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input306_I tholin_riscv_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ net20 _1400_ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _2741_ _2879_ _2882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5899_ _1344_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3339__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput401 net632 net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput412 wbs_stb_i net412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_output525_I net525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5724__C1 net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3250_ _1676_ _1684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3181_ dffram.data\[63\]\[7\] _1632_ _1636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_163_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5822_ _1245_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5558__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4093__I _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5753_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4821__I _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ net546 _2697_ _2698_ _2707_ _2708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_33_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5684_ _1168_ _1169_ net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_72_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_96_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4635_ _2647_ _2648_ _2649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4566_ _2566_ wb_counter\[3\] _2585_ _2586_ _2587_ _2588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_142_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3517_ _1839_ _1860_ _1864_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6305_ _0225_ clknet_leaf_25_wb_clk_i dffram.data\[55\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3741__A1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4497_ _2526_ _2521_ _2527_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_90_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input256_I sid_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ _0156_ clknet_leaf_44_wb_clk_i dffram.data\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3448_ dffram.data\[60\]\[7\] _1811_ _1815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3379_ _1556_ _1769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4268__I _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _0087_ clknet_leaf_24_wb_clk_i dffram.data\[61\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _0619_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_58_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_139_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6098_ _0018_ clknet_leaf_75_wb_clk_i dffram.data\[37\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5341__S1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5049_ _2952_ _2965_ _2968_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3347__I _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output475_I net475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3082__I _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput220 qcpu_oeb[9] net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_145_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput242 sid_do[15] net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput253 sid_do[6] net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput231 qcpu_sram_in[3] net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput286 tbb1143_do[0] net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput297 tholin_riscv_do[15] net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_106_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput264 sn76489_do[15] net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput275 sn76489_do[25] net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_153_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3971__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ _2408_ _2470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4351_ _1521_ _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_165_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3302_ dffram.data\[32\]\[5\] _1716_ _1719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4282_ dffram.data\[18\]\[5\] _2369_ _2371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3233_ _1655_ _1670_ _1673_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6021_ net83 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_146_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3164_ _1624_ _1626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_143_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_143_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3095_ _1576_ _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _1214_ _1268_ _1270_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3997_ _2165_ _2180_ _2184_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5736_ _1206_ _0663_ _1171_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5667_ net191 _1154_ _1156_ net125 _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input373_I wbs_adr_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4618_ net563 _2623_ _2626_ _2634_ _2635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5703__A2 _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input67_I mc14500_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ _0751_ _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4549_ _2545_ _2571_ _2572_ _2573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_40_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6219_ _0139_ clknet_leaf_70_wb_clk_i dffram.data\[34\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3953__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3705__A1 _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3805__I _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4130__A1 _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__B2 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__A1 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3920_ _2132_ _2134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3851_ _2037_ _2082_ _2084_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6570_ _0490_ clknet_leaf_108_wb_clk_i dffram.data\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3782_ dffram.data\[53\]\[4\] _2039_ _2040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4371__I _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5933__A2 _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5521_ _1021_ _1024_ _0924_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput502 net502 io_out[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5452_ dffram.data\[48\]\[4\] dffram.data\[50\]\[4\] dffram.data\[52\]\[4\] dffram.data\[54\]\[4\]
+ _0956_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_140_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput513 net513 qcpu_sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5383_ dffram.data\[24\]\[2\] dffram.data\[26\]\[2\] dffram.data\[28\]\[2\] dffram.data\[30\]\[2\]
+ _0889_ _0890_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xoutput524 net524 rst_mc14500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4403_ _2454_ net604 _2457_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput535 net535 wbs_dat_o[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput546 net546 wbs_dat_o[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4334_ net372 net371 _2403_ _2404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xoutput557 net557 wbs_dat_o[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_157_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4265_ dffram.data\[16\]\[7\] _2353_ _2360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6004_ _1203_ _1440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_105_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3216_ _1661_ _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4196_ _1608_ _1662_ _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_2_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3147_ _1571_ _1610_ _1614_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input121_I pdp11_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input219_I qcpu_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3078_ _1563_ _1564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_46_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5909__C1 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_40_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__S0 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5719_ _1188_ _1195_ net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5688__B2 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__I _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_123_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output438_I net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4112__A1 _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3360__I _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5463__I1 _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4179__A1 _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3926__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5526__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ dffram.data\[4\]\[7\] _2213_ _2217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput6 ay8913_do[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3001_ _1445_ _1509_ _1511_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3270__I _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__S _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4952_ _2898_ _2905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ dffram.data\[51\]\[2\] _2120_ _2123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5197__I _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _2411_ _2854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _0542_ clknet_leaf_124_wb_clk_i wb_counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3834_ dffram.data\[22\]\[7\] _2069_ _2073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5462__S0 _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3765_ _1526_ _1964_ _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_6_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6553_ _0473_ clknet_leaf_115_wb_clk_i net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_132_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6484_ _0404_ clknet_leaf_47_wb_clk_i dffram.data\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5504_ _1007_ _1008_ _0903_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3696_ _1855_ _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _0936_ _0941_ _0905_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ dffram.data\[57\]\[2\] dffram.data\[59\]\[2\] dffram.data\[61\]\[2\] dffram.data\[63\]\[2\]
+ _0872_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input169_I qcpu_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4317_ _2347_ _2388_ _2392_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5297_ dffram.data\[40\]\[1\] dffram.data\[42\]\[1\] dffram.data\[44\]\[1\] dffram.data\[46\]\[1\]
+ _0804_ _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input336_I tholin_riscv_oeb[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4248_ dffram.data\[16\]\[2\] _2343_ _2348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5842__B2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4179_ _2279_ _2302_ _2304_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3081__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output555_I net555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_131_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5508__S1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5833__B2 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__I _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3090__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_140_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3072__A1 _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_155_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3550_ _1856_ _1879_ _1884_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_12_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3481_ _1836_ _1832_ _1837_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5220_ _0725_ _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5372__I0 _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5151_ _0648_ _0665_ net529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_138_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5082_ dffram.data\[9\]\[2\] _2986_ _2989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4102_ _1542_ _1562_ _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6077__A1 _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4033_ _2205_ _2207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4627__A2 _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5984_ _1396_ _1420_ _1421_ net505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_87_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3063__A1 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4935_ net391 _2509_ _1522_ _2894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _2800_ _2838_ _2839_ _2840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3817_ _2061_ _2063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4797_ wb_counter\[5\] _2783_ _2784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6605_ _0525_ clknet_leaf_115_wb_clk_i net557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input286_I tbb1143_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3748_ dffram.data\[23\]\[1\] _2015_ _2017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _0456_ clknet_leaf_128_wb_clk_i net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_162_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6467_ _0387_ clknet_leaf_48_wb_clk_i dffram.data\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3679_ _1838_ _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5418_ _0918_ _0923_ _0924_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4315__A1 _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _0318_ clknet_leaf_24_wb_clk_i dffram.data\[59\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5349_ _0774_ _0847_ _0857_ _0792_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_54_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6068__A1 net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5815__B2 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_84_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5751__C2 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__B1 _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_111_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4306__A1 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__A1 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__A4 _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3045__A1 _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4720_ wb_counter\[24\] _2721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4651_ net537 _2651_ _2652_ _2662_ _2663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput20 ay8913_do[27] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 blinker_do[2] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3602_ _1919_ _1912_ _1920_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput42 io_in_0 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5742__B1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput64 mc14500_do[29] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput53 mc14500_do[19] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4582_ _2557_ wb_counter\[5\] _2600_ _2601_ _2587_ _2602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xinput97 pdp11_do[17] net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3533_ dffram.data\[57\]\[0\] _1874_ _1875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6321_ _0241_ clknet_leaf_19_wb_clk_i dffram.data\[54\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput86 mc14500_sram_in[5] net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput75 mc14500_sram_addr[1] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6252_ _0172_ clknet_leaf_66_wb_clk_i dffram.data\[26\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3464_ _1780_ _1823_ _1825_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_168_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6183_ _0103_ clknet_leaf_95_wb_clk_i dffram.data\[32\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5203_ net378 _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4819__I _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5134_ _0634_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3395_ _1770_ _1781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5065_ _2971_ _2978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4016_ _2163_ _2193_ _2196_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input201_I qcpu_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5967_ _1386_ _1407_ _1408_ _1409_ net500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_118_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _2864_ _2880_ _2881_ _2871_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input97_I pdp11_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ net264 _1345_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__I _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _2664_ _2822_ _2826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_95_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6519_ _0439_ clknet_leaf_106_wb_clk_i dffram.data\[44\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5336__I0 _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A2 wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput402 net648 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput413 wbs_we_i net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output518_I net518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output420_I net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3275__A1 _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__I net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3180_ _1585_ _1631_ _1635_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_163_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5660__C1 net326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__I _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _1257_ _1281_ _1283_ _1284_ net479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_141_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5752_ _0637_ _0638_ _0640_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4766__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ _2699_ _2704_ _2706_ _2707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5683_ net195 _1163_ _1166_ net129 net331 _1164_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_127_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4634_ net416 _2616_ _2637_ _2648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4518__A1 net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _2502_ _2587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3516_ dffram.data\[26\]\[2\] _1861_ _1864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6304_ _0224_ clknet_leaf_99_wb_clk_i dffram.data\[24\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4496_ dffram.data\[27\]\[2\] _2522_ _2527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input151_I pdp11_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6235_ _0155_ clknet_leaf_44_wb_clk_i dffram.data\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3447_ _1786_ _1810_ _1814_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6166_ _0086_ clknet_leaf_24_wb_clk_i dffram.data\[61\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input249_I sid_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3378_ _1722_ _1763_ _1768_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _0017_ clknet_leaf_80_wb_clk_i dffram.data\[37\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5117_ design_select\[1\] _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_97_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5048_ dffram.data\[38\]\[5\] _2966_ _2968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I ay8913_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_49_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__I _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output468_I net468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__I3 dffram.data\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput210 qcpu_oeb[2] net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_145_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput243 sid_do[16] net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput254 sid_do[7] net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput221 qcpu_sram_addr[0] net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput232 qcpu_sram_in[4] net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput287 tbb1143_do[1] net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput265 sn76489_do[16] net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput276 sn76489_do[26] net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5642__C1 net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput298 tholin_riscv_do[16] net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3248__A1 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5753__I _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4350_ net405 _2409_ _2417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3301_ _1581_ _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_165_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__I _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4281_ _2351_ _2368_ _2370_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6020_ _1436_ _1453_ _1454_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3232_ dffram.data\[33\]\[5\] _1671_ _1673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I ay8913_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _1624_ _1625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_169_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3094_ _1477_ _1576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4987__A1 _2519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ net250 _1269_ _1252_ net34 _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4739__A1 _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ dffram.data\[29\]\[2\] _2181_ _2184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5251__I2 dffram.data\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5666_ _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_143_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input199_I qcpu_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4617_ _2627_ _2628_ _2633_ _2634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input366_I ue1_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ net122 _1097_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ wb_rst_override _2562_ _2572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4279__I _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ net406 _2512_ _2515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6218_ _0138_ clknet_leaf_70_wb_clk_i dffram.data\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _0069_ clknet_leaf_20_wb_clk_i dffram.data\[62\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_5_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4978__A1 _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _2544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_121_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5630__A2 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5748__I _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3850_ dffram.data\[52\]\[4\] _2083_ _2084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_158_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3781_ _2027_ _2039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1022_ _1023_ _0810_ _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__A1 _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5451_ _0743_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput503 net503 io_out[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5697__A2 _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput525 net525 rst_pdp11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput514 net514 qcpu_sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5382_ _0833_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4402_ _2434_ _2457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput536 net536 wbs_dat_o[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput558 net558 wbs_dat_o[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput547 net547 wbs_dat_o[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4333_ net412 net379 _2402_ _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_157_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4264_ _1500_ _2359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5854__C1 net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3215_ _1592_ _1505_ _1661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6003_ net81 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4195_ _2298_ _2308_ _2313_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3731__I _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ dffram.data\[0\]\[2\] _1611_ _1614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3077_ _1559_ _1562_ _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input114_I pdp11_do[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3632__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5909__B1 _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ net205 _1190_ _1193_ net139 net341 _1191_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__S1 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3979_ _2169_ _2170_ _2172_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5649_ net219 _1131_ _1135_ net153 net355 _1133_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5527__I3 dffram.data\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3699__A1 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_142_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output500_I net500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_153_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3816__I _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 ay8913_do[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3000_ dffram.data\[35\]\[0\] _1510_ _1511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3614__A1 _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4951_ _2528_ _2899_ _2904_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3902_ _2095_ _2119_ _2122_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ net393 _2844_ _2853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_138_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6621_ _0541_ clknet_leaf_124_wb_clk_i wb_counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ _2043_ _2068_ _2072_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5462__S1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3764_ _1829_ _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ _0472_ clknet_leaf_116_wb_clk_i net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_125_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _0403_ clknet_leaf_47_wb_clk_i dffram.data\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ dffram.data\[0\]\[5\] dffram.data\[2\]\[5\] dffram.data\[4\]\[5\] dffram.data\[6\]\[5\]
+ _0975_ _0976_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_3695_ _1981_ _1976_ _1982_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5434_ _0939_ _0940_ _0903_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5365_ _0730_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4316_ dffram.data\[17\]\[2\] _2389_ _2392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5296_ _0759_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4247_ _1460_ _2347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3461__I _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input329_I tholin_riscv_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A2 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ dffram.data\[46\]\[0\] _2303_ _2304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input231_I qcpu_sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3853__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ _1595_ _1603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4030__A1 _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output450_I net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__I _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__A1 _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A1 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_133_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3480_ dffram.data\[58\]\[1\] _1833_ _1837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5761__I _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _2942_ _2985_ _2988_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6077__A2 _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4101_ _2237_ _2246_ _2251_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4032_ _2205_ _2206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3835__A1 _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ net179 _1413_ _1097_ net113 _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5588__A1 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4934_ _2892_ _2893_ _2605_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4260__A1 _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ net389 _2763_ _2839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3816_ _2061_ _2062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4796_ _2593_ _2778_ _2783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6604_ _0524_ clknet_leaf_114_wb_clk_i net556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3747_ _1962_ _2014_ _2016_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6535_ _0455_ clknet_leaf_135_wb_clk_i net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_67_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input279_I sn76489_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input181_I qcpu_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6466_ _0386_ clknet_leaf_47_wb_clk_i dffram.data\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3678_ _1969_ _1966_ _1970_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5417_ _0706_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6397_ _0317_ clknet_leaf_23_wb_clk_i dffram.data\[59\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input42_I io_in_0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5348_ _0853_ _0856_ _0708_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6068__A2 _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5815__A2 _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _0784_ _0787_ _0788_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output498_I net498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4003__A1 _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5751__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5751__B2 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4197__I _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_109_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5756__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4650_ _2659_ _2661_ _2662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput10 ay8913_do[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput21 ay8913_do[2] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5742__A1 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3601_ dffram.data\[25\]\[7\] _1913_ _1920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput32 diceroll_do[0] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5742__B2 net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput54 mc14500_do[1] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput43 mc14500_do[0] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4581_ _2425_ _2555_ _2577_ _2601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _0240_ clknet_leaf_145_wb_clk_i dffram.data\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput98 pdp11_do[18] net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput65 mc14500_do[2] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3532_ _1872_ _1874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 mc14500_sram_in[6] net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput76 mc14500_sram_addr[2] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_137_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6251_ _0171_ clknet_leaf_66_wb_clk_i dffram.data\[26\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3463_ dffram.data\[5\]\[4\] _1824_ _1825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6182_ _0102_ clknet_leaf_100_wb_clk_i dffram.data\[32\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5202_ _0686_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_36_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5133_ _0648_ _0650_ net524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_97_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3394_ _1576_ _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_23_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5064_ _2946_ _2972_ _2977_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5353__S0 _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3808__A1 _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ dffram.data\[49\]\[1\] _2194_ _2196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4481__A1 net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5966_ net276 _1322_ _1206_ net61 net309 _1366_ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__4233__A1 _2294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5897_ net242 _1247_ _1264_ net49 _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_8_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4917_ net400 _2866_ _2881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4848_ _2821_ _2823_ _2825_ _2814_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_118_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ _2762_ _2766_ _2767_ _2769_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_67_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6518_ _0438_ clknet_leaf_107_wb_clk_i dffram.data\[44\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6449_ _0369_ clknet_leaf_73_wb_clk_i dffram.data\[47\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput403 net624 net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__B2 net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3096__I _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5575__I1 dffram.data\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ net183 _1154_ _1106_ net319 _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5751_ net236 _1215_ _1218_ net43 net291 _1219_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_72_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ net427 _2705_ _2672_ _2706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_33_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5682_ _1159_ _0671_ _1092_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_72_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4633_ _2621_ _2646_ _2647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _2416_ _2556_ _2577_ _2586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_142_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3515_ _1836_ _1860_ _1863_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6303_ _0223_ clknet_leaf_99_wb_clk_i dffram.data\[24\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6234_ _0154_ clknet_leaf_46_wb_clk_i dffram.data\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4495_ _1460_ _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_90_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3446_ dffram.data\[60\]\[6\] _1811_ _1814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6165_ _0085_ clknet_leaf_24_wb_clk_i dffram.data\[61\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3377_ dffram.data\[2\]\[7\] _1764_ _1768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input144_I pdp11_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5116_ _0632_ _0636_ net527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5326__S0 _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _0016_ clknet_leaf_113_wb_clk_i wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5047_ _2948_ _2965_ _2967_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input311_I tholin_riscv_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4454__A1 net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4206__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5949_ _1245_ _1393_ _1394_ _1395_ net496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_66_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output530_I net530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput211 qcpu_oeb[30] net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput200 qcpu_oeb[20] net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput244 sid_do[17] net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput222 qcpu_sram_addr[1] net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput233 qcpu_sram_in[5] net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput288 tbb1143_do[2] net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput255 sid_do[8] net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput266 sn76489_do[17] net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput277 sn76489_do[27] net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4475__I _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput299 tholin_riscv_do[17] net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_106_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__A1 net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3554__I _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3300_ _1714_ _1715_ _1717_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_165_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4280_ dffram.data\[18\]\[4\] _2369_ _2370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3231_ _1651_ _1670_ _1672_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3162_ _1562_ _1623_ _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4385__I _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3093_ _1574_ _1564_ _1575_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4436__A1 net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5803_ _1086_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5936__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ _2163_ _2180_ _2183_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _1204_ _1205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5251__I3 dffram.data\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5665_ _1094_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ net444 _2629_ _2632_ _2633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5596_ _0671_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input261_I sn76489_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _2566_ _2567_ _2569_ _2570_ _2559_ _2571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_input359_I ue1_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4478_ _0633_ _2505_ _2513_ _2514_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6217_ _0137_ clknet_leaf_70_wb_clk_i dffram.data\[34\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3429_ _1434_ _1623_ _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6148_ _0068_ clknet_leaf_37_wb_clk_i dffram.data\[62\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4675__A1 net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _1506_ _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_73_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__A1 net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5927__A1 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5927__B2 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output480_I net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3166__A1 _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_160_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold13_I wbs_dat_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5091__A1 _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_158_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3780_ _2027_ _2038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _0826_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_136_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3157__A1 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ net386 _2455_ _2456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput504 net504 io_out[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput515 net515 qcpu_sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3284__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput526 net526 rst_qcpu vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5381_ _0831_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput559 net559 wbs_dat_o[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput537 net537 wbs_dat_o[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput548 net548 wbs_dat_o[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4332_ wb_feedback_delay _2402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4263_ _2357_ _2352_ _2358_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5854__C2 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5854__B1 _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3214_ _1659_ _1652_ _1660_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6002_ _1437_ _1438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4194_ dffram.data\[46\]\[7\] _2309_ _2313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3145_ _1568_ _1610_ _1613_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4409__A1 net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3076_ _1561_ _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__I _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input107_I pdp11_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5909__B2 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5909__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ dffram.data\[50\]\[4\] _2171_ _2172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5717_ _1188_ _1194_ net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5674__I _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _0617_ clknet_leaf_57_wb_clk_i dffram.data\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5648_ _0642_ _0658_ _1139_ _1140_ _1141_ _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input72_I mc14500_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _1079_ _1081_ _1062_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_142_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_0_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3369__I _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3387__A1 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__A1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4887__A1 net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 ay8913_do[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__A1 _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4950_ dffram.data\[42\]\[3\] _2900_ _2904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3901_ dffram.data\[51\]\[1\] _2120_ _2122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4881_ wb_counter\[21\] _2847_ _2852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_28_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3832_ dffram.data\[22\]\[6\] _2069_ _2072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6620_ _0540_ clknet_leaf_124_wb_clk_i wb_counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3378__A1 _1722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__B1 _2594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6551_ _0471_ clknet_leaf_117_wb_clk_i net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_41_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5502_ dffram.data\[8\]\[5\] dffram.data\[10\]\[5\] dffram.data\[12\]\[5\] dffram.data\[14\]\[5\]
+ _0937_ _0938_ _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3763_ _1983_ _2020_ _2025_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6482_ _0402_ clknet_leaf_67_wb_clk_i dffram.data\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3694_ dffram.data\[55\]\[6\] _1977_ _1982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5433_ dffram.data\[0\]\[3\] dffram.data\[2\]\[3\] dffram.data\[4\]\[3\] dffram.data\[6\]\[3\]
+ _0785_ _0786_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_112_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _0738_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4315_ _2345_ _2388_ _2391_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3550__A1 _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5295_ _0794_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_39_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4246_ _2345_ _2342_ _2346_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4177_ _2301_ _2303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3128_ _1595_ _1602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input224_I qcpu_sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3059_ _1470_ _1544_ _1549_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3189__I _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__B1 _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output443_I net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5597__A2 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_116_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3827__I _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_133_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5080_ dffram.data\[9\]\[1\] _2986_ _2988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4100_ dffram.data\[14\]\[7\] _2247_ _2251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4031_ _2074_ _1559_ _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5037__A1 _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5982_ net315 _1152_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5588__A2 _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3599__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ net380 _2510_ _2893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_72_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4864_ wb_counter\[18\] _2834_ _2838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_59_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3815_ _1740_ _2012_ _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4795_ _2777_ _2779_ _2782_ _2769_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6603_ _0523_ clknet_leaf_114_wb_clk_i net554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3746_ dffram.data\[23\]\[0\] _2015_ _2016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6534_ _0454_ clknet_leaf_136_wb_clk_i net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6465_ _0385_ clknet_leaf_66_wb_clk_i dffram.data\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5416_ _0921_ _0922_ _0879_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3677_ dffram.data\[55\]\[1\] _1967_ _1970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input174_I qcpu_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ _0316_ clknet_leaf_32_wb_clk_i dffram.data\[59\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_81_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5347_ _0854_ _0855_ _0788_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3523__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input341_I tholin_riscv_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _0746_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_54_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input35_I diceroll_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4229_ _2327_ _2335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_90_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5200__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__I _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5751__A2 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output560_I net560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3762__A1 dffram.data\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3382__I _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5303__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 ay8913_do[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 ay8913_do[3] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _0996_ _1011_ _2552_ _2600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3600_ _1855_ _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput33 diceroll_do[1] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5742__A2 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput55 mc14500_do[20] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput44 mc14500_do[10] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3531_ _1872_ _1873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3753__A1 _1973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput66 mc14500_do[30] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput88 mc14500_sram_in[7] net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput77 mc14500_sram_addr[3] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput99 pdp11_do[19] net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_161_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6250_ _0170_ clknet_leaf_66_wb_clk_i dffram.data\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3462_ _1816_ _1824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3393_ _1778_ _1771_ _1779_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6181_ _0101_ clknet_leaf_109_wb_clk_i dffram.data\[32\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5201_ net79 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5132_ _0618_ net578 _0649_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xclkbuf_leaf_106_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5063_ dffram.data\[39\]\[3\] _2973_ _2977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5353__S1 _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4014_ _2158_ _2193_ _2195_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4481__A2 _2504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ net173 _1325_ _1299_ net107 _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5966__C1 net309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5896_ net161 _1262_ _1326_ net7 _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4916_ _2741_ _2879_ _2880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_168_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5718__C1 net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ net385 _2824_ _2825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input291_I tholin_riscv_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_95_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _2768_ _2769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3729_ dffram.data\[54\]\[3\] _2000_ _2004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6517_ _0437_ clknet_leaf_107_wb_clk_i dffram.data\[44\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6448_ _0368_ clknet_leaf_145_wb_clk_i dffram.data\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6379_ _0299_ clknet_leaf_26_wb_clk_i dffram.data\[51\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput404 net627 net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3930__I _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5709__C1 net338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold43_I wbs_dat_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4001__I _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5660__A1 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5660__B2 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5750_ _1117_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_147_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5681_ _1160_ _1167_ net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__3974__A1 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4701_ _2614_ _2705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4632_ wb_counter\[11\] _2646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3726__A1 _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4563_ _0926_ _0943_ _2568_ _2585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_64_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3514_ dffram.data\[26\]\[1\] _1861_ _1863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4494_ _2524_ _2521_ _2525_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6302_ _0222_ clknet_leaf_99_wb_clk_i dffram.data\[24\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6233_ _0153_ clknet_leaf_46_wb_clk_i dffram.data\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3445_ _1784_ _1810_ _1813_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5007__I _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6164_ _0084_ clknet_leaf_34_wb_clk_i dffram.data\[61\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3376_ _1720_ _1763_ _1767_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5326__S1 _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6095_ _0015_ clknet_leaf_87_wb_clk_i dffram.data\[35\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4846__I _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input137_I pdp11_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5046_ dffram.data\[38\]\[4\] _2966_ _2967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input304_I tholin_riscv_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5948_ net305 _1127_ _1363_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xclkbuf_leaf_74_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_66_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__A1 _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5879_ net262 _1287_ _1334_ net93 _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_146_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3717__A1 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4390__A1 net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A1 _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput201 qcpu_oeb[21] net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_145_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output523_I net523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput212 qcpu_oeb[31] net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput245 sid_do[18] net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput223 qcpu_sram_addr[2] net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput234 qcpu_sram_in[6] net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput256 sid_do[9] net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput278 sn76489_do[2] net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput267 sn76489_do[18] net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5642__B2 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__A1 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput289 tbb1143_do[3] net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_106_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_86_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A1 net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3230_ dffram.data\[33\]\[4\] _1671_ _1672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5881__B2 net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ _1622_ _1623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3092_ dffram.data\[7\]\[3\] _1565_ _1575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5802_ net22 _1266_ _1267_ net115 _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3994_ dffram.data\[29\]\[1\] _2181_ _2183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3947__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5492__S0 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5664_ _1102_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_143_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5595_ _1096_ _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3745__I _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4615_ _2631_ _2632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4546_ _2413_ _2556_ _2557_ _2570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_121_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_29_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4477_ _2419_ _2514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4124__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input254_I sid_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3428_ _1788_ _1797_ _1802_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6216_ _0136_ clknet_leaf_98_wb_clk_i dffram.data\[28\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5872__A1 net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _0067_ clknet_leaf_36_wb_clk_i dffram.data\[62\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3359_ _1756_ _1757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_5_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _1504_ _1505_ _1506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5029_ _2954_ _2949_ _2955_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5927__A2 _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3938__A1 _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output473_I net473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__I _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__A1 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__B2 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5311__S _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5110__I _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_138_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4400_ _2431_ _2455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput505 net505 io_out[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_164_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput516 net516 qcpu_sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5380_ _0886_ _0887_ _0836_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput527 net527 rst_sid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput538 net538 wbs_dat_o[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4331_ net413 _2401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput549 net549 wbs_dat_o[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_120_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4106__A1 _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ dffram.data\[16\]\[6\] _2353_ _2358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5854__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5854__B2 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3213_ dffram.data\[62\]\[7\] _1653_ _1660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1100_ _1437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4193_ _2296_ _2308_ _2312_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3144_ dffram.data\[0\]\[1\] _1611_ _1613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_2_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3075_ _1560_ _1505_ _1561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__A1 _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__I _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__S0 _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3977_ _2159_ _2171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5716_ net204 _1190_ _1193_ net138 net340 _1191_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6696_ _0616_ clknet_leaf_98_wb_clk_i dffram.data\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_21_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5647_ net436 _0641_ _0636_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_116_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3475__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4345__A1 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input65_I mc14500_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5578_ _1057_ _1080_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4529_ _0756_ _0793_ _2553_ _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_111_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_142_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A1 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5781__B1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_101_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3139__A2 _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5306__S _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__A1 net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__A4 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput9 ay8913_do[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4811__A2 _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _2089_ _2119_ _2121_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _2846_ _2849_ _2851_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_28_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5447__S0 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3831_ _2041_ _2068_ _2071_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6550_ _0470_ clknet_leaf_117_wb_clk_i net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3762_ dffram.data\[23\]\[7\] _2021_ _2025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_41_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5501_ _1004_ _1005_ _0788_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_41_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6481_ _0401_ clknet_leaf_47_wb_clk_i dffram.data\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3693_ _1852_ _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5432_ dffram.data\[8\]\[3\] dffram.data\[10\]\[3\] dffram.data\[12\]\[3\] dffram.data\[14\]\[3\]
+ _0937_ _0938_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4327__A1 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ dffram.data\[49\]\[2\] dffram.data\[51\]\[2\] dffram.data\[53\]\[2\] dffram.data\[55\]\[2\]
+ _0816_ _0817_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_168_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ dffram.data\[17\]\[1\] _2389_ _2391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5827__B2 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5827__A1 net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5294_ _0798_ _0801_ _0802_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4245_ dffram.data\[16\]\[1\] _2343_ _2346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4176_ _2301_ _2302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3127_ _1574_ _1596_ _1601_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input217_I qcpu_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3058_ dffram.data\[43\]\[3\] _1545_ _1549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__I _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__B1 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6679_ _0599_ clknet_leaf_95_wb_clk_i dffram.data\[38\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output436_I net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3057__A1 _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4557__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4309__A1 _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__B1 _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4030_ _2177_ _2199_ _2204_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5981_ _1387_ _1418_ _1419_ net504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4932_ wb_override_act _2512_ _2892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4863_ _2821_ _2836_ _2837_ _2829_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6602_ _0522_ clknet_leaf_114_wb_clk_i net553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3814_ _2045_ _2055_ _2060_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4794_ net406 _2781_ _2782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3745_ _2013_ _2015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _0453_ clknet_leaf_136_wb_clk_i net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_125_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _0384_ clknet_leaf_137_wb_clk_i dffram.data\[20\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3676_ _1835_ _1969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5415_ dffram.data\[48\]\[3\] dffram.data\[50\]\[3\] dffram.data\[52\]\[3\] dffram.data\[54\]\[3\]
+ _0742_ _0744_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_63_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6395_ _0315_ clknet_leaf_27_wb_clk_i dffram.data\[59\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_28_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5346_ dffram.data\[0\]\[1\] dffram.data\[2\]\[1\] dffram.data\[4\]\[1\] dffram.data\[6\]\[1\]
+ _0785_ _0786_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_input167_I qcpu_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5277_ dffram.data\[0\]\[0\] dffram.data\[2\]\[0\] dffram.data\[4\]\[0\] dffram.data\[6\]\[0\]
+ _0785_ _0786_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_54_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input334_I tholin_riscv_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4228_ _2327_ _2334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input28_I ay8913_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4159_ _2288_ _2281_ _2289_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3039__A1 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3211__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5672__C1 net328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3278__A1 dffram.data\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3838__I _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3450__A1 _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput12 ay8913_do[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 diceroll_do[2] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput23 ay8913_do[4] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput45 mc14500_do[11] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3530_ _1638_ _1662_ _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput89 pdp11_do[0] net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput56 mc14500_do[21] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput67 mc14500_do[3] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput78 mc14500_sram_addr[4] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3461_ _1816_ _1823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3392_ dffram.data\[28\]\[3\] _1772_ _1779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6180_ _0100_ clknet_leaf_71_wb_clk_i dffram.data\[32\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5200_ net226 _0701_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_21_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4702__A1 net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5131_ _0643_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5062_ _2944_ _2972_ _2976_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3269__A1 _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ dffram.data\[49\]\[0\] _2194_ _2195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_146_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_133_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ net19 _1400_ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5966__C2 _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5895_ net366 _1111_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4915_ _2721_ _2735_ _2858_ _2873_ _2879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _2780_ _2824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5194__A1 net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6516_ _0436_ clknet_leaf_93_wb_clk_i dffram.data\[44\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input284_I sn76489_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4777_ _1521_ _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3728_ _1971_ _1999_ _2003_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3659_ _1949_ _1957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6447_ _0367_ clknet_leaf_145_wb_clk_i dffram.data\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6378_ _0298_ clknet_leaf_26_wb_clk_i dffram.data\[51\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5329_ _0831_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput405 net652 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5654__C1 net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5957__B1 _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3658__I _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5575__I3 dffram.data\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4489__I _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3499__A1 _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__S _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4999__A1 _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3671__A1 _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4952__I _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5963__A3 _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5680_ net194 _1163_ _1166_ net128 net330 _1164_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_85_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ wb_counter\[21\] _2704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_155_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1522_ _2645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5783__I _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4562_ net558 _2583_ _2584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3513_ _1830_ _1860_ _1862_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4493_ dffram.data\[27\]\[1\] _2522_ _2525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _0221_ clknet_leaf_99_wb_clk_i dffram.data\[24\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3444_ dffram.data\[60\]\[5\] _1811_ _1813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6232_ _0152_ clknet_leaf_16_wb_clk_i dffram.data\[60\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6163_ _0083_ clknet_leaf_34_wb_clk_i dffram.data\[61\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3375_ dffram.data\[2\]\[6\] _1764_ _1767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _0625_ _0634_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_104_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6094_ _0014_ clknet_leaf_86_wb_clk_i dffram.data\[35\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5045_ _2958_ _2966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5947_ net272 _1322_ _1114_ net169 net57 _1206_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__3414__A1 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3478__I _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input95_I pdp11_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _1155_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_43_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ net381 _2800_ _2810_ _2811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput202 qcpu_oeb[22] net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3941__I _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput213 qcpu_oeb[32] net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput224 qcpu_sram_addr[3] net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput235 qcpu_sram_in[7] net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output516_I net516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput257 sid_oeb net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput246 sid_do[19] net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput279 sn76489_do[3] net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput268 sn76489_do[19] net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_106_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__I _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3653__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__I _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__B1 net519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5158__A1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4012__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3160_ _1540_ _0754_ _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5618__C1 net335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3091_ _1573_ _1574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold1 wbs_dat_i[10] net581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5633__A2 _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3644__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5801_ _1095_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3298__I _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_138_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3993_ _2158_ _2180_ _2182_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5732_ _0712_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5492__S1 _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_44_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5663_ net327 _1152_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_115_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5594_ _1095_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4614_ _2630_ _2631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4545_ _0825_ _0858_ _2568_ _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_142_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_147_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ net405 _2512_ _2513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3427_ dffram.data\[34\]\[7\] _1798_ _1802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6215_ _0135_ clknet_leaf_98_wb_clk_i dffram.data\[28\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6146_ _0066_ clknet_leaf_36_wb_clk_i dffram.data\[62\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3358_ _1608_ _1755_ _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input247_I sid_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3289_ _1708_ _1705_ _1709_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6077_ _0702_ _0705_ _1431_ _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input10_I ay8913_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ dffram.data\[3\]\[6\] _2950_ _2955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_156_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4060__A1 _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output466_I net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_165_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5863__A2 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__A1 _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A1 _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__B _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput506 net506 io_out[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput517 net517 qcpu_sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput528 net528 rst_sn76489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput539 net539 wbs_dat_o[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4330_ net414 _2400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4261_ _1493_ _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _1435_ _1436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3212_ _1587_ _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input2_I ay8913_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ dffram.data\[46\]\[6\] _2309_ _2312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3143_ _1557_ _1610_ _1612_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_2_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3074_ _0827_ _0829_ _1560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5301__I _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_46_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5465__S1 _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3976_ _2159_ _2170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5790__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5715_ _1177_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6695_ _0615_ clknet_leaf_98_wb_clk_i dffram.data\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5646_ net436 _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA_input197_I qcpu_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_21_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ dffram.data\[16\]\[7\] dffram.data\[18\]\[7\] dffram.data\[20\]\[7\] dffram.data\[22\]\[7\]
+ _0956_ _0957_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input364_I ue1_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4528_ _2552_ _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I mc14500_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4459_ _2497_ net625 _2491_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_142_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6129_ _0049_ clknet_leaf_35_wb_clk_i dffram.data\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3608__A1 _1899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4281__A1 _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5781__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5781__B2 net313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__A1 _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3075__A2 _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5447__S1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4024__A1 _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3830_ dffram.data\[22\]\[5\] _2069_ _2071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5772__A1 net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3761_ _1981_ _2020_ _2024_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5772__B2 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3576__I _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ dffram.data\[1\]\[5\] dffram.data\[3\]\[5\] dffram.data\[5\]\[5\] dffram.data\[7\]\[5\]
+ _0897_ _0898_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _0400_ clknet_leaf_109_wb_clk_i dffram.data\[46\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3692_ _1979_ _1976_ _1980_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _0777_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _0864_ _0869_ _0814_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _2340_ _2388_ _2390_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5827__A2 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5293_ _0692_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_22_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5383__S0 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4244_ _1452_ _2345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ _2300_ _1640_ _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3126_ dffram.data\[8\]\[3\] _1597_ _1601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input112_I pdp11_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3057_ _1461_ _1544_ _1548_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4263__A1 _2357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5763__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5763__B2 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3486__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _2115_ _2152_ _2157_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6678_ _0598_ clknet_leaf_94_wb_clk_i dffram.data\[38\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5629_ _1120_ _1128_ net476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_103_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3829__A1 _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output429_I net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3396__I _1770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5980_ net66 _1218_ _1343_ net112 net314 _1118_ _1419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_91_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A1 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ _2846_ _2890_ _2891_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_87_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ net388 _2824_ _2837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3813_ dffram.data\[13\]\[7\] _2056_ _2060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6601_ _0521_ clknet_leaf_114_wb_clk_i net552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5745__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4793_ _2780_ _2781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3744_ _2013_ _2014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6532_ _0452_ clknet_leaf_137_wb_clk_i net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_141_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3675_ _1962_ _1966_ _1968_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6463_ _0383_ clknet_leaf_139_wb_clk_i dffram.data\[20\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ dffram.data\[56\]\[3\] dffram.data\[58\]\[3\] dffram.data\[60\]\[3\] dffram.data\[62\]\[3\]
+ _0919_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5227__S _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _0314_ clknet_leaf_33_wb_clk_i dffram.data\[59\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5345_ dffram.data\[8\]\[1\] dffram.data\[10\]\[1\] dffram.data\[12\]\[1\] dffram.data\[14\]\[1\]
+ _0782_ _0783_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5276_ _0726_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_68_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4227_ _2288_ _2328_ _2333_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5520__I1 _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input327_I tholin_riscv_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__A1 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4158_ dffram.data\[15\]\[3\] _2282_ _2289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _2225_ _2240_ _2244_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ _1587_ _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4227__A1 _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3450__A2 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 ay8913_do[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 diceroll_do[3] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput24 ay8913_do[5] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 mc14500_do[12] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput57 mc14500_do[22] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput68 mc14500_do[4] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput79 mc14500_sram_addr[5] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3460_ _1778_ _1817_ _1822_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3391_ _1573_ _1778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ _0631_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_122_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5061_ dffram.data\[39\]\[2\] _2973_ _2976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4012_ _2192_ _2194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5510__S _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _1386_ _1404_ _1405_ _1406_ net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5966__A1 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5966__B2 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4914_ _2864_ _2877_ _2878_ _2871_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5894_ _1340_ _1341_ _1342_ _1348_ net488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5718__A1 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5718__B2 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4845_ wb_counter\[14\] _2822_ _2823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_16_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_115_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_145_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4776_ net391 _2764_ _2767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_95_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6515_ _0435_ clknet_leaf_93_wb_clk_i dffram.data\[44\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3727_ dffram.data\[54\]\[2\] _2000_ _2003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__A2 _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3658_ _1949_ _1956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__S0 _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input277_I sn76489_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6446_ _0366_ clknet_leaf_145_wb_clk_i dffram.data\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6377_ _0297_ clknet_leaf_26_wb_clk_i dffram.data\[51\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_73_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3589_ _1844_ _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5328_ _0830_ _0835_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input40_I diceroll_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput406 net650 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4595__I net562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _0692_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4457__A1 net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A1 net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output496_I net496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__B2 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__A1 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__S0 _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_167_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__B1 _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4696__A1 net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3849__I _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4620__A1 _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__A4 _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4630_ _1523_ _2644_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6300_ _0220_ clknet_leaf_65_wb_clk_i dffram.data\[24\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4561_ _2582_ _2583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3512_ dffram.data\[26\]\[0\] _1861_ _1862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _1452_ _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6231_ _0151_ clknet_leaf_15_wb_clk_i dffram.data\[60\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3443_ _1780_ _1810_ _1812_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _0082_ clknet_leaf_34_wb_clk_i dffram.data\[61\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__S _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3374_ _1718_ _1763_ _1766_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_51_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ design_select\[4\] _0633_ _0618_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_139_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ _0013_ clknet_leaf_86_wb_clk_i dffram.data\[35\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5304__I _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A1 net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _2958_ _2965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3111__A1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5240__S _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5946_ net15 _1312_ _1116_ net103 _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_66_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5877_ net159 _1325_ _1326_ net5 _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_91_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4828_ _2796_ _2806_ _2809_ _2810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_29_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3178__A1 _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input88_I mc14500_sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4759_ _2734_ _2753_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_83_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6429_ _0349_ clknet_leaf_5_wb_clk_i dffram.data\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_12_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput203 qcpu_oeb[23] net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput214 qcpu_oeb[3] net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput236 sid_do[0] net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput225 qcpu_sram_addr[4] net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput247 sid_do[1] net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput269 sn76489_do[1] net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput258 sn76489_do[0] net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output509_I net509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4850__A1 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A1 net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3341__A1 _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3090_ _1468_ _1573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold2 net620 net579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4963__I _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__A1 net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5800_ _1224_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3992_ dffram.data\[29\]\[0\] _2181_ _2182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5731_ _1186_ _1202_ net471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5662_ _1132_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5593_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4613_ _2546_ _2551_ _2630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4544_ _2552_ _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5857__B1 _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6214_ _0134_ clknet_leaf_98_wb_clk_i dffram.data\[28\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4475_ _2504_ _2512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3426_ _1786_ _1797_ _1801_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5034__I _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6145_ _0065_ clknet_leaf_37_wb_clk_i dffram.data\[62\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3357_ _1754_ _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input142_I pdp11_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _0827_ _1503_ _1504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3288_ dffram.data\[32\]\[1\] _1706_ _1709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5085__A1 _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _1493_ _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_68_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_130_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_130_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5929_ _1377_ _1378_ _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4113__I _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__A1 net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_8_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output459_I net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3323__A1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold96_I wbs_dat_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput507 net507 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput518 net518 qcpu_sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3562__A1 _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5839__B1 _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput529 net529 rst_tbb1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3862__I _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4260_ _2355_ _2352_ _2356_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3211_ _1657_ _1652_ _1658_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _2294_ _2308_ _2311_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3142_ dffram.data\[0\]\[0\] _1611_ _1612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3073_ _1558_ _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A1 _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3975_ _2103_ _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5790__A2 _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _1188_ _1192_ net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_116_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6694_ _0614_ clknet_leaf_57_wb_clk_i dffram.data\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _1138_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_61_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _0844_ _1078_ _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4868__I _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _2551_ _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input357_I ue1_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4458_ net403 _2489_ _2498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3409_ _1790_ _1791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_142_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _0048_ clknet_leaf_12_wb_clk_i dffram.data\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4389_ _2422_ _2447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5058__A1 _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ net87 _1489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_139_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3792__A1 _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3544__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4778__I _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_131_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__A1 _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4811__A4 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3760_ dffram.data\[23\]\[6\] _2021_ _2024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3783__A1 _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _0781_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3691_ dffram.data\[55\]\[5\] _1977_ _1980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _0867_ _0868_ _0811_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5292_ dffram.data\[33\]\[1\] dffram.data\[35\]\[1\] dffram.data\[37\]\[1\] dffram.data\[39\]\[1\]
+ _0799_ _0800_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_4312_ dffram.data\[17\]\[0\] _2389_ _2390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4243_ _2340_ _2342_ _2344_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_39_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5383__S1 _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5513__S _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _1541_ _2300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3125_ _1571_ _1596_ _1600_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3056_ dffram.data\[43\]\[2\] _1545_ _1548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input105_I pdp11_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3767__I _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3958_ dffram.data\[59\]\[7\] _2153_ _2157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6677_ _0597_ clknet_leaf_71_wb_clk_i dffram.data\[38\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3889_ dffram.data\[21\]\[6\] _2106_ _2113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5628_ net210 _1122_ _1124_ net144 net346 _1127_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_131_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input70_I mc14500_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5920__C1 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3526__A1 dffram.data\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ _0706_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_113_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__A1 net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3765__A1 _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3517__A1 _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ net404 _2850_ _2891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _2834_ _2835_ _2836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_157_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3812_ _2043_ _2055_ _2059_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6600_ _0520_ clknet_leaf_119_wb_clk_i net551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5745__A2 _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4792_ _2760_ _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3743_ _1724_ _2012_ _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_82_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6531_ _0451_ clknet_leaf_137_wb_clk_i net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XPHY_EDGE_ROW_41_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3674_ dffram.data\[55\]\[0\] _1967_ _1968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6462_ _0382_ clknet_leaf_137_wb_clk_i dffram.data\[20\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6393_ _0313_ clknet_leaf_33_wb_clk_i dffram.data\[59\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5413_ _0730_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5344_ _0850_ _0851_ _0852_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4181__A1 _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5275_ _0781_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_54_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4226_ dffram.data\[45\]\[3\] _2329_ _2333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4157_ _2100_ _2288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_71_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3108_ _1499_ _1587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input222_I qcpu_sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4088_ dffram.data\[14\]\[2\] _2241_ _2244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3039_ _1479_ _1534_ _1536_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3995__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__S0 _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3747__A1 _1962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5418__S _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_150_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5217__I _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output441_I net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5672__A1 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__B2 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6048__I _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_147_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5975__A2 _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5328__S _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3738__A1 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 ay8913_do[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput25 ay8913_do[6] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput36 diceroll_do[4] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput58 mc14500_do[23] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput47 mc14500_do[13] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput69 mc14500_do[5] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_123_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3390_ _1776_ _1771_ _1777_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3910__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5060_ _2942_ _2972_ _2975_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A1 net327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _2192_ _2193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ net275 _1278_ _1370_ net60 net308 _1357_ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4913_ net399 _2866_ _2878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ net94 _1343_ _1219_ net296 _1347_ _1348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ wb_counter\[11\] wb_counter\[12\] wb_counter\[13\] _2808_ _2822_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5274__S0 _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4775_ _2549_ _2567_ _2766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_99_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5238__S _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3726_ _1969_ _1999_ _2002_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6514_ _0434_ clknet_leaf_93_wb_clk_i dffram.data\[44\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3657_ _1909_ _1950_ _1955_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__S1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input172_I qcpu_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _0365_ clknet_leaf_145_wb_clk_i dffram.data\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3588_ _1909_ _1902_ _1910_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _0296_ clknet_leaf_143_wb_clk_i dffram.data\[21\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _0735_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3780__I _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput407 net649 net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input33_I diceroll_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__B2 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A1 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ dffram.data\[16\]\[0\] dffram.data\[18\]\[0\] dffram.data\[20\]\[0\] dffram.data\[22\]\[0\]
+ _0762_ _0763_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5189_ _0695_ _0698_ _0693_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4209_ dffram.data\[1\]\[4\] _2322_ _2323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__A1 _2163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__I _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output489_I net489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5265__S0 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4393__A1 net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5568__S1 _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__B2 net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_141_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3959__A1 _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3865__I _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3187__A2 _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A1 net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ _2541_ _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_7_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3511_ _1859_ _1861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4491_ _2519_ _2521_ _2523_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6230_ _0150_ clknet_leaf_15_wb_clk_i dffram.data\[60\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3442_ dffram.data\[60\]\[4\] _1811_ _1812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6161_ _0081_ clknet_leaf_34_wb_clk_i dffram.data\[61\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3373_ dffram.data\[2\]\[5\] _1764_ _1766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ design_select\[1\] _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6092_ _0012_ clknet_leaf_87_wb_clk_i dffram.data\[35\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5043_ _2946_ _2959_ _2964_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5521__S _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5320__I _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__S0 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5945_ _1387_ _1388_ _1392_ net495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5876_ _1285_ _1327_ _1328_ _1332_ net486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_66_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__B _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4827_ _2808_ _2809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__A1 net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ net556 _2739_ _2740_ _2752_ _2753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3709_ _1973_ _1986_ _1991_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ _2627_ _2693_ _2694_ _2695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6428_ _0348_ clknet_leaf_34_wb_clk_i dffram.data\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5875__A1 net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6359_ _0279_ clknet_leaf_142_wb_clk_i dffram.data\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput204 qcpu_oeb[24] net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput215 qcpu_oeb[4] net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput226 qcpu_sram_addr[5] net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_162_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput248 sid_do[20] net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput237 sid_do[10] net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_76_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput259 sn76489_do[10] net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_162_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6052__A1 net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__A2 _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4366__A1 net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__A1 _2233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__S0 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A1 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5618__B2 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold3 _2449_ net580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_18_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__I _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6043__A1 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3991_ _2179_ _2181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5477__S0 _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5730_ net211 _1197_ _1183_ net145 net347 _1198_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_85_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _1148_ _1151_ net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_128_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5592_ _0619_ net578 _0661_ _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_128_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4612_ _2614_ _2629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ wb_counter\[1\] _2567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5857__B2 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5857__A1 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5401__S0 _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ _0133_ clknet_leaf_98_wb_clk_i dffram.data\[28\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _2506_ _2511_ _2501_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3425_ dffram.data\[34\]\[6\] _1798_ _1801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3356_ _1504_ _1432_ _1754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6144_ _0064_ clknet_leaf_22_wb_clk_i dffram.data\[63\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3287_ _1567_ _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6075_ _0829_ _1503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input135_I pdp11_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5026_ _2952_ _2949_ _2953_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_68_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input302_I tholin_riscv_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6034__A1 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5468__S0 _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ net165 _1365_ _1366_ net301 _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_119_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5859_ net361 _1111_ _1239_ _1317_ _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_119_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4348__A1 _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__S _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5848__A1 net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5225__I _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_160_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output521_I net521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__S0 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_88_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4587__A1 net561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold89_I wbs_dat_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_136_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3011__A1 _1479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput508 net508 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__5336__S _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput519 net519 qcpu_sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_97_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3210_ dffram.data\[62\]\[6\] _1653_ _1658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4190_ dffram.data\[46\]\[5\] _2309_ _2311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4511__A1 _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3141_ _1609_ _1611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4974__I _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3072_ _1423_ _0980_ _1558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3974_ _2167_ _2160_ _2168_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_63_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5713_ net203 _1190_ _1178_ net137 net339 _1191_ _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6693_ _0613_ clknet_leaf_66_wb_clk_i dffram.data\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ _0651_ _0649_ _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ dffram.data\[24\]\[7\] dffram.data\[26\]\[7\] dffram.data\[28\]\[7\] dffram.data\[30\]\[7\]
+ _1058_ _1059_ _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4526_ _2550_ net369 _2551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4750__A1 _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5045__I _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4457_ net437 _2492_ _2497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3408_ _1703_ _1755_ _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_input252_I sid_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6127_ _0047_ clknet_leaf_10_wb_clk_i dffram.data\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4388_ _2443_ net589 _2446_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3339_ _1702_ _1742_ _1744_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _1472_ _1487_ _1488_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3069__A1 _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5009_ _2937_ _2939_ _2941_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_83_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output471_I net471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5384__I3 dffram.data\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3963__I _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3203__I _1641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3690_ _1849_ _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__I _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ dffram.data\[32\]\[2\] dffram.data\[34\]\[2\] dffram.data\[36\]\[2\] dffram.data\[38\]\[2\]
+ _0807_ _0808_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__4732__A1 net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4311_ _2387_ _2389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5291_ _0796_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4242_ dffram.data\[16\]\[0\] _2343_ _2344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_39_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4173_ _2298_ _2291_ _2299_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3124_ dffram.data\[8\]\[2\] _1597_ _1600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3055_ _1453_ _1544_ _1547_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3223__A1 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3957_ _2112_ _2152_ _2156_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _0596_ clknet_leaf_76_wb_clk_i dffram.data\[38\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _2111_ _2112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5627_ _1126_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_147_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input63_I mc14500_do[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5920__C2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5558_ _1057_ _1060_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4509_ _1493_ _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _0992_ _0993_ _0879_ _0994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_137_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__B _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3214__A1 _1659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4789__I _2776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4714__A1 net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4860_ wb_counter\[16\] _2830_ wb_counter\[17\] _2835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3205__A1 _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ dffram.data\[13\]\[6\] _2056_ _2059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4791_ _2593_ _2778_ _2779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6530_ _0450_ clknet_leaf_133_wb_clk_i net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3742_ _2011_ _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3673_ _1965_ _1967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _0381_ clknet_leaf_137_wb_clk_i dffram.data\[20\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5902__B1 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5412_ _0738_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_88_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6392_ _0312_ clknet_leaf_138_wb_clk_i dffram.data\[19\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5343_ _0692_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_58_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3108__I _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ dffram.data\[8\]\[0\] dffram.data\[10\]\[0\] dffram.data\[12\]\[0\] dffram.data\[14\]\[0\]
+ _0782_ _0783_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_103_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ _2286_ _2328_ _2332_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_71_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4156_ _2286_ _2281_ _2287_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_71_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3107_ _1585_ _1578_ _1586_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3692__A1 _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5969__B1 _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ _2223_ _2240_ _2243_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input215_I qcpu_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3038_ dffram.data\[37\]\[4\] _1535_ _1536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4383__B _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5984__A3 _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_77_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5736__A3 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _2524_ _2925_ _2928_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5292__S1 _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6659_ _0579_ clknet_leaf_86_wb_clk_i dffram.data\[40\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5434__S _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3018__I net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5121__A1 _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__I _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output434_I net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3435__A1 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A1 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput37 diceroll_do[5] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput15 ay8913_do[22] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 ay8913_do[7] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput59 mc14500_do[24] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput48 mc14500_do[14] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__C _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5143__I _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _1900_ _2117_ _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4466__A3 _2503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5961_ net172 _1249_ _1299_ net106 _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__3426__A1 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4912_ _2735_ _2874_ _2877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5892_ _1344_ _1346_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4843_ _2761_ _2821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_16_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5274__S1 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _2549_ _2762_ _2765_ _2514_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_160_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_95_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6513_ _0433_ clknet_leaf_93_wb_clk_i dffram.data\[44\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3725_ dffram.data\[54\]\[1\] _2000_ _2002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6444_ _0364_ clknet_leaf_53_wb_clk_i dffram.data\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5318__I _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3656_ dffram.data\[24\]\[3\] _1951_ _1955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3587_ dffram.data\[25\]\[3\] _1903_ _1910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6375_ _0295_ clknet_leaf_143_wb_clk_i dffram.data\[21\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5326_ dffram.data\[25\]\[1\] dffram.data\[27\]\[1\] dffram.data\[29\]\[1\] dffram.data\[31\]\[1\]
+ _0832_ _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input165_I qcpu_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_124_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5103__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ dffram.data\[24\]\[0\] dffram.data\[26\]\[0\] dffram.data\[28\]\[0\] dffram.data\[30\]\[0\]
+ _0762_ _0763_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xinput408 net646 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input332_I tholin_riscv_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ _2314_ _2322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input26_I ay8913_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5188_ dffram.data\[32\]\[0\] dffram.data\[34\]\[0\] dffram.data\[36\]\[0\] dffram.data\[38\]\[0\]
+ _0696_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3665__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ dffram.data\[20\]\[5\] _2274_ _2276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3417__A1 dffram.data\[34\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5429__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4917__A1 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__I _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5164__S _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5893__A2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4081__A1 _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5581__A1 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3510_ _1859_ _1860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4042__I _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ dffram.data\[27\]\[0\] _2522_ _2523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3441_ _1803_ _1811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6160_ _0080_ clknet_leaf_89_wb_clk_i dffram.data\[33\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3372_ _1714_ _1763_ _1765_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _0628_ _0632_ net521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_51_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6091_ _0011_ clknet_leaf_78_wb_clk_i dffram.data\[35\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_51_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ dffram.data\[38\]\[3\] _2960_ _2964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3647__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_108_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5944_ net56 _1233_ _1250_ net14 _1391_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__S1 _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ net363 _1098_ _1331_ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_146_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4826_ _2793_ _2628_ _2790_ _2807_ _2808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_32_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_117_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input282_I sn76489_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4757_ _2750_ _2751_ _2752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3708_ dffram.data\[12\]\[3\] _1987_ _1991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ net424 _2665_ _2672_ _2694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6427_ _0347_ clknet_leaf_31_wb_clk_i dffram.data\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ dffram.data\[11\]\[4\] _1944_ _1945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _0278_ clknet_leaf_142_wb_clk_i dffram.data\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5309_ dffram.data\[49\]\[1\] dffram.data\[51\]\[1\] dffram.data\[53\]\[1\] dffram.data\[55\]\[1\]
+ _0816_ _0817_ _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_80_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3886__A1 _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_145_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput205 qcpu_oeb[25] net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6289_ _0209_ clknet_leaf_49_wb_clk_i dffram.data\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput216 qcpu_oeb[5] net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput227 qcpu_sram_gwe net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_145_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_126_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput238 sid_do[11] net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput249 sid_do[2] net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_162_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_123_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4063__A1 _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3810__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_169_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__S1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold34_I wbs_dat_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5618__A2 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__S0 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold4 wbs_dat_i[14] net584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _2179_ _2180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5477__S1 _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ net190 _1144_ _1149_ net124 net326 _1146_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_84_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4611_ wb_counter\[8\] _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_44_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5591_ _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_81_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _2547_ _2566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4473_ net402 _2510_ _2511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6212_ _0132_ clknet_leaf_67_wb_clk_i dffram.data\[28\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5401__S1 _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3424_ _1784_ _1797_ _1800_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3868__A1 _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6143_ _0063_ clknet_leaf_22_wb_clk_i dffram.data\[63\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5532__S _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3355_ _1722_ _1748_ _1753_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3286_ _1702_ _1705_ _1707_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6074_ _1472_ _1501_ _1502_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5025_ dffram.data\[3\]\[5\] _2950_ _2953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input128_I pdp11_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4045__A1 _2169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5468__S1 _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ net53 _1315_ _1267_ net99 _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_101_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input93_I pdp11_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5858_ _1314_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5789_ net65 _1254_ _1255_ net111 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5396__I1 _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ wb_counter\[7\] _2793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_134_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3026__I _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold4_I wbs_dat_i[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output514_I net514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__S1 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5784__B2 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput509 net509 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5839__A2 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__I _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_152_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3140_ _1609_ _1610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3071_ _1556_ _1557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_161_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5775__A1 net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5712_ _1145_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3973_ dffram.data\[50\]\[3\] _2161_ _2168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6692_ _0612_ clknet_leaf_64_wb_clk_i dffram.data\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ _1109_ _1137_ net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_116_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5574_ _1075_ _1076_ _0736_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4525_ net370 _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4456_ _2495_ net633 _2491_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3407_ _1788_ _1781_ _1789_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4387_ _2434_ _2446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3338_ dffram.data\[30\]\[0\] _1743_ _1744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input245_I sid_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6126_ _0046_ clknet_leaf_10_wb_clk_i dffram.data\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3269_ _1649_ _1690_ _1695_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6057_ dffram.data\[36\]\[5\] _1480_ _1488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input412_I wbs_stb_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ dffram.data\[3\]\[0\] _2940_ _2941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4018__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5310__S0 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output464_I net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5236__I _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4257__A1 _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4009__A1 _2177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_41_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5347__S _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4310_ _2387_ _2388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5290_ _0794_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_77_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ _2341_ _2343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4985__I _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4496__A1 dffram.data\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4172_ dffram.data\[15\]\[7\] _2292_ _2299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3123_ _1568_ _1596_ _1599_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3054_ dffram.data\[43\]\[1\] _1545_ _1547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5540__S0 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4934__B _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3956_ dffram.data\[59\]\[6\] _2153_ _2156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6675_ _0595_ clknet_leaf_76_wb_clk_i dffram.data\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5626_ _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input195_I qcpu_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3887_ _1492_ _2111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5920__A1 net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__B2 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5056__I _2971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ dffram.data\[48\]\[7\] dffram.data\[50\]\[7\] dffram.data\[52\]\[7\] dffram.data\[54\]\[7\]
+ _1058_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_input362_I ue1_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5359__S0 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4508_ _2534_ _2531_ _2535_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5488_ dffram.data\[48\]\[5\] dffram.data\[50\]\[5\] dffram.data\[52\]\[5\] dffram.data\[54\]\[5\]
+ _0956_ _0957_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_input56_I mc14500_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4439_ net431 _2481_ _2484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4487__A1 _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4239__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6109_ _0029_ clknet_leaf_87_wb_clk_i dffram.data\[43\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5436__B1 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__S0 _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__A1 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4135__I _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__A2 _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3810_ _2041_ _2055_ _2058_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4790_ wb_counter\[0\] wb_counter\[1\] wb_counter\[2\] wb_counter\[3\] _2778_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_157_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _1423_ _0963_ _2011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6460_ _0380_ clknet_leaf_60_wb_clk_i dffram.data\[20\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3672_ _1965_ _1966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5902__A1 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__B2 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5411_ _0916_ _0917_ _0875_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6391_ _0311_ clknet_leaf_138_wb_clk_i dffram.data\[19\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5342_ dffram.data\[1\]\[1\] dffram.data\[3\]\[1\] dffram.data\[5\]\[1\] dffram.data\[7\]\[1\]
+ _0776_ _0778_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_58_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5273_ _0777_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4224_ dffram.data\[45\]\[2\] _2329_ _2332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4155_ dffram.data\[15\]\[2\] _2282_ _2287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3106_ dffram.data\[7\]\[6\] _1579_ _1586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5969__A1 net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4086_ dffram.data\[14\]\[1\] _2241_ _2243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input110_I pdp11_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3037_ _1527_ _1535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input208_I qcpu_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4988_ dffram.data\[40\]\[1\] _2926_ _2928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3939_ _2131_ _1638_ _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6658_ _0578_ clknet_leaf_85_wb_clk_i dffram.data\[40\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5609_ _0671_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_144_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_46_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _0509_ clknet_leaf_120_wb_clk_i net539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3380__A1 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output427_I net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5432__I0 dffram.data\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput27 ay8913_do[8] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput16 ay8913_do[23] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 diceroll_do[6] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_162_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput49 mc14500_do[15] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5648__B1 _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3123__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3879__I _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ net18 _1400_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__B1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5891_ net263 _1345_ _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _2412_ _2876_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4842_ _2802_ _2819_ _2820_ _2814_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5179__A2 _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4773_ net380 _2764_ _2765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3724_ _1962_ _1999_ _2001_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4503__I _2520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _0432_ clknet_leaf_103_wb_clk_i dffram.data\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3655_ _1907_ _1950_ _1954_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6443_ _0363_ clknet_leaf_50_wb_clk_i dffram.data\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3119__I _1595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__S _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3586_ _1841_ _1909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3362__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6374_ _0294_ clknet_leaf_143_wb_clk_i dffram.data\[21\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5325_ _0833_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_73_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5103__A2 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _0761_ _0764_ _0765_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput409 net647 net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input158_I qcpu_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4207_ _2314_ _2321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input325_I tholin_riscv_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5270__S _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _0682_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4862__A1 net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4138_ _2229_ _2273_ _2275_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input19_I ay8913_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4069_ _2219_ _2231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_88_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3353__A1 _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output544_I net544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5496__I3 dffram.data\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3408__A2 _1755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4081__A2 _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3440_ _1803_ _1810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3371_ dffram.data\[2\]\[4\] _1764_ _1765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5110_ _0631_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6090_ _0010_ clknet_leaf_78_wb_clk_i dffram.data\[35\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_51_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _2944_ _2959_ _2963_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5943_ _1389_ _1390_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5874_ _1274_ _1329_ _1330_ _1331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_103_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4825_ wb_counter\[9\] wb_counter\[10\] _2807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4756_ net437 _2629_ _2632_ _2751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ _1971_ _1986_ _1990_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ wb_counter\[19\] _2693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6426_ _0346_ clknet_leaf_31_wb_clk_i dffram.data\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3638_ _1936_ _1944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input275_I sn76489_do[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3335__A1 _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3569_ dffram.data\[10\]\[6\] _1894_ _1897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6357_ _0277_ clknet_leaf_143_wb_clk_i dffram.data\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _0726_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput206 qcpu_oeb[26] net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput217 qcpu_oeb[6] net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6288_ _0208_ clknet_leaf_11_wb_clk_i dffram.data\[56\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_145_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5239_ _0707_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput239 sid_do[12] net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput228 qcpu_sram_in[0] net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__B _1363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output494_I net494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5012__A1 _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__I _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__C1 net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__A1 _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__S1 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold5 net584 net582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_134_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5149__I _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5003__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _2619_ _2627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_44_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5590_ _0652_ _1091_ _1092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ net544 _2542_ _2565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ _2509_ _2510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6211_ _0131_ clknet_leaf_67_wb_clk_i dffram.data\[28\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3317__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3423_ dffram.data\[34\]\[5\] _1798_ _1800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6142_ _0062_ clknet_leaf_25_wb_clk_i dffram.data\[63\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3354_ dffram.data\[30\]\[7\] _1749_ _1753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__I _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3285_ dffram.data\[32\]\[0\] _1706_ _1707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6073_ dffram.data\[36\]\[7\] _1480_ _1502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4817__A1 net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5024_ _1486_ _2952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4228__I _2327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5242__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ net246 _1282_ _1260_ net268 net287 _0664_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_101_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ net259 _1222_ _1315_ net44 _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5788_ _1115_ _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input86_I mc14500_sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _2777_ _2791_ _2792_ _2786_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_161_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3556__A1 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4739_ _2619_ _2735_ _2736_ _2737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _0329_ clknet_leaf_64_wb_clk_i dffram.data\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output507_I net507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__I _2159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5784__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__I _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3070_ _1443_ _1556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__I _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5711_ _1162_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3972_ _2100_ _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3786__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6691_ _0611_ clknet_leaf_65_wb_clk_i dffram.data\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ net218 _1131_ _1135_ net152 net354 _1133_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_128_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5932__C1 net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3538__A1 _1839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5573_ dffram.data\[25\]\[7\] dffram.data\[27\]\[7\] dffram.data\[29\]\[7\] dffram.data\[31\]\[7\]
+ _0678_ _0683_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_41_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ wb_counter\[0\] _2549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ net401 _2489_ _2496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ dffram.data\[28\]\[7\] _1782_ _1789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4386_ net382 _2444_ _2445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3337_ _1741_ _1743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6125_ _0045_ clknet_leaf_12_wb_clk_i dffram.data\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input140_I pdp11_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input238_I sid_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3268_ dffram.data\[6\]\[3\] _1691_ _1695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6056_ _1486_ _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5007_ _2938_ _2940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3199_ dffram.data\[62\]\[3\] _1643_ _1650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5310__S1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5909_ net244 _1230_ _1287_ net266 net288 _0664_ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_76_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3529__A1 _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3037__I _1527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__S _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output457_I net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__A1 net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3500__I _1492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold94_I wbs_dat_i[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4193__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4331__I net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4240_ _2341_ _2342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4171_ _2114_ _2298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3122_ dffram.data\[8\]\[1\] _1597_ _1599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3053_ _1445_ _1544_ _1546_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5996__A2 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5540__S1 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3410__I _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3955_ _2109_ _2152_ _2155_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3759__A1 _1979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _0594_ clknet_leaf_76_wb_clk_i dffram.data\[38\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _1104_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3886_ _2109_ _2105_ _2110_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_152_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4241__I _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5337__I _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input188_I qcpu_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5556_ _0743_ _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__S1 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5487_ dffram.data\[56\]\[5\] dffram.data\[58\]\[5\] dffram.data\[60\]\[5\] dffram.data\[62\]\[5\]
+ _0919_ _0920_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4507_ dffram.data\[27\]\[5\] _2532_ _2535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input355_I tholin_riscv_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4438_ _2482_ _2483_ _2480_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input49_I mc14500_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4369_ _2431_ _2432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6108_ _0028_ clknet_leaf_79_wb_clk_i dffram.data\[43\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5800__I _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6039_ _1436_ _1470_ _1471_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__S1 _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3990__I _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__A1 _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5978__A2 _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3989__A1 _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3740_ _1983_ _2005_ _2010_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3671_ _1724_ _1964_ _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_24_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5410_ dffram.data\[57\]\[3\] dffram.data\[59\]\[3\] dffram.data\[61\]\[3\] dffram.data\[63\]\[3\]
+ _0872_ _0873_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_11_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6390_ _0310_ clknet_leaf_138_wb_clk_i dffram.data\[19\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5341_ dffram.data\[9\]\[1\] dffram.data\[11\]\[1\] dffram.data\[13\]\[1\] dffram.data\[15\]\[1\]
+ _0848_ _0849_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_58_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5272_ _0781_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_128_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _2284_ _2328_ _2331_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4154_ _2097_ _2286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_71_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4085_ _2218_ _2240_ _2242_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3105_ _1584_ _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5969__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3036_ _1527_ _1534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A2 wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3140__I _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input103_I pdp11_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_154_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4987_ _2519_ _2925_ _2927_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3938_ _2115_ _2139_ _2144_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_150_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3869_ _1459_ _2097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_78_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6657_ _0577_ clknet_leaf_111_wb_clk_i dffram.data\[41\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _0663_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6588_ _0508_ clknet_leaf_120_wb_clk_i net538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3904__A1 _2098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5539_ _0707_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3315__I _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3050__I _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4590__B _2608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4396__A1 net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput17 ay8913_do[24] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 ay8913_do[9] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 diceroll_do[7] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A1 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__B2 net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold57_I wbs_dat_i[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5648__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5648__B2 _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__B2 net319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5820__A1 net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _1221_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4910_ net398 _2800_ _2875_ _2876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4841_ net384 _2804_ _2820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__I _1963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4772_ _2763_ _2764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_95_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3723_ dffram.data\[54\]\[0\] _2000_ _2001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6511_ _0431_ clknet_leaf_104_wb_clk_i dffram.data\[18\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3654_ dffram.data\[24\]\[2\] _1951_ _1954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6442_ _0362_ clknet_leaf_53_wb_clk_i dffram.data\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5887__B2 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5887__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5615__I _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3585_ _1907_ _1902_ _1908_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6373_ _0293_ clknet_leaf_143_wb_clk_i dffram.data\[21\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5324_ _0681_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5255_ _0735_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5551__S _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4206_ _2288_ _2315_ _2320_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_147_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5186_ _0677_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_108_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input220_I qcpu_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ dffram.data\[20\]\[4\] _2274_ _2275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input318_I tholin_riscv_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _2219_ _2230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5811__B2 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5811__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3019_ _1521_ _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_133_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A1 net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput490 net490 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_128_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4302__A1 _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmultiplexer_570 irq[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5802__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__I1 dffram.data\[34\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3041__A1 _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5169__I0 net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3370_ _1756_ _1764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A1 net544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ dffram.data\[38\]\[2\] _2960_ _2963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4844__A2 wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5942_ net290 _0662_ _1177_ net102 _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5873_ net46 _1232_ _1105_ net294 _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_103_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4824_ wb_counter\[9\] _2797_ wb_counter\[10\] _2806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4755_ _2548_ wb_counter\[30\] _2750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3706_ dffram.data\[12\]\[2\] _1987_ _1990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_146_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5404__S0 _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4686_ _2669_ _2692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _0345_ clknet_leaf_31_wb_clk_i dffram.data\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3637_ _1936_ _1943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input170_I qcpu_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _0276_ clknet_leaf_55_wb_clk_i dffram.data\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3568_ _1850_ _1893_ _1896_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input268_I sn76489_do[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _0723_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_45_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput207 qcpu_oeb[27] net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput218 qcpu_oeb[7] net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3499_ _1850_ _1846_ _1851_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6287_ _0207_ clknet_leaf_11_wb_clk_i dffram.data\[56\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input31_I blinker_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5238_ _0741_ _0745_ _0747_ _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3099__A1 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput229 qcpu_sram_in[1] net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ net375 net76 _0673_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_123_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output487_I net487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_169_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_169_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_30_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5255__I _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold6 _2453_ net583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4826__A2 _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4540_ _2543_ _2564_ _2501_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__A1 net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _2507_ _2508_ _2403_ _2509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_150_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6210_ _0130_ clknet_leaf_68_wb_clk_i dffram.data\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3422_ _1780_ _1797_ _1799_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4514__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _0061_ clknet_leaf_24_wb_clk_i dffram.data\[63\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3353_ _1720_ _1748_ _1752_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3284_ _1704_ _1706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__I0 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6072_ _1500_ _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5023_ _2948_ _2949_ _2951_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_85_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5925_ _1246_ _1371_ _1375_ net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_101_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _1205_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_81_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4807_ net409 _2781_ _2792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ _1205_ _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3005__A1 _1461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2999_ _1508_ _1510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ net433 _2615_ _2710_ _2736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_39_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input79_I mc14500_sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4669_ _2653_ wb_counter\[16\] _2678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4505__A1 _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _0328_ clknet_leaf_7_wb_clk_i dffram.data\[50\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5803__I _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _0259_ clknet_leaf_27_wb_clk_i dffram.data\[53\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_48_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3244__A1 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3971_ _2165_ _2160_ _2166_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3235__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ _1188_ _1189_ net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_63_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _0610_ clknet_leaf_64_wb_clk_i dffram.data\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_75_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _1109_ _1136_ net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ dffram.data\[17\]\[7\] dffram.data\[19\]\[7\] dffram.data\[21\]\[7\] dffram.data\[23\]\[7\]
+ _0762_ _0763_ _1075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_81_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _2547_ _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5696__C1 net334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4454_ net435 _2492_ _2495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5160__A1 _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3405_ _1587_ _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4385_ _2431_ _2444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3336_ _1741_ _1742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6124_ _0044_ clknet_leaf_41_wb_clk_i dffram.data\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_84_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6055_ _1485_ _1486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input133_I pdp11_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _2938_ _2939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3267_ _1647_ _1690_ _1694_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3198_ _1573_ _1649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input300_I tholin_riscv_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_93_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5908_ _1245_ _1355_ _1356_ _1360_ net490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5839_ net72 _1264_ _1299_ net120 _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_146_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold87_I wbs_dat_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3228__I _1663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__I0 _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5142__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A2 _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _2296_ _2291_ _2297_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3121_ _1557_ _1596_ _1598_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3456__A1 _1774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3052_ dffram.data\[43\]\[0\] _1545_ _1546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3898__I _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput390 net585 net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3208__A1 _1655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3954_ dffram.data\[59\]\[5\] _2153_ _2155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6673_ _0593_ clknet_leaf_57_wb_clk_i dffram.data\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3885_ dffram.data\[21\]\[5\] _2106_ _2110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5624_ _1123_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__A1 net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5555_ _0826_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_113_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5486_ _0989_ _0990_ _0875_ _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4506_ _1486_ _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5133__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4437_ net396 _2478_ _2483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input348_I tholin_riscv_oeb[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input250_I sid_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__I3 dffram.data\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6107_ _0027_ clknet_leaf_80_wb_clk_i dffram.data\[43\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3695__A1 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4368_ _2430_ _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3319_ _1708_ _1728_ _1731_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4299_ _2374_ _2381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6038_ dffram.data\[36\]\[3\] _1446_ _1471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3447__A1 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4947__A1 _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4175__A2 _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5464__S _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4588__B _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3511__I _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_169_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3610__A1 _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3670_ _1963_ _1964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5340_ _0682_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_58_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5271_ _0722_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4222_ dffram.data\[45\]\[1\] _2329_ _2331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4153_ _2284_ _2281_ _2285_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4084_ dffram.data\[14\]\[0\] _2241_ _2242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3429__A1 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3104_ _1492_ _1584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3035_ _1470_ _1528_ _1533_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4986_ dffram.data\[40\]\[0\] _2926_ _2927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3937_ dffram.data\[19\]\[7\] _2140_ _2144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input298_I tholin_riscv_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3868_ _2095_ _2091_ _2096_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_78_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6656_ _0576_ clknet_leaf_111_wb_clk_i dffram.data\[41\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5607_ _0652_ _1089_ _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_132_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3799_ dffram.data\[13\]\[1\] _2050_ _2052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _0507_ clknet_leaf_120_wb_clk_i net537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1026_ _1041_ net518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_input61_I mc14500_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5469_ _0723_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_126_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4162__I _2280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 ay8913_do[25] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput29 blinker_do[0] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_150_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3831__A1 _2041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ wb_counter\[13\] _2818_ _2819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_158_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_99_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__I _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4771_ _2759_ _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_136_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6510_ _0430_ clknet_leaf_104_wb_clk_i dffram.data\[18\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3722_ _1998_ _2000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3653_ _1905_ _1950_ _1953_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _0361_ clknet_leaf_52_wb_clk_i dffram.data\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _0292_ clknet_leaf_55_wb_clk_i dffram.data\[21\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3584_ dffram.data\[25\]\[2\] _1903_ _1908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5323_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_110_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5254_ dffram.data\[25\]\[0\] dffram.data\[27\]\[0\] dffram.data\[29\]\[0\] dffram.data\[31\]\[0\]
+ _0762_ _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4205_ dffram.data\[1\]\[3\] _2316_ _2320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5185_ dffram.data\[40\]\[0\] dffram.data\[42\]\[0\] dffram.data\[44\]\[0\] dffram.data\[46\]\[0\]
+ _0678_ _0683_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_147_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4136_ _2266_ _2274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input213_I qcpu_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3151__I _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4067_ _2103_ _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5811__A2 _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3822__A1 dffram.data\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3018_ net368 _1521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__S _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4969_ dffram.data\[41\]\[2\] _2913_ _2916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6639_ _0559_ clknet_4_8_0_wb_clk_i wb_override_act vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_104_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput480 net480 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_167_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput491 net491 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_128_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output432_I net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__A1 _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3061__I _1543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmultiplexer_571 irq[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_158_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5189__S _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5169__I1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5451__I _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4057__A1 _2218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5941_ net271 _1345_ _1102_ net168 _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_88_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3804__A1 _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ net239 _1269_ _1329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_103_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _2802_ _2803_ _2805_ _2786_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4754_ _2734_ _2749_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3705_ _1969_ _1986_ _1989_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5404__S1 _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ _2670_ _2691_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4530__I net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3636_ _1909_ _1937_ _1942_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _0344_ clknet_leaf_5_wb_clk_i dffram.data\[49\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6355_ _0275_ clknet_leaf_50_wb_clk_i dffram.data\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3567_ dffram.data\[10\]\[5\] _1894_ _1896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5306_ _0803_ _0812_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6286_ _0206_ clknet_leaf_11_wb_clk_i dffram.data\[56\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input163_I qcpu_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput208 qcpu_oeb[28] net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3498_ dffram.data\[58\]\[5\] _1847_ _1851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5237_ _0746_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input330_I tholin_riscv_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput219 qcpu_oeb[8] net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input24_I ay8913_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5168_ _0677_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4119_ dffram.data\[47\]\[6\] _2260_ _2263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5099_ design_select\[1\] design_select\[4\] _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3023__A2 _1505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_104_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5720__B2 net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__A1 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5472__S _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5271__I _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold7 wbs_dat_i[15] net587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4039__A1 _2165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_18_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5331__S0 _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_122_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4470_ net413 _2508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3421_ dffram.data\[34\]\[4\] _1798_ _1799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6140_ _0060_ clknet_leaf_33_wb_clk_i dffram.data\[63\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3352_ dffram.data\[30\]\[6\] _1749_ _1752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3283_ _1704_ _1705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5475__B1 _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6071_ _1499_ _1500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5022_ dffram.data\[3\]\[4\] _2950_ _2951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5924_ net245 _1230_ _1103_ net164 _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4525__I net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5855_ net156 _1114_ _1267_ net90 _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ wb_counter\[7\] _2790_ _2791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5786_ net278 _1222_ _1252_ net33 _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4202__A1 _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ _1508_ _1509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input280_I sn76489_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ wb_counter\[27\] _2735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input378_I wbs_adr_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4668_ _2625_ _2677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3619_ dffram.data\[56\]\[5\] _1930_ _1932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6407_ _0327_ clknet_leaf_8_wb_clk_i dffram.data\[50\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4599_ _2553_ _2617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_164_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6338_ _0258_ clknet_leaf_26_wb_clk_i dffram.data\[53\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _0189_ clknet_leaf_10_wb_clk_i dffram.data\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5769__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__I _2408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__S _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5941__B2 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5941__A1 net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__I _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3180__A1 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5552__S0 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ dffram.data\[50\]\[2\] _2161_ _2166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4432__A1 net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__A2 _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ net217 _1131_ _1135_ net151 net353 _1133_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_130_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5932__B2 net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5932__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _1042_ _1068_ _1073_ _0719_ _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5176__I _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4522_ _2546_ _2547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ _2493_ net639 _2491_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A1 dffram.data\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3404_ _1786_ _1781_ _1787_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5160__A2 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4384_ net416 _2436_ _2443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6123_ _0043_ clknet_leaf_51_wb_clk_i dffram.data\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3335_ _1740_ _1726_ _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ dffram.data\[6\]\[2\] _1691_ _1694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6054_ net233 _1473_ _1484_ _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5005_ _2131_ _1559_ _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5543__S0 _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3197_ _1647_ _1642_ _1648_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input126_I pdp11_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4255__I _2341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ net243 _1215_ _1357_ net298 _1359_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_113_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input91_I pdp11_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _1155_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_10_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5769_ net41 _0653_ _0655_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__I _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5526__I1 dffram.data\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3162__A1 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output512_I net512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3217__A2 _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__A1 net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3153__A1 _1577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ dffram.data\[8\]\[0\] _1597_ _1598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3051_ _1543_ _1545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput380 net651 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput391 net653 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4405__A1 net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3953_ _2104_ _2152_ _2154_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ _0592_ clknet_leaf_58_wb_clk_i dffram.data\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3884_ _2108_ _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5623_ _1095_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5905__A1 net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3419__I _1790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5554_ _0734_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5485_ dffram.data\[57\]\[5\] dffram.data\[59\]\[5\] dffram.data\[61\]\[5\] dffram.data\[63\]\[5\]
+ _0872_ _0873_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4505_ _2530_ _2531_ _2533_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4436_ net430 _2481_ _2482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4367_ net370 _2401_ _2404_ _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3318_ dffram.data\[31\]\[1\] _1729_ _1731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6106_ _0026_ clknet_leaf_80_wb_clk_i dffram.data\[43\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input243_I sid_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_127_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4298_ _2349_ _2375_ _2380_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5516__S0 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _1469_ _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3249_ _1676_ _1683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__B1 _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output462_I net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5124__A2 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3135__A1 _1585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5832__B1 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5060__A1 _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3239__I _1676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3374__A1 _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5270_ _0775_ _0779_ _0693_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3126__A1 dffram.data\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _2279_ _2328_ _2330_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4152_ dffram.data\[15\]\[1\] _2282_ _2285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4083_ _2239_ _2241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3103_ _1582_ _1578_ _1583_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5823__B1 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3034_ dffram.data\[37\]\[3\] _1529_ _1533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4626__A1 _2621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4985_ _2924_ _2926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5051__A1 _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _2112_ _2139_ _2143_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input193_I qcpu_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3867_ dffram.data\[21\]\[1\] _2092_ _2096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5565__S _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ _0575_ clknet_leaf_112_wb_clk_i dffram.data\[41\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ _1089_ _1093_ _1099_ _1107_ net474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_116_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3798_ _2026_ _2049_ _2051_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6586_ _0506_ clknet_leaf_120_wb_clk_i net536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5364__I _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5537_ _0963_ _1033_ _1040_ _0980_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA_input360_I ue1_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input54_I mc14500_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3117__A1 _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ dffram.data\[8\]\[4\] dffram.data\[10\]\[4\] dffram.data\[12\]\[4\] dffram.data\[14\]\[4\]
+ _0937_ _0938_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5399_ _0774_ _0895_ _0906_ _0792_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_79_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4865__A1 net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4419_ _2465_ net586 _2469_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__I _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 ay8913_do[26] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__A1 net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5281__A1 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4353__I _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4770_ _2761_ _2762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3721_ _1998_ _1999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3652_ dffram.data\[24\]\[1\] _1951_ _1953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6440_ _0360_ clknet_leaf_9_wb_clk_i dffram.data\[48\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3583_ _1838_ _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6371_ _0291_ clknet_leaf_55_wb_clk_i dffram.data\[21\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5322_ _0676_ _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _0682_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4847__A1 net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4204_ _2286_ _2315_ _2319_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5184_ _0684_ _0685_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_147_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4528__I _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4135_ _2266_ _2273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4066_ _2227_ _2220_ _2228_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3017_ _1501_ _1515_ _1520_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input206_I qcpu_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_159_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ _2524_ _2912_ _2915_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5980__C1 net314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3919_ _2132_ _2133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4899_ net396 _2866_ _2867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6638_ _0558_ clknet_leaf_135_wb_clk_i wb_counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__B1 _2554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _0489_ clknet_leaf_73_wb_clk_i dffram.data\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_142_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_142_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_168_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_167_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5822__I _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput470 net470 io_oeb[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput492 net492 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput481 net481 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_128_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output425_I net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__A1 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmultiplexer_572 irq[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_97_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5015__A1 _2944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_13_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3329__A1 _1718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4829__A1 net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5940_ net304 _1152_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_158_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5871_ net261 _1287_ _1156_ net92 _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_146_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4083__I _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ net411 _2804_ _2805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5962__C1 net308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3568__A1 _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4753_ net554 _2739_ _2740_ _2748_ _2749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_160_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3704_ dffram.data\[12\]\[1\] _1987_ _1989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6423_ _0343_ clknet_leaf_7_wb_clk_i dffram.data\[49\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ net542 _2676_ _2677_ _2690_ _2691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_144_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ dffram.data\[11\]\[3\] _1938_ _1942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ _0274_ clknet_leaf_54_wb_clk_i dffram.data\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3566_ _1845_ _1893_ _1895_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_149_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5305_ _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6285_ _0205_ clknet_leaf_11_wb_clk_i dffram.data\[56\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3497_ _1849_ _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3740__A1 _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput209 qcpu_oeb[29] net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5236_ _0691_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input156_I qcpu_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_162_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input323_I tholin_riscv_do[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5167_ _0676_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5098_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_98_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4118_ _2233_ _2259_ _2262_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input17_I ay8913_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4049_ _2175_ _2212_ _2216_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_140_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__A2 _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__C1 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_169_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3337__I _1741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__B _2796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold8 net605 net585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_89_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5331__S1 _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3798__A1 _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4631__I _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3420_ _1790_ _1798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3351_ _1718_ _1748_ _1751_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I ay8913_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3282_ _1703_ _1594_ _1704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6070_ net235 _1473_ _1498_ _1499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_29_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5021_ _2938_ _2950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3789__A1 _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3710__I _1985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5923_ _1344_ _1372_ _1373_ _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5854_ net237 _1230_ _1312_ net2 net292 _1106_ _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_150_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4805_ wb_counter\[4\] wb_counter\[5\] wb_counter\[6\] _2778_ _2790_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_146_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5785_ _1090_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2997_ _1425_ _1507_ _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4736_ _2669_ _2734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3961__A1 _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4667_ _2582_ _2676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3618_ _1911_ _1929_ _1931_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6406_ _0326_ clknet_leaf_8_wb_clk_i dffram.data\[50\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input273_I sn76489_do[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6337_ _0257_ clknet_leaf_27_wb_clk_i dffram.data\[53\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4598_ _2615_ _2616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3713__A1 _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3549_ dffram.data\[57\]\[7\] _1880_ _1884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6268_ _0188_ clknet_leaf_39_wb_clk_i dffram.data\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _0119_ clknet_leaf_96_wb_clk_i dffram.data\[30\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5219_ _0723_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5769__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output492_I net492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__C1 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold25_I wbs_dat_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__S1 _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_100_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4196__A1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _1070_ _1072_ _1062_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__A1 _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ net371 _2546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ net400 _2489_ _2494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5696__B2 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A1 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3403_ dffram.data\[28\]\[6\] _1782_ _1787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4383_ _2441_ net619 _2435_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6122_ _0042_ clknet_leaf_40_wb_clk_i dffram.data\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3334_ _1639_ _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3265_ _1645_ _1690_ _1693_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6053_ _1482_ _1464_ _1483_ _1457_ _1484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_147_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5004_ _1444_ _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5999__A2 _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__S1 _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4120__A1 _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3196_ dffram.data\[62\]\[2\] _1643_ _1648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3440__I _1803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input119_I pdp11_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5906_ _1344_ _1358_ _1359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5620__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5837_ _1293_ _1294_ _1298_ net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_147_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5367__I _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5768_ _1110_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_134_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input84_I mc14500_sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4719_ _2624_ _2720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3934__A1 _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _1172_ _1180_ net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_135_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__S0 _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3615__I _1922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output505_I net505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__I _2430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5611__A1 net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5222__S0 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3050_ _1543_ _1544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A1 net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput381 net618 net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput370 net642 net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__B2 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3260__I _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput392 net591 net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5289__S0 _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5453__I1 _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3952_ dffram.data\[59\]\[4\] _2153_ _2154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _0591_ clknet_leaf_58_wb_clk_i dffram.data\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3883_ _1485_ _2108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ _1121_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5553_ _0802_ _1055_ _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5461__S0 _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3916__A1 _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4504_ dffram.data\[27\]\[4\] _2532_ _2533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5484_ dffram.data\[49\]\[5\] dffram.data\[51\]\[5\] dffram.data\[53\]\[5\] dffram.data\[55\]\[5\]
+ _0729_ _0731_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_158_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4435_ _2408_ _2481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_130_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4366_ net443 _2423_ _2429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3317_ _1702_ _1728_ _1730_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6105_ _0025_ clknet_leaf_80_wb_clk_i dffram.data\[43\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4297_ dffram.data\[44\]\[3\] _2376_ _2380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5516__S1 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input236_I sid_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3248_ _1649_ _1677_ _1682_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6036_ _1468_ _1469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5841__A1 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5841__B2 net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3179_ dffram.data\[63\]\[6\] _1632_ _1635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5097__I _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5452__S0 _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output455_I net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5832__A1 net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__I _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4399__A1 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold92_I wbs_dat_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4938__A3 _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5443__S0 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4220_ dffram.data\[45\]\[0\] _2329_ _2330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4323__A1 _2351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4151_ _2094_ _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5470__I _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ _2239_ _2240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3102_ dffram.data\[7\]\[5\] _1579_ _1583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__B2 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A1 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3033_ _1461_ _1528_ _1532_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4984_ _2924_ _2925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_154_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3935_ dffram.data\[19\]\[6\] _2140_ _2143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _0574_ clknet_leaf_111_wb_clk_i dffram.data\[41\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ net188 _1103_ _1106_ net324 _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_116_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3866_ _2094_ _2095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3797_ dffram.data\[13\]\[0\] _2050_ _2051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6585_ _0505_ clknet_leaf_121_wb_clk_i net535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5536_ _1036_ _1039_ _0749_ _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4562__A1 net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input186_I qcpu_do[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5467_ _0971_ _0972_ _0852_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input353_I tholin_riscv_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3117__A2 _1594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _2468_ _2469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input47_I mc14500_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5398_ _0900_ _0904_ _0905_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4865__A2 _2763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ net439 _2416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6019_ dffram.data\[36\]\[1\] _1446_ _1454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4617__A2 _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5555__I _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3356__A2 _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5281__A2 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3292__A1 _1710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _1740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_16_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _1740_ _1964_ _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _1899_ _1950_ _1952_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3582_ _1905_ _1902_ _1906_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6370_ _0290_ clknet_leaf_55_wb_clk_i dffram.data\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5321_ dffram.data\[17\]\[1\] dffram.data\[19\]\[1\] dffram.data\[21\]\[1\] dffram.data\[23\]\[1\]
+ _0827_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_139_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5252_ _0757_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4203_ dffram.data\[1\]\[2\] _2316_ _2319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5183_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_147_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4134_ _2227_ _2267_ _2272_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4065_ dffram.data\[48\]\[3\] _2221_ _2228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3016_ dffram.data\[35\]\[7\] _1516_ _1520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__I _2552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input101_I pdp11_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3035__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4967_ dffram.data\[41\]\[1\] _2913_ _2915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5980__B1 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ _2131_ _2012_ _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_62_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4898_ _2760_ _2866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2999__I _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__I _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3849_ _2075_ _2083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6637_ _0557_ clknet_leaf_135_wb_clk_i wb_counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6568_ _0488_ clknet_leaf_73_wb_clk_i dffram.data\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__A1 _2548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5519_ dffram.data\[48\]\[6\] dffram.data\[50\]\[6\] dffram.data\[52\]\[6\] dffram.data\[54\]\[6\]
+ _0956_ _0957_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6499_ _0419_ clknet_leaf_73_wb_clk_i dffram.data\[16\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_167_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput471 net471 io_oeb[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput460 net460 io_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput493 net493 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput482 net482 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_121_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4719__I _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5799__B1 _1181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5263__A2 _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output418_I net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmultiplexer_573 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_167_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5994__B _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_94_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__I _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4526__A1 _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3265__A1 _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5870_ net158 _1325_ _1326_ net4 _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_76_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4821_ _2780_ _2804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5396__S _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3017__A1 _1501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4752_ _2746_ _2747_ _2748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4765__A1 _2754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3703_ _1962_ _1986_ _1988_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4683_ _2687_ _2689_ _2690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3634_ _1907_ _1937_ _1941_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6422_ _0342_ clknet_leaf_5_wb_clk_i dffram.data\[49\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _0273_ clknet_leaf_49_wb_clk_i dffram.data\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3565_ dffram.data\[10\]\[4\] _1894_ _1895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5190__A1 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6284_ _0204_ clknet_leaf_41_wb_clk_i dffram.data\[56\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5304_ _0706_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3496_ _1485_ _1849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5235_ dffram.data\[48\]\[0\] dffram.data\[50\]\[0\] dffram.data\[52\]\[0\] dffram.data\[54\]\[0\]
+ _0742_ _0744_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input149_I pdp11_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5166_ _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5097_ _0618_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4117_ dffram.data\[47\]\[5\] _2260_ _2262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input316_I tholin_riscv_do[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3256__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ dffram.data\[4\]\[6\] _2213_ _2216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5999_ _1425_ _1434_ _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_52_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4756__A1 net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4508__A1 _2534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_18_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3495__A1 _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold9 _2467_ net586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_96_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_27_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3350_ dffram.data\[30\]\[5\] _1749_ _1751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5020_ _2938_ _2949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3281_ _1424_ _1703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_144_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3238__A1 _1526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5632__C1 net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5922_ net10 _1224_ _1117_ net300 _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_152_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5853_ _1224_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_119_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5784_ net177 _1249_ _1250_ net21 _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_4804_ _2777_ _2788_ _2789_ _2786_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4738__A1 net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _2714_ _2733_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4666_ _2670_ _2675_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3617_ dffram.data\[56\]\[4\] _1930_ _1931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6405_ _0325_ clknet_leaf_7_wb_clk_i dffram.data\[50\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4597_ _2614_ _2615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3548_ _1853_ _1879_ _1883_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input266_I sn76489_do[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4910__A1 net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ _0256_ clknet_leaf_144_wb_clk_i dffram.data\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4269__I _2361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3479_ _1835_ _1836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6267_ _0187_ clknet_leaf_39_wb_clk_i dffram.data\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3173__I _1624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3477__A1 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ dffram.data\[49\]\[0\] dffram.data\[51\]\[0\] dffram.data\[53\]\[0\] dffram.data\[55\]\[0\]
+ _0724_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6198_ _0118_ clknet_leaf_100_wb_clk_i dffram.data\[30\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5149_ _0663_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_4_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5769__A3 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output485_I net485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3401__A1 _1784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3468__A1 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_145_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__A2 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_35_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3640__A1 _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4196__A2 _1662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _2544_ _2545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_44_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ net434 _2492_ _2493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3402_ _1584_ _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5160__A4 _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6121_ _0041_ clknet_leaf_51_wb_clk_i dffram.data\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4382_ net381 _2432_ _2442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3333_ _1722_ _1734_ _1739_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3264_ dffram.data\[6\]\[1\] _1691_ _1693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6052_ net407 _1465_ _1483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_42_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5003_ _2538_ _2931_ _2936_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3195_ _1570_ _1647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3721__I _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4959__A1 _2536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ net265 _1345_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5620__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5836_ net358 _1236_ _1239_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_57_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5767_ net54 _1233_ _1234_ net302 _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_118_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5698_ net200 _1174_ _1178_ net134 net336 _1175_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_118_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4718_ _2544_ _2719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_135_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input77_I mc14500_sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4649_ net418 _2655_ _2660_ _2661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5687__A2 _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__S1 _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_9_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3698__A1 _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _0239_ clknet_leaf_9_wb_clk_i dffram.data\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_18_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_71_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3622__A1 _1917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3078__I _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__S _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5222__S1 _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3806__I _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3689__A1 _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4102__A2 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput360 ue1_do[3] net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3541__I _1872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput371 net623 net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput393 net597 net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput382 net588 net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5289__S1 _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3951_ _2145_ _2153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _0590_ clknet_leaf_56_wb_clk_i dffram.data\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _2104_ _2105_ _2107_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1113_ _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ dffram.data\[56\]\[7\] dffram.data\[58\]\[7\] dffram.data\[60\]\[7\] dffram.data\[62\]\[7\]
+ _0883_ _0828_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__5461__S1 _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _2520_ _2532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5669__A2 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5483_ _0984_ _0987_ _0914_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5508__I3 dffram.data\[47\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4434_ _2477_ _2479_ _2480_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_130_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4365_ _2427_ _2423_ _2428_ _2420_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3316_ dffram.data\[31\]\[0\] _1729_ _1730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6104_ _0024_ clknet_leaf_88_wb_clk_i dffram.data\[37\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4296_ _2347_ _2375_ _2379_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6035_ net231 _1438_ _1467_ _1468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA_input131_I pdp11_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3451__I _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3247_ dffram.data\[61\]\[3\] _1678_ _1682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3178_ _1582_ _1631_ _1634_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input229_I qcpu_sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_136_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5819_ net252 _1282_ _1233_ net69 _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_88_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__S1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output448_I net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3843__A1 _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__S _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5288__I _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold85_I wbs_adr_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5443__S1 _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__A1 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_58_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4150_ _2279_ _2281_ _2283_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3101_ _1581_ _1582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4087__A1 _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _1591_ _1640_ _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__3271__I _1689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3032_ dffram.data\[37\]\[2\] _1529_ _1532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput190 qcpu_oeb[11] net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5587__A1 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__I _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _2300_ _1594_ _2924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_53_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3934_ _2109_ _2139_ _2142_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3865_ _1451_ _2094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6653_ _0573_ clknet_leaf_85_wb_clk_i dffram.data\[41\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5604_ _1105_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3796_ _2048_ _2050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6584_ _0504_ clknet_leaf_123_wb_clk_i net534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5535_ _1037_ _1038_ _0747_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5466_ dffram.data\[1\]\[4\] dffram.data\[3\]\[4\] dffram.data\[5\]\[4\] dffram.data\[7\]\[4\]
+ _0897_ _0898_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input179_I qcpu_do[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4417_ _2418_ _2468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input346_I tholin_riscv_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _0707_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4348_ _1140_ _2407_ _2415_ _2412_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4279_ _2361_ _2369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6018_ _1452_ _1453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3825__A1 _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_92_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6058__A2 _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4187__I _2301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5746__I _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3650_ dffram.data\[24\]\[0\] _1951_ _1952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ dffram.data\[25\]\[1\] _1903_ _1906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_77_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer1 _0621_ net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_144_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5320_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_110_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5251_ dffram.data\[17\]\[0\] dffram.data\[19\]\[0\] dffram.data\[21\]\[0\] dffram.data\[23\]\[0\]
+ _0758_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_51_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ _2284_ _2315_ _2318_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5182_ _0691_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_147_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4133_ dffram.data\[20\]\[3\] _2268_ _2272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _2100_ _2227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_108_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3015_ _1494_ _1515_ _1519_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__A1 _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4966_ _2519_ _2912_ _2914_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5980__B2 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3917_ _1506_ _2131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4897_ wb_counter\[24\] _2859_ _2865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input296_I tholin_riscv_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _2075_ _2082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6636_ _0556_ clknet_leaf_105_wb_clk_i wb_counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6567_ _0487_ clknet_leaf_73_wb_clk_i dffram.data\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3779_ _1844_ _2037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_104_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5518_ dffram.data\[56\]\[6\] dffram.data\[58\]\[6\] dffram.data\[60\]\[6\] dffram.data\[62\]\[6\]
+ _0919_ _0920_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6498_ _0418_ clknet_leaf_93_wb_clk_i dffram.data\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_167_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5449_ dffram.data\[56\]\[4\] dffram.data\[58\]\[4\] dffram.data\[60\]\[4\] dffram.data\[62\]\[4\]
+ _0919_ _0920_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput450 net450 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput461 net461 io_oeb[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput494 net494 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput483 net483 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_121_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput472 net472 io_oeb[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__A1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__B2 net317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmultiplexer_574 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_167_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__C _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4223__A1 _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__I net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3086__I _1459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5574__I1 _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4526__A2 net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5334__S0 _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ wb_counter\[9\] _2797_ _2803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_111_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4214__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5962__B2 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5962__A1 net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ net435 _2629_ _2726_ _2747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3702_ dffram.data\[12\]\[0\] _1987_ _1988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4682_ net423 _2688_ _2660_ _2689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ dffram.data\[11\]\[2\] _1938_ _1941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6421_ _0341_ clknet_leaf_4_wb_clk_i dffram.data\[49\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3564_ _1886_ _1894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6352_ _0272_ clknet_leaf_140_wb_clk_i dffram.data\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5190__A2 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6283_ _0203_ clknet_leaf_45_wb_clk_i dffram.data\[56\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5303_ _0806_ _0809_ _0811_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3495_ _1845_ _1846_ _1848_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _0743_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5573__S0 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ net222 _0674_ _0646_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4116_ _2229_ _2259_ _2261_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_162_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5096_ design_select\[0\] _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_123_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4047_ _2173_ _2212_ _2215_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input309_I tholin_riscv_do[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input211_I qcpu_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _1433_ _1434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_52_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__A1 net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5953__B2 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _2526_ _2899_ _2903_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__I _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6619_ _0539_ clknet_leaf_129_wb_clk_i wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__A2 _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__I _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5564__S0 _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output430_I net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output528_I net528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_135_wb_clk_i_I clknet_4_9_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5497__S _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5944__B2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5944__A1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3280_ _1556_ _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_144_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5921_ net286 _0663_ _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_85_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_100_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _1306_ _1307_ _1311_ net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_76_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5783_ _1139_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ net408 _2781_ _2789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ net551 _2719_ _2720_ _2732_ _2733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4665_ net539 _2651_ _2652_ _2674_ _2675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_25_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ _0324_ clknet_leaf_29_wb_clk_i dffram.data\[50\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3616_ _1922_ _1930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4596_ _2550_ _2614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3547_ dffram.data\[57\]\[6\] _1880_ _1883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6335_ _0255_ clknet_leaf_144_wb_clk_i dffram.data\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input161_I qcpu_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input259_I sn76489_do[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3478_ _1451_ _1835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6266_ _0186_ clknet_leaf_40_wb_clk_i dffram.data\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5217_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6197_ _0117_ clknet_leaf_100_wb_clk_i dffram.data\[30\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input22_I ay8913_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__B1 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5148_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_4_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5079_ _2937_ _2985_ _2987_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5926__B2 net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output478_I net478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4450_ _2408_ _2492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3401_ _1784_ _1781_ _1785_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4381_ net415 _2436_ _2441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _0040_ clknet_leaf_15_wb_clk_i dffram.data\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3332_ dffram.data\[31\]\[7\] _1735_ _1739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3263_ _1637_ _1690_ _1692_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6051_ net86 _1482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3194_ _1645_ _1642_ _1646_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5002_ dffram.data\[40\]\[7\] _2932_ _2936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5605__B1 _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4408__A1 net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__A1 _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _1117_ _1357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4833__I _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5835_ _1295_ _1296_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5908__A1 _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ _1132_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _1172_ _1179_ net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_118_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4717_ _2714_ _2718_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input376_I wbs_adr_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _2631_ _2660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3147__A1 _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3184__I _1622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4579_ net560 _2583_ _2599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6318_ _0238_ clknet_leaf_145_wb_clk_i dffram.data\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5519__S0 _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6249_ _0169_ clknet_leaf_66_wb_clk_i dffram.data\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5072__A1 _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4743__I _2624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5462__I3 dffram.data\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3359__I _1756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5127__A2 _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3094__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput361 ue1_do[4] net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput350 tholin_riscv_oeb[3] net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput372 net621 net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_117_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput383 net579 net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput394 net612 net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold90 wbs_dat_i[0] net668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _2145_ _2152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_133_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3881_ dffram.data\[21\]\[4\] _2106_ _2107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _0623_ _0658_ _1108_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_73_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5551_ _1052_ _1053_ _0736_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4502_ _2520_ _2531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5482_ _0985_ _0986_ _0769_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4433_ _2468_ _2480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_130_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4364_ net408 _2406_ _2428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3315_ _1727_ _1729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4295_ dffram.data\[44\]\[2\] _2376_ _2379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6103_ _0023_ clknet_leaf_86_wb_clk_i dffram.data\[37\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3732__I _1998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5826__B1 _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3246_ _1647_ _1677_ _1681_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6034_ _1463_ _1464_ _1466_ _1457_ _1467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_83_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3177_ dffram.data\[63\]\[5\] _1632_ _1634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input124_I pdp11_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _1229_ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_107_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5749_ _1217_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3368__A1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3907__I _2118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__A2 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_105_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3540__A1 _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output510_I net510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4556__B1 _2576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold78_I wbs_cyc_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3817__I _2061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4859__A1 _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__B1 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ _1485_ _1581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4080_ _2237_ _2230_ _2238_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3031_ _1453_ _1528_ _1531_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput180 qcpu_do[32] net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput191 qcpu_oeb[12] net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A2 _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _2538_ _2918_ _2923_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_3_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3933_ dffram.data\[19\]\[5\] _2140_ _2142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_154_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6652_ _0572_ clknet_leaf_79_wb_clk_i dffram.data\[41\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3864_ _2089_ _2091_ _2093_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5603_ _1104_ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4547__B1 _2569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3795_ _2048_ _2049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _0503_ clknet_leaf_121_wb_clk_i net564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_132_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5534_ dffram.data\[0\]\[6\] dffram.data\[2\]\[6\] dffram.data\[4\]\[6\] dffram.data\[6\]\[6\]
+ _0975_ _0976_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_5465_ dffram.data\[9\]\[4\] dffram.data\[11\]\[4\] dffram.data\[13\]\[4\] dffram.data\[15\]\[4\]
+ _0848_ _0849_ _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_30_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ net390 _2466_ _2467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5396_ _0901_ _0902_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3522__A1 dffram.data\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input241_I sid_do[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3462__I _1816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4347_ net402 _2409_ _2415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input339_I tholin_riscv_oeb[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4278_ _2361_ _2368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_158_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _1451_ _1452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3229_ _1663_ _1671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_129_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__I _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3637__I _1936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output558_I net558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3761__A1 _1981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output460_I net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3513__A1 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_73_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5018__A1 _2946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__A2 _1071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5974__C1 net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_15_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5726__C1 net344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A2 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3580_ _1835_ _1905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5250_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4201_ dffram.data\[1\]\[1\] _2316_ _2318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5181_ net224 _0647_ _0690_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_147_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4132_ _2225_ _2267_ _2271_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4063_ _2225_ _2220_ _2226_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3014_ dffram.data\[35\]\[6\] _1516_ _1519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A1 _2937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4965_ dffram.data\[41\]\[0\] _2913_ _2914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5280__I1 _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _2115_ _2125_ _2130_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5980__A2 _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _2761_ _2864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3847_ _2035_ _2076_ _2081_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _0555_ clknet_leaf_105_wb_clk_i wb_counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input289_I tbb1143_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _0486_ clknet_leaf_74_wb_clk_i dffram.data\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input191_I qcpu_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3778_ _2035_ _2028_ _2036_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3743__A1 _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _1019_ _1020_ _0735_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6497_ _0417_ clknet_leaf_73_wb_clk_i dffram.data\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_167_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input52_I mc14500_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _0952_ _0953_ _0875_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput462 net462 io_oeb[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput451 net451 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput440 net440 custom_settings[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput495 net495 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput484 net484 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5379_ dffram.data\[25\]\[2\] dffram.data\[27\]\[2\] dffram.data\[29\]\[2\] dffram.data\[31\]\[2\]
+ _0832_ _0834_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput473 net473 io_oeb[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5799__A2 _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__I _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmultiplexer_575 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__6008__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_120_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_146_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A1 _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_94_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3734__A1 _1975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_155_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4198__I _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5334__S1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_164_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_158_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__C1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A2 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _2548_ wb_counter\[29\] _2746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ _1985_ _1987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4681_ _2615_ _2688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _1905_ _1937_ _1940_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6420_ _0340_ clknet_leaf_28_wb_clk_i dffram.data\[49\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _0271_ clknet_leaf_141_wb_clk_i dffram.data\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _0810_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3563_ _1886_ _1893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6282_ _0202_ clknet_leaf_45_wb_clk_i dffram.data\[56\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3494_ dffram.data\[58\]\[4\] _1847_ _1848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _0725_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4150__A1 _2279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__S1 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ net374 net75 _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4115_ dffram.data\[47\]\[4\] _2260_ _2261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5095_ _2956_ _2991_ _2996_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4046_ dffram.data\[4\]\[5\] _2213_ _2215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input204_I qcpu_oeb[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _1427_ _1432_ _1433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5953__A2 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4948_ dffram.data\[42\]\[2\] _2900_ _2903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ net392 _2850_ _2851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6618_ _0538_ clknet_leaf_129_wb_clk_i wb_counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6549_ _0469_ clknet_leaf_117_wb_clk_i net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5564__S1 _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output423_I net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3097__I _1563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__A1 _2109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3707__A1 _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold60_I wbs_dat_i[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4132__A1 _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5880__A1 net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5632__B2 net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ net267 _1260_ _1370_ net52 net98 _1343_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_85_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5851_ _1214_ _1308_ _1309_ _1310_ _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__A2 _1507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5935__A2 _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5782_ _1102_ _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ wb_counter\[6\] _2787_ _2788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_145_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4733_ _2730_ _2731_ _2732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6403_ _0323_ clknet_leaf_30_wb_clk_i dffram.data\[50\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ _2627_ _2671_ _2673_ _2674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3615_ _1922_ _1929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4595_ net562 _2613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3546_ _1850_ _1879_ _1882_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6334_ _0254_ clknet_leaf_144_wb_clk_i dffram.data\[23\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6265_ _0185_ clknet_leaf_39_wb_clk_i dffram.data\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input154_I pdp11_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5950__I _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3477_ _1830_ _1832_ _1834_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5216_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5871__A1 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _0116_ clknet_leaf_69_wb_clk_i dffram.data\[30\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input321_I tholin_riscv_do[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5147_ _0658_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_4_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5078_ dffram.data\[9\]\[0\] _2986_ _2987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input15_I ay8913_do[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ dffram.data\[49\]\[7\] _2200_ _2204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5397__I _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5862__A1 net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5100__I net578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3928__A1 _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3400_ dffram.data\[28\]\[5\] _1782_ _1785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4380_ _2439_ net601 _2435_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3331_ _1720_ _1734_ _1738_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3262_ dffram.data\[6\]\[0\] _1691_ _1692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6050_ _1472_ _1479_ _1481_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I ay8913_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3193_ dffram.data\[62\]\[1\] _1643_ _1646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5001_ _2536_ _2931_ _2935_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4656__A2 _2664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__B2 net324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A1 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5903_ net8 _1312_ _1334_ net96 _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_152_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ net254 _1229_ _1232_ net71 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_14_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5765_ _1232_ _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5696_ net198 _1174_ _1178_ net132 net334 _1175_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_20_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4592__A1 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ net548 _2697_ _2698_ _2717_ _2718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_135_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4647_ _2653_ wb_counter\[13\] _2659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input271_I sn76489_do[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4578_ _2591_ _2598_ _2574_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_9_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _0237_ clknet_leaf_9_wb_clk_i dffram.data\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _1856_ _1866_ _1871_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5519__S1 _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _0168_ clknet_leaf_21_wb_clk_i dffram.data\[58\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5844__A1 net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _0099_ clknet_leaf_71_wb_clk_i dffram.data\[32\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_98_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output490_I net490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_27_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4583__A1 _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4335__A1 net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput362 ue1_do[5] net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput340 tholin_riscv_oeb[24] net340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput351 tholin_riscv_oeb[4] net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput384 net594 net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput395 net641 net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput373 wbs_adr_i[2] net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold91 wbs_dat_i[8] net669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_37_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5446__S0 _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3880_ _2090_ _2106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5550_ dffram.data\[57\]\[7\] dffram.data\[59\]\[7\] dffram.data\[61\]\[7\] dffram.data\[63\]\[7\]
+ _0724_ _0727_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_152_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ dffram.data\[32\]\[5\] dffram.data\[34\]\[5\] dffram.data\[36\]\[5\] dffram.data\[38\]\[5\]
+ _0758_ _0760_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_4501_ _1478_ _2530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4602__C _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4432_ net395 _2478_ _2479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_113_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4363_ net442 _2427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3314_ _1727_ _1728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4294_ _2345_ _2375_ _2378_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6102_ _0022_ clknet_leaf_86_wb_clk_i dffram.data\[37\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5826__B2 net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5826__A1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3245_ dffram.data\[61\]\[2\] _1678_ _1681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6033_ net405 _1465_ _1466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3176_ _1577_ _1631_ _1633_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_159_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input117_I pdp11_do[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5054__A2 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3065__A1 _1487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5817_ net281 _1278_ _1266_ net24 _1280_ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_137_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5748_ _1216_ _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input82_I mc14500_sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5679_ _1123_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_145_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_145_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5817__A1 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5817__B2 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output503_I net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__S0 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4859__A2 _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5808__B2 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__A1 net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3295__A1 _1712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ dffram.data\[37\]\[1\] _1529_ _1531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput181 qcpu_do[3] net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput170 qcpu_do[23] net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput192 qcpu_oeb[13] net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4981_ dffram.data\[41\]\[7\] _2919_ _2923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_13_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3932_ _2104_ _2139_ _2141_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _0571_ clknet_leaf_84_wb_clk_i dffram.data\[41\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3863_ dffram.data\[21\]\[0\] _2092_ _2093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5602_ _0651_ _0667_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6582_ _0502_ clknet_leaf_121_wb_clk_i net563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3794_ _2047_ _1935_ _2048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5533_ dffram.data\[8\]\[6\] dffram.data\[10\]\[6\] dffram.data\[12\]\[6\] dffram.data\[14\]\[6\]
+ _0937_ _0938_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_27_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _0966_ _0969_ _0846_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5395_ _0746_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4415_ _2430_ _2466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_169_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4346_ _2413_ _2407_ _2414_ _2412_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4277_ _2349_ _2362_ _2367_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3286__A1 _1702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3228_ _1663_ _1670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input234_I qcpu_sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ net229 _1438_ _1450_ _1451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5680__C1 net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3159_ _1588_ _1616_ _1621_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5983__B1 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output453_I net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3277__A1 _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_42_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3029__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold90_I wbs_dat_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__I0 dffram.data\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I _2418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4200_ _2279_ _2315_ _2317_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3563__I _1886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _0687_ _0689_ _0646_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_147_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4131_ dffram.data\[20\]\[2\] _2268_ _2271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4062_ dffram.data\[48\]\[2\] _2221_ _2226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_108_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3013_ _1487_ _1515_ _1518_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__B1 _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _2911_ _2913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3915_ dffram.data\[51\]\[7\] _2126_ _2130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4895_ _2841_ _2862_ _2863_ _2854_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_144_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3846_ dffram.data\[52\]\[3\] _2077_ _2081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6634_ _0554_ clknet_leaf_116_wb_clk_i wb_counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3777_ dffram.data\[53\]\[3\] _2029_ _2036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6565_ _0485_ clknet_leaf_147_wb_clk_i design_select\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3743__A2 _2012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ dffram.data\[57\]\[6\] dffram.data\[59\]\[6\] dffram.data\[61\]\[6\] dffram.data\[63\]\[6\]
+ _0739_ _0740_ _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _0416_ clknet_leaf_91_wb_clk_i dffram.data\[45\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input184_I qcpu_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ dffram.data\[57\]\[4\] dffram.data\[59\]\[4\] dffram.data\[61\]\[4\] dffram.data\[63\]\[4\]
+ _0872_ _0873_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_input351_I tholin_riscv_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput430 net430 custom_settings[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput441 net441 custom_settings[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput452 net452 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput485 net485 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput496 net496 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input45_I mc14500_do[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ dffram.data\[17\]\[2\] dffram.data\[19\]\[2\] dffram.data\[21\]\[2\] dffram.data\[23\]\[2\]
+ _0884_ _0885_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput463 net463 io_oeb[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput474 net474 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_35_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4329_ _2359_ _2394_ _2399_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3259__A1 _1608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xmultiplexer_565 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmultiplexer_576 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_TAPCELL_ROW_2_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__A3 _2403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A3 _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3648__I _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5947__B1 _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4942__I _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _1985_ _1986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3422__A1 _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4680_ _2686_ wb_counter\[18\] _2687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3631_ dffram.data\[11\]\[1\] _1938_ _1940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3562_ _1842_ _1887_ _1892_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6350_ _0270_ clknet_leaf_141_wb_clk_i dffram.data\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5301_ _0691_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I _2422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _0201_ clknet_leaf_41_wb_clk_i dffram.data\[56\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3493_ _1831_ _1847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3489__A1 _1842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _0738_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5163_ _0659_ design_select\[2\] design_select\[0\] _0621_ _0673_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_127_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4114_ _2252_ _2260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5094_ dffram.data\[9\]\[7\] _2992_ _2996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4989__A1 _2524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4045_ _2169_ _2212_ _2214_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5650__A2 _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3661__A1 _1911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__I _2768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _1062_ _1431_ _1432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3413__A1 dffram.data\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4947_ _2524_ _2899_ _2902_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _2763_ _2850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_160_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6617_ _0537_ clknet_leaf_125_wb_clk_i wb_counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3829_ _2037_ _2068_ _2070_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4913__A1 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4299__I _2374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _0468_ clknet_leaf_126_wb_clk_i net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6479_ _0399_ clknet_leaf_109_wb_clk_i dffram.data\[46\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output416_I net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3404__A1 _1786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5593__I _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5632__A2 _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5850_ net256 _1269_ _1254_ net73 _1310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__C _1522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ net249 _1247_ _1181_ net313 _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_14_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4801_ _2593_ wb_counter\[5\] _2778_ _2787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_72_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4732_ net432 _2688_ _2726_ _2731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4663_ net420 _2665_ _2672_ _2673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5699__A2 _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3614_ _1909_ _1923_ _1928_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6402_ _0322_ clknet_leaf_39_wb_clk_i dffram.data\[50\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ _2606_ _2612_ _2605_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3545_ dffram.data\[57\]\[5\] _1880_ _1882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6333_ _0253_ clknet_leaf_144_wb_clk_i dffram.data\[23\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_164_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3476_ dffram.data\[58\]\[0\] _1833_ _1834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6264_ _0184_ clknet_leaf_21_wb_clk_i dffram.data\[57\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5215_ _0680_ _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6195_ _0115_ clknet_leaf_69_wb_clk_i dffram.data\[30\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input147_I pdp11_oeb[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__A2 _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5146_ _0660_ design_select\[2\] _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3882__A1 _2104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _2984_ _2986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input314_I tholin_riscv_do[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ _2175_ _2199_ _2203_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3634__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ net178 _1413_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_133_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__A1 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output533_I net533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_100_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3330_ dffram.data\[31\]\[6\] _1735_ _1738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4667__I _2582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3261_ _1689_ _1691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5000_ dffram.data\[40\]\[6\] _2932_ _2935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3192_ _1567_ _1645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3864__A1 _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A2 _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5902_ net162 _1262_ _1264_ net50 _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_53_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5833_ net26 _1225_ _1170_ net38 _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_53_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5764_ _1205_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4041__A1 _2167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5695_ _1177_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_60_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4715_ _2699_ _2715_ _2716_ _2717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _2645_ _2658_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4577_ _2592_ _2596_ _2597_ _2598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_124_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6316_ _0236_ clknet_leaf_53_wb_clk_i dffram.data\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_9_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input264_I sn76489_do[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3528_ dffram.data\[26\]\[7\] _1867_ _1871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3459_ dffram.data\[5\]\[3\] _1818_ _1822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6247_ _0167_ clknet_leaf_20_wb_clk_i dffram.data\[58\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6178_ _0098_ clknet_leaf_71_wb_clk_i dffram.data\[32\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3855__A1 _2043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _0632_ _0647_ net526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_58_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_40_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5201__I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_12_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output483_I net483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4099__A1 _2235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput330 tholin_riscv_oeb[15] net330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5835__A2 _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__S0 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput341 tholin_riscv_oeb[25] net341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput352 tholin_riscv_oeb[5] net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput363 ue1_do[6] net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold16_I wbs_dat_i[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput385 net582 net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold70 net670 net647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput396 net645 net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold92 wbs_dat_i[7] net670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput374 wbs_adr_i[3] net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4271__A1 _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A2 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5446__S1 _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4500_ _2528_ _2521_ _2529_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5480_ dffram.data\[40\]\[5\] dffram.data\[42\]\[5\] dffram.data\[44\]\[5\] dffram.data\[46\]\[5\]
+ _0865_ _0866_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_152_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4431_ _2430_ _2478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_1 _2219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _2425_ _2423_ _2426_ _2420_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4293_ dffram.data\[44\]\[1\] _2376_ _2378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3313_ _1724_ _1726_ _1727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6101_ _0021_ clknet_leaf_87_wb_clk_i dffram.data\[37\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3244_ _1645_ _1677_ _1680_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6032_ _1203_ _1465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__A1 _2074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3175_ dffram.data\[63\]\[4\] _1632_ _1633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_159_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5021__I _2938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5816_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_137_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4014__A1 _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5747_ _1204_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_130_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_144_wb_clk_i_I clknet_4_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5678_ _1160_ _1165_ net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input75_I mc14500_sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ net534 _2623_ _2626_ _2643_ _2644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5817__A2 _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3828__A1 dffram.data\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_114_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_135_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__I _2761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__S1 _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4005__A1 _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5106__I _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3819__A1 _2026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput160 qcpu_do[14] net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput171 qcpu_do[24] net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_37_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput193 qcpu_oeb[14] net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput182 qcpu_do[4] net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_37_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4980_ _2536_ _2918_ _2922_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3931_ dffram.data\[19\]\[4\] _2140_ _2141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _0570_ clknet_leaf_79_wb_clk_i dffram.data\[41\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3862_ _2090_ _2092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5744__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5601_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_129_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6581_ _0501_ clknet_leaf_128_wb_clk_i net562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_144_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3793_ _1525_ _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5532_ _1034_ _1035_ _0788_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__I1 _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _0967_ _0968_ _0893_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5394_ dffram.data\[0\]\[2\] dffram.data\[2\]\[2\] dffram.data\[4\]\[2\] dffram.data\[6\]\[2\]
+ _0785_ _0786_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ net424 _2458_ _2465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4345_ net391 _2409_ _2414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4276_ dffram.data\[18\]\[3\] _2363_ _2367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3227_ _1649_ _1664_ _1669_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6015_ _1448_ _1216_ _1449_ _1101_ _1450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4483__A1 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3158_ dffram.data\[0\]\[7\] _1617_ _1621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input227_I qcpu_sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3089_ _1571_ _1564_ _1572_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4235__A1 _2296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5983__A1 net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output446_I net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5974__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__B2 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__I _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_82_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5726__A1 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold83_I wbs_dat_i[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__B2 net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__I1 dffram.data\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4130_ _2223_ _2267_ _2270_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_147_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4061_ _2097_ _2225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_108_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3012_ dffram.data\[35\]\[5\] _1516_ _1518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4217__A1 _2047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__A1 net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4963_ _2911_ _2912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3914_ _2112_ _2125_ _2129_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4894_ net395 _2844_ _2863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6633_ _0553_ clknet_leaf_135_wb_clk_i wb_counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _2033_ _2076_ _2080_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3776_ _1841_ _2035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6564_ _0484_ clknet_leaf_147_wb_clk_i design_select\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6495_ _0415_ clknet_leaf_89_wb_clk_i dffram.data\[45\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5515_ dffram.data\[49\]\[6\] dffram.data\[51\]\[6\] dffram.data\[53\]\[6\] dffram.data\[55\]\[6\]
+ _0729_ _0731_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__3754__I _2013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5446_ dffram.data\[49\]\[4\] dffram.data\[51\]\[4\] dffram.data\[53\]\[4\] dffram.data\[55\]\[4\]
+ _0816_ _0817_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xoutput420 net420 custom_settings[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input177_I qcpu_do[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput431 net431 custom_settings[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput453 net453 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput442 net442 custom_settings[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input344_I tholin_riscv_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput486 net486 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_160_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5377_ _0833_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xoutput464 net464 io_oeb[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_1_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput475 net475 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_35_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput497 net497 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4328_ dffram.data\[17\]\[7\] _2395_ _2399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input38_I diceroll_do[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _2419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4259_ dffram.data\[16\]\[5\] _2353_ _2356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3259__A2 _1640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmultiplexer_566 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_167_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xmultiplexer_577 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__5956__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5500__S0 _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__I _2132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5971__A4 _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_34_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__I _1435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_69_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4447__A1 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__A1 net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5947__B2 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3839__I _2075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3630_ _1899_ _1937_ _1939_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_78_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3561_ dffram.data\[10\]\[3\] _1888_ _1892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ dffram.data\[32\]\[1\] dffram.data\[34\]\[1\] dffram.data\[36\]\[1\] dffram.data\[38\]\[1\]
+ _0807_ _0808_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_110_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_149_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _1831_ _1846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6280_ _0200_ clknet_leaf_103_wb_clk_i dffram.data\[25\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_166_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ dffram.data\[56\]\[0\] dffram.data\[58\]\[0\] dffram.data\[60\]\[0\] dffram.data\[62\]\[0\]
+ _0739_ _0740_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_45_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _0666_ _0672_ net531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_127_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_87_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5093_ _2954_ _2991_ _2995_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4113_ _2252_ _2259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3110__A1 dffram.data\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4044_ dffram.data\[4\]\[4\] _2213_ _2214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5238__I0 _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5995_ _1428_ _0751_ _1429_ _1430_ net368 _1431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_96_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4946_ dffram.data\[42\]\[1\] _2900_ _2902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _2847_ _2848_ _2796_ _2849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input294_I tholin_riscv_do[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6616_ _0536_ clknet_leaf_128_wb_clk_i wb_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ dffram.data\[22\]\[4\] _2069_ _2070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6547_ _0467_ clknet_leaf_122_wb_clk_i net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_132_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3759_ _1979_ _2020_ _2023_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6478_ _0398_ clknet_leaf_110_wb_clk_i dffram.data\[46\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ _0934_ _0935_ _0852_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__B _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__I _1949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3168__A1 _1568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold46_I wbs_adr_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__S _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_105_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5093__A1 _2954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_122_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__I _2898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_122_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _2777_ _2784_ _2785_ _2786_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_146_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ _1229_ _1247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_127_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4731_ _2686_ wb_counter\[26\] _2730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4662_ _2630_ _2672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3613_ dffram.data\[56\]\[3\] _1924_ _1928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6401_ _0321_ clknet_leaf_29_wb_clk_i dffram.data\[50\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3159__A1 _1588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4593_ _2592_ _2610_ _2611_ _2612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6332_ _0252_ clknet_leaf_54_wb_clk_i dffram.data\[23\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3544_ _1845_ _1879_ _1881_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3475_ _1831_ _1833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6263_ _0183_ clknet_leaf_20_wb_clk_i dffram.data\[57\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5214_ _0723_ _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6194_ _0114_ clknet_leaf_72_wb_clk_i dffram.data\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3331__A1 _1720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5145_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5076_ _2984_ _2985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4027_ dffram.data\[49\]\[6\] _2200_ _2203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input307_I tholin_riscv_do[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _1387_ _1416_ _1417_ net503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_137_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__I _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3398__A1 _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_139_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_139_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4929_ wb_counter\[31\] _2888_ _2889_ _2890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4103__I _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3570__A1 _1853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5847__B1 _1097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output526_I net526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A1 _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__I _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4822__A1 net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3260_ _1689_ _1690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3313__A1 _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3191_ _1637_ _1642_ _1644_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5779__I _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ _1349_ _1350_ _1351_ _1354_ net489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_89_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5832_ net185 _1210_ _1097_ net119 _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_147_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5763_ net247 _1230_ _1122_ net166 _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_84_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_134_wb_clk_i_I clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4714_ net429 _2705_ _2710_ _2716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5694_ _1095_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4645_ net536 _2651_ _2652_ _2657_ _2658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _0624_ _2561_ _2597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6315_ _0235_ clknet_leaf_52_wb_clk_i dffram.data\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3552__A1 _1591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3527_ _1853_ _1866_ _1870_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input257_I sid_oeb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3458_ _1776_ _1817_ _1821_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6246_ _0166_ clknet_leaf_20_wb_clk_i dffram.data\[58\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3389_ dffram.data\[28\]\[2\] _1772_ _1777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6177_ _0097_ clknet_leaf_72_wb_clk_i dffram.data\[32\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input20_I ay8913_do[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_135_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ dffram.data\[39\]\[1\] _2973_ _2975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output476_I net476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3672__I _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput320 tholin_riscv_do[6] net320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput342 tholin_riscv_oeb[26] net342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput331 tholin_riscv_oeb[16] net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput353 tholin_riscv_oeb[6] net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5391__S1 _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput364 ue1_do[7] net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5599__I _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput386 net603 net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold71 net629 net648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput397 net643 net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold60 wbs_dat_i[25] net640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput375 wbs_adr_i[4] net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold82 _2404_ net660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold93 wbs_dat_i[29] net671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_37_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6494__CLK clknet_4_14_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4430_ net429 _2470_ _2477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_2 _2239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3534__A1 _1830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _0020_ clknet_leaf_80_wb_clk_i dffram.data\[37\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4361_ net407 _2406_ _2426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_130_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4292_ _2340_ _2375_ _2377_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3312_ _1725_ _1726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3243_ dffram.data\[61\]\[1\] _1678_ _1680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6031_ _1204_ _1464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_94_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _2942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3174_ _1624_ _1632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5302__I _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5815_ net117 _1115_ _1170_ net36 _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ _1086_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_88_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5677_ net193 _1163_ _1149_ net127 net329 _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_60_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input374_I wbs_adr_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4628_ _2641_ _2642_ _2643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input68_I mc14500_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3525__A1 _1850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3492__I _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _2575_ _2581_ _2574_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _0149_ clknet_leaf_16_wb_clk_i dffram.data\[60\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__I _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_97_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput150 pdp11_oeb[5] net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput161 qcpu_do[15] net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput172 qcpu_do[25] net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput194 qcpu_oeb[15] net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput183 qcpu_do[5] net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5977__C1 net312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _2132_ _2140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_154_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3577__I _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3861_ _2090_ _2091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5744__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5600_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3792_ _2045_ _2038_ _2046_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6580_ _0500_ clknet_leaf_130_wb_clk_i net561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_109_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5531_ dffram.data\[1\]\[6\] dffram.data\[3\]\[6\] dffram.data\[5\]\[6\] dffram.data\[7\]\[6\]
+ _0782_ _0783_ _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_54_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3507__A1 _1856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ dffram.data\[16\]\[4\] dffram.data\[18\]\[4\] dffram.data\[20\]\[4\] dffram.data\[22\]\[4\]
+ _0795_ _0797_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5393_ dffram.data\[8\]\[2\] dffram.data\[10\]\[2\] dffram.data\[12\]\[2\] dffram.data\[14\]\[2\]
+ _0782_ _0783_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_68_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4413_ _2463_ net610 _2457_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4344_ net425 _2413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4275_ _2347_ _2362_ _2366_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6014_ net391 _1440_ _1449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5680__A1 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3226_ dffram.data\[33\]\[3\] _1665_ _1669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5680__B2 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3157_ _1585_ _1616_ _1620_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input122_I pdp11_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3088_ dffram.data\[7\]\[2\] _1565_ _1572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4871__I _2780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5729_ _1186_ _1201_ net470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3746__A1 dffram.data\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_107_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _2145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output439_I net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5974__A2 _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3985__A1 _2175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_125_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_51_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_110_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4021__I _2192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4060_ _2223_ _2220_ _2224_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3011_ _1479_ _1515_ _1517_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5965__A2 _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4962_ _2300_ _1662_ _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_74_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3913_ dffram.data\[51\]\[6\] _2126_ _2129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4893_ _2859_ _2861_ _2862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3844_ dffram.data\[52\]\[2\] _2077_ _2080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3100__I _1485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6632_ _0552_ clknet_leaf_116_wb_clk_i wb_counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3728__A1 _1971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3775_ _2033_ _2028_ _2034_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6563_ _0483_ clknet_leaf_147_wb_clk_i design_select\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _1014_ _1017_ _0914_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _0414_ clknet_4_14_0_wb_clk_i dffram.data\[45\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_160_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5445_ _0947_ _0950_ _0914_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4153__A1 _2284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput432 net432 custom_settings[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput421 net421 custom_settings[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput443 net443 custom_settings[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput487 net487 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3900__A1 _2089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput465 net465 io_oeb[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput476 net476 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_22_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput454 net454 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput498 net498 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_61_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4327_ _2357_ _2394_ _2398_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input337_I tholin_riscv_oeb[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4258_ _1486_ _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3209_ _1584_ _1657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xmultiplexer_567 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_4189_ _2290_ _2308_ _2310_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5500__S1 _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3719__A1 _1983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4144__A1 _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5495__I1 dffram.data\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ _1839_ _1887_ _1891_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5230_ _0730_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3491_ _1844_ _1845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_166_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5883__A1 net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5161_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__3590__I _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4112_ _2227_ _2253_ _2258_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5092_ dffram.data\[9\]\[6\] _2992_ _2995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_142_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_127_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _2205_ _2213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__B1 _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5994_ wb_sram_we _0624_ _0658_ _0660_ _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3949__A1 _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4945_ _2519_ _2899_ _2901_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__A1 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4876_ _2693_ _2842_ _2700_ _2848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3827_ _2061_ _2069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6615_ _0535_ clknet_leaf_128_wb_clk_i wb_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input287_I tbb1143_do[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6546_ _0466_ clknet_leaf_122_wb_clk_i net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3758_ dffram.data\[23\]\[5\] _2021_ _2023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6477_ _0397_ clknet_leaf_108_wb_clk_i dffram.data\[46\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3689_ _1975_ _1976_ _1978_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input50_I mc14500_do[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ dffram.data\[1\]\[3\] dffram.data\[3\]\[3\] dffram.data\[5\]\[3\] dffram.data\[7\]\[3\]
+ _0897_ _0898_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_100_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5874__A1 _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5359_ dffram.data\[40\]\[2\] dffram.data\[42\]\[2\] dffram.data\[44\]\[2\] dffram.data\[46\]\[2\]
+ _0865_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4596__I _2550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4545__B _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__I _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5929__A2 _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5485__S0 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__I _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5165__I0 net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A1 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__B2 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5130__I _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_10_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ _2714_ _2729_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4661_ wb_counter\[15\] _2671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_154_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3612_ _1907_ _1923_ _1927_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6400_ _0320_ clknet_leaf_23_wb_clk_i dffram.data\[59\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _0251_ clknet_leaf_54_wb_clk_i dffram.data\[23\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _0639_ _2561_ _2611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3543_ dffram.data\[57\]\[4\] _1880_ _1881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3474_ _1831_ _1832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4108__A1 _2223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6262_ _0182_ clknet_leaf_21_wb_clk_i dffram.data\[57\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6193_ _0113_ clknet_leaf_72_wb_clk_i dffram.data\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5213_ _0722_ _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__I _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5144_ design_select\[3\] _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5608__A1 _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__I1 dffram.data\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5075_ _1591_ _1900_ _2984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4026_ _2173_ _2199_ _2202_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input202_I qcpu_oeb[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A1 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5977_ net64 _1218_ _1116_ net110 net312 _1118_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_17_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ wb_counter\[31\] _2888_ _2763_ _2889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input98_I pdp11_do[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4859_ _2664_ _2671_ _2822_ _2833_ _2834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4347__A1 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5416__S _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6529_ _0449_ clknet_leaf_137_wb_clk_i net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_160_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__I _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output421_I net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output519_I net519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _1900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_67_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6046__I _1477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 _1455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__S0 _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__I0 _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3190_ dffram.data\[62\]\[0\] _1643_ _1644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4964__I _2911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3077__A1 _1559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ net95 _1255_ _1219_ net297 _1353_ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__A2 _2628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__S0 _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6015__A1 _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ net283 _1223_ _1234_ net321 _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5795__I _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ _1229_ _1230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_57_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4713_ wb_counter\[23\] _2715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_155_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5693_ _1172_ _1176_ net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_115_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4644_ _2654_ _2656_ _2657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3001__A1 _1445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4575_ _2566_ _2593_ _2594_ _2595_ _2587_ _2596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6314_ _0234_ clknet_leaf_40_wb_clk_i dffram.data\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3552__A2 _1885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3526_ dffram.data\[26\]\[6\] _1867_ _1870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5829__A1 net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6245_ _0165_ clknet_leaf_21_wb_clk_i dffram.data\[58\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input152_I pdp11_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3457_ dffram.data\[5\]\[2\] _1818_ _1821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5035__I _2958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3388_ _1570_ _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6176_ _0096_ clknet_leaf_23_wb_clk_i dffram.data\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5127_ _0643_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5058_ _2937_ _2972_ _2974_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I ay8913_do[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ _2177_ _2186_ _2191_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6006__A1 _1439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__I _2252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output469_I net469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput310 tholin_riscv_do[27] net310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput321 tholin_riscv_do[7] net321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput343 tholin_riscv_oeb[27] net343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput332 tholin_riscv_oeb[17] net332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput354 tholin_riscv_oeb[7] net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold50 net637 net627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput365 ue1_do[8] net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold61 net672 net638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput387 net615 net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold72 net664 net649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput376 wbs_adr_i[5] net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold83 wbs_dat_i[30] net661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3059__A1 _1470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput398 net644 net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold94 wbs_dat_i[28] net672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_98_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5548__C _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3231__A1 _1651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6639__CLK clknet_4_8_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_152_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_3 net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ net441 _2425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_130_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3311_ _1540_ _0773_ _1725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4291_ dffram.data\[44\]\[0\] _2376_ _2377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3242_ _1637_ _1677_ _1679_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6030_ net84 _1463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA_input5_I ay8913_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__C1 net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3173_ _1624_ _1631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4694__I _2618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__A1 net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3470__A1 _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5814_ _1259_ _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5745_ net29 _0627_ _1213_ _1214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5676_ _1145_ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__A1 _2526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4627_ net415 _2616_ _2637_ _2642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input367_I ue1_oeb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4722__A1 _2619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4558_ _2545_ _2579_ _2580_ _2581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_25_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4489_ _2520_ _2522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3509_ _1858_ _1755_ _1859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_38_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6228_ _0148_ clknet_leaf_36_wb_clk_i dffram.data\[60\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3289__A1 _1708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__C1 net331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6159_ _0079_ clknet_leaf_92_wb_clk_i dffram.data\[33\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__B _2605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4553__B _2568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5738__B1 _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_97_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4961__A1 _2538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput140 pdp11_oeb[26] net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput151 pdp11_oeb[6] net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput162 qcpu_do[16] net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput195 qcpu_oeb[16] net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput173 qcpu_do[26] net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput184 qcpu_do[6] net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_76_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3858__I _1443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4463__B _2501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _2047_ _2012_ _2090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3791_ dffram.data\[53\]\[7\] _2039_ _2046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5744__A3 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5530_ dffram.data\[9\]\[6\] dffram.data\[11\]\[6\] dffram.data\[13\]\[6\] dffram.data\[15\]\[6\]
+ _0776_ _0778_ _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_15_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5461_ dffram.data\[24\]\[4\] dffram.data\[26\]\[4\] dffram.data\[28\]\[4\] dffram.data\[30\]\[4\]
+ _0889_ _0890_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_48_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4412_ net389 _2455_ _2464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5392_ _0896_ _0899_ _0852_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4343_ _2400_ _2407_ _2410_ _2412_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_169_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4274_ dffram.data\[18\]\[2\] _2363_ _2366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3225_ _1647_ _1664_ _1668_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6013_ net82 _1448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_119_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3156_ dffram.data\[0\]\[6\] _1617_ _1620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3087_ _1570_ _1571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input115_I pdp11_do[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3443__A1 _1780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4373__B _2435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A1 _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ net209 _1197_ _1183_ net143 net345 _1198_ _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_116_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3989_ _2047_ _1858_ _2179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_73_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input80_I mc14500_sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4599__I _2553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _1148_ _1150_ net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3008__I _1508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__A1 _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output501_I net501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_91_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__C _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_147_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3010_ dffram.data\[35\]\[4\] _1516_ _1517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _2538_ _2905_ _2910_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3912_ _2109_ _2125_ _2128_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4892_ _2715_ _2860_ _2861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3843_ _2031_ _2076_ _2079_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6631_ _0551_ clknet_leaf_127_wb_clk_i wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5568__I3 dffram.data\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4925__A1 net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3774_ dffram.data\[53\]\[2\] _2029_ _2034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _0482_ clknet_leaf_147_wb_clk_i design_select\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5308__I _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5513_ _1015_ _1016_ _0769_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _0413_ clknet_leaf_89_wb_clk_i dffram.data\[45\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5444_ _0948_ _0949_ _0769_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput433 net433 custom_settings[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput422 net422 custom_settings[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput444 net444 custom_settings[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_5375_ _0826_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput466 net466 io_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput477 net477 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_35_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput455 net455 io_oeb[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput499 net499 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput488 net488 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4326_ dffram.data\[17\]\[6\] _2395_ _2398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4257_ _2351_ _2352_ _2354_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3208_ _1655_ _1652_ _1656_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4188_ dffram.data\[46\]\[4\] _2309_ _2310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input232_I qcpu_sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3139_ _1608_ _1594_ _1609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xmultiplexer_568 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3416__A1 _1776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output451_I net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__I _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3655__A1 _1907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3407__A1 _1788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_11_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4080__A1 _2237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__I _2205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3490_ _1477_ _1844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_149_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5160_ _0660_ _0642_ _0638_ _0644_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__3894__A1 _2115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4111_ dffram.data\[47\]\[3\] _2254_ _2258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5091_ _2952_ _2991_ _2994_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_127_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4042_ _2205_ _2212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A1 _1919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5993_ net80 _1203_ _1429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4944_ dffram.data\[42\]\[0\] _2900_ _2901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4207__I _2314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__A1 _2229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ wb_counter\[18\] wb_counter\[19\] wb_counter\[20\] _2834_ _2847_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_117_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6614_ _0534_ clknet_leaf_128_wb_clk_i wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3826_ _2061_ _2068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6545_ _0465_ clknet_leaf_122_wb_clk_i net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3757_ _1975_ _2020_ _2022_ _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input182_I qcpu_do[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _0396_ clknet_leaf_83_wb_clk_i dffram.data\[46\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3688_ dffram.data\[55\]\[4\] _1977_ _1978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5427_ dffram.data\[9\]\[3\] dffram.data\[11\]\[3\] dffram.data\[13\]\[3\] dffram.data\[15\]\[3\]
+ _0848_ _0849_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3781__I _2027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input43_I mc14500_do[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _0759_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4309_ _1900_ _2265_ _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_138_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5289_ dffram.data\[41\]\[1\] dffram.data\[43\]\[1\] dffram.data\[45\]\[1\] dffram.data\[47\]\[1\]
+ _0795_ _0797_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__S1 _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output499_I net499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5562__A1 _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3876__A1 _2101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4053__A1 _1921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3800__A1 _2031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ _2669_ _2670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3611_ dffram.data\[56\]\[2\] _1924_ _1927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5553__A1 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6330_ _0250_ clknet_leaf_54_wb_clk_i dffram.data\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4591_ _2557_ wb_counter\[6\] _2607_ _2609_ _2587_ _2610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3542_ _1872_ _1880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3473_ _1638_ _1755_ _1831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6261_ _0181_ clknet_leaf_21_wb_clk_i dffram.data\[57\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5212_ _0675_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6192_ _0112_ clknet_leaf_100_wb_clk_i dffram.data\[31\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5143_ _0645_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _2956_ _2978_ _2983_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4292__A1 _2340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4025_ dffram.data\[49\]\[5\] _2200_ _2202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5976_ net176 _1413_ _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_87_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5792__A1 _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4927_ _2741_ wb_counter\[29\] wb_counter\[30\] _2879_ _2888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_90_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ wb_counter\[16\] wb_counter\[17\] _2833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5544__A1 _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3809_ dffram.data\[13\]\[5\] _2056_ _2058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4789_ _2776_ _2777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _0448_ clknet_leaf_104_wb_clk_i dffram.data\[17\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _0379_ clknet_leaf_63_wb_clk_i dffram.data\[20\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5847__A2 _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4400__I _2431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4283__A1 _2355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output414_I net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_67_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A2 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__S1 _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4035__A1 _2158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3686__I _1965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__I _2387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3077__A2 _1562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__A2 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _1285_ _1286_ _1288_ _1292_ net480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_147_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5449__S1 _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__A1 _2173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5761_ _1086_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4712_ _2669_ _2714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5692_ net197 _1174_ _1166_ net131 net333 _1175_ _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_127_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5517__S _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ net417 _2655_ _2637_ _2656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_135_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _2421_ _2555_ _2577_ _2595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6313_ _0233_ clknet_leaf_52_wb_clk_i dffram.data\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3525_ _1850_ _1866_ _1869_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6244_ _0164_ clknet_leaf_40_wb_clk_i dffram.data\[58\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3456_ _1774_ _1817_ _1820_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3387_ _1774_ _1771_ _1775_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _0095_ clknet_leaf_21_wb_clk_i dffram.data\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input145_I pdp11_oeb[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5126_ _0618_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5057_ dffram.data\[39\]\[0\] _2973_ _2974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input312_I tholin_riscv_do[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4008_ dffram.data\[29\]\[7\] _2187_ _2191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4265__A1 dffram.data\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__A2 _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5959_ _1396_ _1401_ _1402_ _1403_ net498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_149_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5226__I _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output531_I net531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput311 tholin_riscv_do[28] net311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput300 tholin_riscv_do[18] net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput344 tholin_riscv_oeb[28] net344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput333 tholin_riscv_oeb[18] net333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput322 tholin_riscv_do[8] net322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_101_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold40 wbs_dat_i[12] net620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput366 ue1_do[9] net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput355 tholin_riscv_oeb[8] net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput388 net630 net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xhold73 net662 net650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput377 wbs_adr_i[6] net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold51 _2500_ net628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold62 _2494_ net639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold84 wbs_dat_i[4] net662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold95 wbs_dat_i[27] net673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput399 net635 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4008__A1 dffram.data\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5300__S0 _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_4 _1901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3310_ _1561_ _1724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _2374_ _2376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3241_ dffram.data\[61\]\[0\] _1678_ _1679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3172_ _1574_ _1625_ _1630_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__B2 _1430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _1272_ _1273_ _1277_ net511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_119_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5744_ net41 _0653_ _0656_ _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_18_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5675_ _1162_ _1163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _2621_ wb_counter\[10\] _2641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input262_I sn76489_do[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ _0620_ _2562_ _2580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4488_ _2520_ _2521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3508_ _1725_ _1858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_38_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3439_ _1778_ _1804_ _1809_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6227_ _0147_ clknet_leaf_36_wb_clk_i dffram.data\[60\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _0078_ clknet_leaf_92_wb_clk_i dffram.data\[33\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_55_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ wb_override_act net42 _0630_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6089_ _0009_ clknet_leaf_78_wb_clk_i dffram.data\[35\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__S0 _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5738__A1 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__B2 net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4125__I _2266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output481_I net481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_75_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput141 pdp11_oeb[27] net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput152 pdp11_oeb[7] net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput130 pdp11_oeb[17] net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput163 qcpu_do[17] net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput196 qcpu_oeb[17] net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput174 qcpu_do[27] net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput185 qcpu_do[7] net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5977__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5977__B2 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3790_ _1855_ _2045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4401__A1 net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5460_ _0964_ _0965_ _0765_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_132_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4411_ net423 _2458_ _2463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5391_ dffram.data\[1\]\[2\] dffram.data\[3\]\[2\] dffram.data\[5\]\[2\] dffram.data\[7\]\[2\]
+ _0897_ _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_112_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4342_ _2411_ _2412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_169_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4273_ _2345_ _2362_ _2365_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5504__I1 _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3224_ dffram.data\[33\]\[2\] _1665_ _1668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6012_ _1436_ _1445_ _1447_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4468__A1 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

