VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_qcpu
  CLASS BLOCK ;
  FOREIGN wrapped_qcpu ;
  ORIGIN 0.000 0.000 ;
  SIZE 575.000 BY 600.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.000 4.000 56.560 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.000 4.000 224.560 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 240.800 4.000 241.360 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.400 4.000 274.960 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.200 4.000 291.760 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.000 4.000 308.560 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.400 4.000 358.960 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.200 4.000 375.760 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.000 4.000 392.560 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 408.800 4.000 409.360 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 425.600 4.000 426.160 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 442.400 4.000 442.960 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 459.200 4.000 459.760 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 492.800 4.000 493.360 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 526.400 4.000 526.960 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 543.200 4.000 543.760 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.600 4.000 90.160 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 576.800 4.000 577.360 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.200 4.000 123.760 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.400 4.000 190.960 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END custom_settings[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 596.000 33.040 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 596.000 111.440 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 596.000 119.280 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 596.000 127.120 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 596.000 134.960 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 596.000 142.800 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 596.000 150.640 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 596.000 158.480 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 596.000 166.320 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 596.000 174.160 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 596.000 182.000 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 596.000 40.880 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 596.000 189.840 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 596.000 197.680 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 596.000 205.520 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 596.000 213.360 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 596.000 221.200 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 596.000 229.040 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 596.000 236.880 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 596.000 244.720 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 596.000 252.560 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 596.000 260.400 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 596.000 48.720 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 596.000 268.240 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 596.000 276.080 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 596.000 283.920 600.000 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 596.000 56.560 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 596.000 64.400 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 596.000 72.240 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 596.000 80.080 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 596.000 87.920 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 596.000 95.760 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 596.000 103.600 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 22.400 575.000 22.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 123.200 575.000 123.760 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 133.280 575.000 133.840 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 143.360 575.000 143.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 153.440 575.000 154.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 163.520 575.000 164.080 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 173.600 575.000 174.160 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 183.680 575.000 184.240 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 193.760 575.000 194.320 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 203.840 575.000 204.400 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 213.920 575.000 214.480 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 32.480 575.000 33.040 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 224.000 575.000 224.560 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 234.080 575.000 234.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 244.160 575.000 244.720 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 254.240 575.000 254.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 264.320 575.000 264.880 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 274.400 575.000 274.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 284.480 575.000 285.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 294.560 575.000 295.120 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 304.640 575.000 305.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 314.720 575.000 315.280 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 42.560 575.000 43.120 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 324.800 575.000 325.360 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 334.880 575.000 335.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 344.960 575.000 345.520 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 52.640 575.000 53.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 62.720 575.000 63.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 72.800 575.000 73.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 82.880 575.000 83.440 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 92.960 575.000 93.520 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 103.040 575.000 103.600 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 113.120 575.000 113.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 596.000 291.760 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 596.000 370.160 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 596.000 378.000 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 596.000 385.840 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 596.000 393.680 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 596.000 401.520 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 596.000 409.360 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 596.000 417.200 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 596.000 425.040 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 596.000 432.880 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 596.000 440.720 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 596.000 299.600 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 596.000 448.560 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 596.000 456.400 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 596.000 464.240 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 596.000 472.080 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 596.000 479.920 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 596.000 487.760 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 596.000 495.600 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 596.000 503.440 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 596.000 511.280 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 596.000 519.120 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 596.000 307.440 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 596.000 526.960 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 596.000 534.800 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 596.000 542.640 600.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 596.000 315.280 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 596.000 323.120 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 596.000 330.960 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 596.000 338.800 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 596.000 346.640 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 596.000 354.480 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 596.000 362.320 600.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END rst_n
  PIN sram_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 355.040 575.000 355.600 ;
    END
  END sram_addr[0]
  PIN sram_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 365.120 575.000 365.680 ;
    END
  END sram_addr[1]
  PIN sram_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 375.200 575.000 375.760 ;
    END
  END sram_addr[2]
  PIN sram_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 385.280 575.000 385.840 ;
    END
  END sram_addr[3]
  PIN sram_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 395.360 575.000 395.920 ;
    END
  END sram_addr[4]
  PIN sram_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 405.440 575.000 406.000 ;
    END
  END sram_addr[5]
  PIN sram_gwe
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 576.800 575.000 577.360 ;
    END
  END sram_gwe
  PIN sram_in[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 415.520 575.000 416.080 ;
    END
  END sram_in[0]
  PIN sram_in[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 425.600 575.000 426.160 ;
    END
  END sram_in[1]
  PIN sram_in[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 435.680 575.000 436.240 ;
    END
  END sram_in[2]
  PIN sram_in[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 445.760 575.000 446.320 ;
    END
  END sram_in[3]
  PIN sram_in[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 455.840 575.000 456.400 ;
    END
  END sram_in[4]
  PIN sram_in[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 465.920 575.000 466.480 ;
    END
  END sram_in[5]
  PIN sram_in[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 476.000 575.000 476.560 ;
    END
  END sram_in[6]
  PIN sram_in[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 486.080 575.000 486.640 ;
    END
  END sram_in[7]
  PIN sram_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 496.160 575.000 496.720 ;
    END
  END sram_out[0]
  PIN sram_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 506.240 575.000 506.800 ;
    END
  END sram_out[1]
  PIN sram_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 516.320 575.000 516.880 ;
    END
  END sram_out[2]
  PIN sram_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 526.400 575.000 526.960 ;
    END
  END sram_out[3]
  PIN sram_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 536.480 575.000 537.040 ;
    END
  END sram_out[4]
  PIN sram_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 546.560 575.000 547.120 ;
    END
  END sram_out[5]
  PIN sram_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 556.640 575.000 557.200 ;
    END
  END sram_out[6]
  PIN sram_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 571.000 566.720 575.000 567.280 ;
    END
  END sram_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.400 4.000 22.960 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 15.250 568.270 584.510 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 567.840 585.050 ;
      LAYER Metal2 ;
        RECT 0.140 595.700 32.180 596.820 ;
        RECT 33.340 595.700 40.020 596.820 ;
        RECT 41.180 595.700 47.860 596.820 ;
        RECT 49.020 595.700 55.700 596.820 ;
        RECT 56.860 595.700 63.540 596.820 ;
        RECT 64.700 595.700 71.380 596.820 ;
        RECT 72.540 595.700 79.220 596.820 ;
        RECT 80.380 595.700 87.060 596.820 ;
        RECT 88.220 595.700 94.900 596.820 ;
        RECT 96.060 595.700 102.740 596.820 ;
        RECT 103.900 595.700 110.580 596.820 ;
        RECT 111.740 595.700 118.420 596.820 ;
        RECT 119.580 595.700 126.260 596.820 ;
        RECT 127.420 595.700 134.100 596.820 ;
        RECT 135.260 595.700 141.940 596.820 ;
        RECT 143.100 595.700 149.780 596.820 ;
        RECT 150.940 595.700 157.620 596.820 ;
        RECT 158.780 595.700 165.460 596.820 ;
        RECT 166.620 595.700 173.300 596.820 ;
        RECT 174.460 595.700 181.140 596.820 ;
        RECT 182.300 595.700 188.980 596.820 ;
        RECT 190.140 595.700 196.820 596.820 ;
        RECT 197.980 595.700 204.660 596.820 ;
        RECT 205.820 595.700 212.500 596.820 ;
        RECT 213.660 595.700 220.340 596.820 ;
        RECT 221.500 595.700 228.180 596.820 ;
        RECT 229.340 595.700 236.020 596.820 ;
        RECT 237.180 595.700 243.860 596.820 ;
        RECT 245.020 595.700 251.700 596.820 ;
        RECT 252.860 595.700 259.540 596.820 ;
        RECT 260.700 595.700 267.380 596.820 ;
        RECT 268.540 595.700 275.220 596.820 ;
        RECT 276.380 595.700 283.060 596.820 ;
        RECT 284.220 595.700 290.900 596.820 ;
        RECT 292.060 595.700 298.740 596.820 ;
        RECT 299.900 595.700 306.580 596.820 ;
        RECT 307.740 595.700 314.420 596.820 ;
        RECT 315.580 595.700 322.260 596.820 ;
        RECT 323.420 595.700 330.100 596.820 ;
        RECT 331.260 595.700 337.940 596.820 ;
        RECT 339.100 595.700 345.780 596.820 ;
        RECT 346.940 595.700 353.620 596.820 ;
        RECT 354.780 595.700 361.460 596.820 ;
        RECT 362.620 595.700 369.300 596.820 ;
        RECT 370.460 595.700 377.140 596.820 ;
        RECT 378.300 595.700 384.980 596.820 ;
        RECT 386.140 595.700 392.820 596.820 ;
        RECT 393.980 595.700 400.660 596.820 ;
        RECT 401.820 595.700 408.500 596.820 ;
        RECT 409.660 595.700 416.340 596.820 ;
        RECT 417.500 595.700 424.180 596.820 ;
        RECT 425.340 595.700 432.020 596.820 ;
        RECT 433.180 595.700 439.860 596.820 ;
        RECT 441.020 595.700 447.700 596.820 ;
        RECT 448.860 595.700 455.540 596.820 ;
        RECT 456.700 595.700 463.380 596.820 ;
        RECT 464.540 595.700 471.220 596.820 ;
        RECT 472.380 595.700 479.060 596.820 ;
        RECT 480.220 595.700 486.900 596.820 ;
        RECT 488.060 595.700 494.740 596.820 ;
        RECT 495.900 595.700 502.580 596.820 ;
        RECT 503.740 595.700 510.420 596.820 ;
        RECT 511.580 595.700 518.260 596.820 ;
        RECT 519.420 595.700 526.100 596.820 ;
        RECT 527.260 595.700 533.940 596.820 ;
        RECT 535.100 595.700 541.780 596.820 ;
        RECT 542.940 595.700 567.700 596.820 ;
        RECT 0.140 15.490 567.700 595.700 ;
      LAYER Metal3 ;
        RECT 0.090 577.660 571.620 590.660 ;
        RECT 4.300 576.500 570.700 577.660 ;
        RECT 0.090 567.580 571.620 576.500 ;
        RECT 0.090 566.420 570.700 567.580 ;
        RECT 0.090 560.860 571.620 566.420 ;
        RECT 4.300 559.700 571.620 560.860 ;
        RECT 0.090 557.500 571.620 559.700 ;
        RECT 0.090 556.340 570.700 557.500 ;
        RECT 0.090 547.420 571.620 556.340 ;
        RECT 0.090 546.260 570.700 547.420 ;
        RECT 0.090 544.060 571.620 546.260 ;
        RECT 4.300 542.900 571.620 544.060 ;
        RECT 0.090 537.340 571.620 542.900 ;
        RECT 0.090 536.180 570.700 537.340 ;
        RECT 0.090 527.260 571.620 536.180 ;
        RECT 4.300 526.100 570.700 527.260 ;
        RECT 0.090 517.180 571.620 526.100 ;
        RECT 0.090 516.020 570.700 517.180 ;
        RECT 0.090 510.460 571.620 516.020 ;
        RECT 4.300 509.300 571.620 510.460 ;
        RECT 0.090 507.100 571.620 509.300 ;
        RECT 0.090 505.940 570.700 507.100 ;
        RECT 0.090 497.020 571.620 505.940 ;
        RECT 0.090 495.860 570.700 497.020 ;
        RECT 0.090 493.660 571.620 495.860 ;
        RECT 4.300 492.500 571.620 493.660 ;
        RECT 0.090 486.940 571.620 492.500 ;
        RECT 0.090 485.780 570.700 486.940 ;
        RECT 0.090 476.860 571.620 485.780 ;
        RECT 4.300 475.700 570.700 476.860 ;
        RECT 0.090 466.780 571.620 475.700 ;
        RECT 0.090 465.620 570.700 466.780 ;
        RECT 0.090 460.060 571.620 465.620 ;
        RECT 4.300 458.900 571.620 460.060 ;
        RECT 0.090 456.700 571.620 458.900 ;
        RECT 0.090 455.540 570.700 456.700 ;
        RECT 0.090 446.620 571.620 455.540 ;
        RECT 0.090 445.460 570.700 446.620 ;
        RECT 0.090 443.260 571.620 445.460 ;
        RECT 4.300 442.100 571.620 443.260 ;
        RECT 0.090 436.540 571.620 442.100 ;
        RECT 0.090 435.380 570.700 436.540 ;
        RECT 0.090 426.460 571.620 435.380 ;
        RECT 4.300 425.300 570.700 426.460 ;
        RECT 0.090 416.380 571.620 425.300 ;
        RECT 0.090 415.220 570.700 416.380 ;
        RECT 0.090 409.660 571.620 415.220 ;
        RECT 4.300 408.500 571.620 409.660 ;
        RECT 0.090 406.300 571.620 408.500 ;
        RECT 0.090 405.140 570.700 406.300 ;
        RECT 0.090 396.220 571.620 405.140 ;
        RECT 0.090 395.060 570.700 396.220 ;
        RECT 0.090 392.860 571.620 395.060 ;
        RECT 4.300 391.700 571.620 392.860 ;
        RECT 0.090 386.140 571.620 391.700 ;
        RECT 0.090 384.980 570.700 386.140 ;
        RECT 0.090 376.060 571.620 384.980 ;
        RECT 4.300 374.900 570.700 376.060 ;
        RECT 0.090 365.980 571.620 374.900 ;
        RECT 0.090 364.820 570.700 365.980 ;
        RECT 0.090 359.260 571.620 364.820 ;
        RECT 4.300 358.100 571.620 359.260 ;
        RECT 0.090 355.900 571.620 358.100 ;
        RECT 0.090 354.740 570.700 355.900 ;
        RECT 0.090 345.820 571.620 354.740 ;
        RECT 0.090 344.660 570.700 345.820 ;
        RECT 0.090 342.460 571.620 344.660 ;
        RECT 4.300 341.300 571.620 342.460 ;
        RECT 0.090 335.740 571.620 341.300 ;
        RECT 0.090 334.580 570.700 335.740 ;
        RECT 0.090 325.660 571.620 334.580 ;
        RECT 4.300 324.500 570.700 325.660 ;
        RECT 0.090 315.580 571.620 324.500 ;
        RECT 0.090 314.420 570.700 315.580 ;
        RECT 0.090 308.860 571.620 314.420 ;
        RECT 4.300 307.700 571.620 308.860 ;
        RECT 0.090 305.500 571.620 307.700 ;
        RECT 0.090 304.340 570.700 305.500 ;
        RECT 0.090 295.420 571.620 304.340 ;
        RECT 0.090 294.260 570.700 295.420 ;
        RECT 0.090 292.060 571.620 294.260 ;
        RECT 4.300 290.900 571.620 292.060 ;
        RECT 0.090 285.340 571.620 290.900 ;
        RECT 0.090 284.180 570.700 285.340 ;
        RECT 0.090 275.260 571.620 284.180 ;
        RECT 4.300 274.100 570.700 275.260 ;
        RECT 0.090 265.180 571.620 274.100 ;
        RECT 0.090 264.020 570.700 265.180 ;
        RECT 0.090 258.460 571.620 264.020 ;
        RECT 4.300 257.300 571.620 258.460 ;
        RECT 0.090 255.100 571.620 257.300 ;
        RECT 0.090 253.940 570.700 255.100 ;
        RECT 0.090 245.020 571.620 253.940 ;
        RECT 0.090 243.860 570.700 245.020 ;
        RECT 0.090 241.660 571.620 243.860 ;
        RECT 4.300 240.500 571.620 241.660 ;
        RECT 0.090 234.940 571.620 240.500 ;
        RECT 0.090 233.780 570.700 234.940 ;
        RECT 0.090 224.860 571.620 233.780 ;
        RECT 4.300 223.700 570.700 224.860 ;
        RECT 0.090 214.780 571.620 223.700 ;
        RECT 0.090 213.620 570.700 214.780 ;
        RECT 0.090 208.060 571.620 213.620 ;
        RECT 4.300 206.900 571.620 208.060 ;
        RECT 0.090 204.700 571.620 206.900 ;
        RECT 0.090 203.540 570.700 204.700 ;
        RECT 0.090 194.620 571.620 203.540 ;
        RECT 0.090 193.460 570.700 194.620 ;
        RECT 0.090 191.260 571.620 193.460 ;
        RECT 4.300 190.100 571.620 191.260 ;
        RECT 0.090 184.540 571.620 190.100 ;
        RECT 0.090 183.380 570.700 184.540 ;
        RECT 0.090 174.460 571.620 183.380 ;
        RECT 4.300 173.300 570.700 174.460 ;
        RECT 0.090 164.380 571.620 173.300 ;
        RECT 0.090 163.220 570.700 164.380 ;
        RECT 0.090 157.660 571.620 163.220 ;
        RECT 4.300 156.500 571.620 157.660 ;
        RECT 0.090 154.300 571.620 156.500 ;
        RECT 0.090 153.140 570.700 154.300 ;
        RECT 0.090 144.220 571.620 153.140 ;
        RECT 0.090 143.060 570.700 144.220 ;
        RECT 0.090 140.860 571.620 143.060 ;
        RECT 4.300 139.700 571.620 140.860 ;
        RECT 0.090 134.140 571.620 139.700 ;
        RECT 0.090 132.980 570.700 134.140 ;
        RECT 0.090 124.060 571.620 132.980 ;
        RECT 4.300 122.900 570.700 124.060 ;
        RECT 0.090 113.980 571.620 122.900 ;
        RECT 0.090 112.820 570.700 113.980 ;
        RECT 0.090 107.260 571.620 112.820 ;
        RECT 4.300 106.100 571.620 107.260 ;
        RECT 0.090 103.900 571.620 106.100 ;
        RECT 0.090 102.740 570.700 103.900 ;
        RECT 0.090 93.820 571.620 102.740 ;
        RECT 0.090 92.660 570.700 93.820 ;
        RECT 0.090 90.460 571.620 92.660 ;
        RECT 4.300 89.300 571.620 90.460 ;
        RECT 0.090 83.740 571.620 89.300 ;
        RECT 0.090 82.580 570.700 83.740 ;
        RECT 0.090 73.660 571.620 82.580 ;
        RECT 4.300 72.500 570.700 73.660 ;
        RECT 0.090 63.580 571.620 72.500 ;
        RECT 0.090 62.420 570.700 63.580 ;
        RECT 0.090 56.860 571.620 62.420 ;
        RECT 4.300 55.700 571.620 56.860 ;
        RECT 0.090 53.500 571.620 55.700 ;
        RECT 0.090 52.340 570.700 53.500 ;
        RECT 0.090 43.420 571.620 52.340 ;
        RECT 0.090 42.260 570.700 43.420 ;
        RECT 0.090 40.060 571.620 42.260 ;
        RECT 4.300 38.900 571.620 40.060 ;
        RECT 0.090 33.340 571.620 38.900 ;
        RECT 0.090 32.180 570.700 33.340 ;
        RECT 0.090 23.260 571.620 32.180 ;
        RECT 4.300 22.100 570.700 23.260 ;
        RECT 0.090 15.540 571.620 22.100 ;
      LAYER Metal4 ;
        RECT 42.700 584.680 562.660 588.470 ;
        RECT 42.700 80.730 98.740 584.680 ;
        RECT 100.940 80.730 175.540 584.680 ;
        RECT 177.740 80.730 252.340 584.680 ;
        RECT 254.540 80.730 329.140 584.680 ;
        RECT 331.340 80.730 405.940 584.680 ;
        RECT 408.140 80.730 482.740 584.680 ;
        RECT 484.940 80.730 559.540 584.680 ;
        RECT 561.740 80.730 562.660 584.680 ;
  END
END wrapped_qcpu
END LIBRARY

