magic
tech gf180mcuD
magscale 1 10
timestamp 1699956016
<< nwell >>
rect 1258 22304 24726 22822
rect 1258 21575 5789 21600
rect 1258 20761 24726 21575
rect 1258 20736 2989 20761
rect 1258 19193 24726 20032
rect 1258 19168 12087 19193
rect 1258 18439 2541 18464
rect 1258 17625 24726 18439
rect 1258 17600 6344 17625
rect 1258 16871 11837 16896
rect 1258 16057 24726 16871
rect 1258 16032 18109 16057
rect 1258 15303 10381 15328
rect 1258 14489 24726 15303
rect 1258 14464 8477 14489
rect 1258 13735 21133 13760
rect 1258 12921 24726 13735
rect 1258 12896 2541 12921
rect 1258 12167 2765 12192
rect 1258 11328 24726 12167
rect 1258 10599 5565 10624
rect 1258 9785 24726 10599
rect 1258 9760 2541 9785
rect 1258 9031 14456 9056
rect 1258 8217 24726 9031
rect 1258 8192 2541 8217
rect 1258 7463 15800 7488
rect 1258 6649 24726 7463
rect 1258 6624 17885 6649
rect 1258 5895 4109 5920
rect 1258 5081 24726 5895
rect 1258 5056 7805 5081
rect 1258 3488 24726 4352
<< pwell >>
rect 1258 21600 24726 22304
rect 1258 20032 24726 20736
rect 1258 18464 24726 19168
rect 1258 16896 24726 17600
rect 1258 15328 24726 16032
rect 1258 13760 24726 14464
rect 1258 12192 24726 12896
rect 1258 10624 24726 11328
rect 1258 9056 24726 9760
rect 1258 7488 24726 8192
rect 1258 5920 24726 6624
rect 1258 4352 24726 5056
rect 1258 3050 24726 3488
<< obsm1 >>
rect 1344 3076 24800 22796
<< metal2 >>
rect 4256 25200 4368 26000
rect 12768 25200 12880 26000
rect 21280 25200 21392 26000
<< obsm2 >>
rect 1820 25140 4196 25200
rect 4428 25140 12708 25200
rect 12940 25140 21220 25200
rect 21452 25140 24948 25200
rect 1820 1810 24948 25140
<< metal3 >>
rect 25200 23968 26000 24080
rect 25200 21952 26000 22064
rect 25200 19936 26000 20048
rect 25200 17920 26000 18032
rect 25200 15904 26000 16016
rect 25200 13888 26000 14000
rect 25200 11872 26000 11984
rect 25200 9856 26000 9968
rect 25200 7840 26000 7952
rect 25200 5824 26000 5936
rect 25200 3808 26000 3920
rect 25200 1792 26000 1904
<< obsm3 >>
rect 1810 23908 25140 24052
rect 1810 22124 25284 23908
rect 1810 21892 25140 22124
rect 1810 20108 25284 21892
rect 1810 19876 25140 20108
rect 1810 18092 25284 19876
rect 1810 17860 25140 18092
rect 1810 16076 25284 17860
rect 1810 15844 25140 16076
rect 1810 14060 25284 15844
rect 1810 13828 25140 14060
rect 1810 12044 25284 13828
rect 1810 11812 25140 12044
rect 1810 10028 25284 11812
rect 1810 9796 25140 10028
rect 1810 8012 25284 9796
rect 1810 7780 25140 8012
rect 1810 5996 25284 7780
rect 1810 5764 25140 5996
rect 1810 3980 25284 5764
rect 1810 3748 25140 3980
rect 1810 1964 25284 3748
rect 1810 1820 25140 1964
<< metal4 >>
rect 4096 3076 4416 22796
rect 7008 3076 7328 22796
rect 9920 3076 10240 22796
rect 12832 3076 13152 22796
rect 15744 3076 16064 22796
rect 18656 3076 18976 22796
rect 21568 3076 21888 22796
rect 24480 3076 24800 22796
<< obsm4 >>
rect 16604 7634 18596 20142
rect 19036 7634 21508 20142
rect 21948 7634 24276 20142
<< labels >>
rlabel metal3 s 25200 1792 26000 1904 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 25200 21952 26000 22064 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 25200 23968 26000 24080 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 25200 3808 26000 3920 6 custom_settings[1]
port 4 nsew signal input
rlabel metal3 s 25200 5824 26000 5936 6 custom_settings[2]
port 5 nsew signal input
rlabel metal3 s 25200 7840 26000 7952 6 custom_settings[3]
port 6 nsew signal input
rlabel metal3 s 25200 9856 26000 9968 6 custom_settings[4]
port 7 nsew signal input
rlabel metal3 s 25200 11872 26000 11984 6 custom_settings[5]
port 8 nsew signal input
rlabel metal3 s 25200 13888 26000 14000 6 custom_settings[6]
port 9 nsew signal input
rlabel metal3 s 25200 15904 26000 16016 6 custom_settings[7]
port 10 nsew signal input
rlabel metal3 s 25200 17920 26000 18032 6 custom_settings[8]
port 11 nsew signal input
rlabel metal3 s 25200 19936 26000 20048 6 custom_settings[9]
port 12 nsew signal input
rlabel metal2 s 21280 25200 21392 26000 6 io_out
port 13 nsew signal output
rlabel metal2 s 12768 25200 12880 26000 6 rst_n
port 14 nsew signal input
rlabel metal4 s 4096 3076 4416 22796 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 9920 3076 10240 22796 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 15744 3076 16064 22796 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 21568 3076 21888 22796 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 7008 3076 7328 22796 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 12832 3076 13152 22796 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 18656 3076 18976 22796 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 24480 3076 24800 22796 6 vss
port 16 nsew ground bidirectional
rlabel metal2 s 4256 25200 4368 26000 6 wb_clk_i
port 17 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 26000 26000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 581954
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/hellorld/runs/23_11_14_10_58/results/signoff/hellorld.magic.gds
string GDS_START 190832
<< end >>

