magic
tech gf180mcuD
magscale 1 5
timestamp 1698956690
<< obsm1 >>
rect 672 1415 59304 48369
<< metal2 >>
rect 2016 49600 2072 50000
rect 2688 49600 2744 50000
rect 3360 49600 3416 50000
rect 4032 49600 4088 50000
rect 4704 49600 4760 50000
rect 5376 49600 5432 50000
rect 6048 49600 6104 50000
rect 6720 49600 6776 50000
rect 7392 49600 7448 50000
rect 8064 49600 8120 50000
rect 8736 49600 8792 50000
rect 9408 49600 9464 50000
rect 10080 49600 10136 50000
rect 10752 49600 10808 50000
rect 11424 49600 11480 50000
rect 12096 49600 12152 50000
rect 12768 49600 12824 50000
rect 13440 49600 13496 50000
rect 14112 49600 14168 50000
rect 14784 49600 14840 50000
rect 15456 49600 15512 50000
rect 16128 49600 16184 50000
rect 16800 49600 16856 50000
rect 17472 49600 17528 50000
rect 18144 49600 18200 50000
rect 18816 49600 18872 50000
rect 19488 49600 19544 50000
rect 20160 49600 20216 50000
rect 20832 49600 20888 50000
rect 21504 49600 21560 50000
rect 22176 49600 22232 50000
rect 22848 49600 22904 50000
rect 23520 49600 23576 50000
rect 24192 49600 24248 50000
rect 24864 49600 24920 50000
rect 25536 49600 25592 50000
rect 26208 49600 26264 50000
rect 26880 49600 26936 50000
rect 27552 49600 27608 50000
rect 28224 49600 28280 50000
rect 28896 49600 28952 50000
rect 29568 49600 29624 50000
rect 30240 49600 30296 50000
rect 30912 49600 30968 50000
rect 31584 49600 31640 50000
rect 32256 49600 32312 50000
rect 32928 49600 32984 50000
rect 33600 49600 33656 50000
rect 34272 49600 34328 50000
rect 34944 49600 35000 50000
rect 35616 49600 35672 50000
rect 36288 49600 36344 50000
rect 36960 49600 37016 50000
rect 37632 49600 37688 50000
rect 38304 49600 38360 50000
rect 38976 49600 39032 50000
rect 39648 49600 39704 50000
rect 40320 49600 40376 50000
rect 40992 49600 41048 50000
rect 41664 49600 41720 50000
rect 42336 49600 42392 50000
rect 43008 49600 43064 50000
rect 43680 49600 43736 50000
rect 44352 49600 44408 50000
rect 45024 49600 45080 50000
rect 45696 49600 45752 50000
rect 46368 49600 46424 50000
rect 47040 49600 47096 50000
rect 47712 49600 47768 50000
rect 48384 49600 48440 50000
rect 49056 49600 49112 50000
rect 49728 49600 49784 50000
rect 50400 49600 50456 50000
rect 51072 49600 51128 50000
rect 51744 49600 51800 50000
rect 52416 49600 52472 50000
rect 53088 49600 53144 50000
rect 53760 49600 53816 50000
rect 54432 49600 54488 50000
rect 55104 49600 55160 50000
rect 55776 49600 55832 50000
rect 56448 49600 56504 50000
rect 57120 49600 57176 50000
rect 57792 49600 57848 50000
rect 112 0 168 400
rect 560 0 616 400
rect 1008 0 1064 400
rect 1456 0 1512 400
rect 1904 0 1960 400
rect 2352 0 2408 400
rect 2800 0 2856 400
rect 3248 0 3304 400
rect 3696 0 3752 400
rect 4144 0 4200 400
rect 4592 0 4648 400
rect 5040 0 5096 400
rect 5488 0 5544 400
rect 5936 0 5992 400
rect 6384 0 6440 400
rect 6832 0 6888 400
rect 7280 0 7336 400
rect 7728 0 7784 400
rect 8176 0 8232 400
rect 8624 0 8680 400
rect 9072 0 9128 400
rect 9520 0 9576 400
rect 9968 0 10024 400
rect 10416 0 10472 400
rect 10864 0 10920 400
rect 11312 0 11368 400
rect 11760 0 11816 400
rect 12208 0 12264 400
rect 12656 0 12712 400
rect 13104 0 13160 400
rect 13552 0 13608 400
rect 14000 0 14056 400
rect 14448 0 14504 400
rect 14896 0 14952 400
rect 15344 0 15400 400
rect 15792 0 15848 400
rect 16240 0 16296 400
rect 16688 0 16744 400
rect 17136 0 17192 400
rect 17584 0 17640 400
rect 18032 0 18088 400
rect 18480 0 18536 400
rect 18928 0 18984 400
rect 19376 0 19432 400
rect 19824 0 19880 400
rect 20272 0 20328 400
rect 20720 0 20776 400
rect 21168 0 21224 400
rect 21616 0 21672 400
rect 22064 0 22120 400
rect 22512 0 22568 400
rect 22960 0 23016 400
rect 23408 0 23464 400
rect 23856 0 23912 400
rect 24304 0 24360 400
rect 24752 0 24808 400
rect 25200 0 25256 400
rect 25648 0 25704 400
rect 26096 0 26152 400
rect 26544 0 26600 400
rect 26992 0 27048 400
rect 27440 0 27496 400
rect 27888 0 27944 400
rect 28336 0 28392 400
rect 28784 0 28840 400
rect 29232 0 29288 400
rect 29680 0 29736 400
rect 30128 0 30184 400
rect 30576 0 30632 400
rect 31024 0 31080 400
rect 31472 0 31528 400
rect 31920 0 31976 400
rect 32368 0 32424 400
rect 32816 0 32872 400
rect 33264 0 33320 400
rect 33712 0 33768 400
rect 34160 0 34216 400
rect 34608 0 34664 400
rect 35056 0 35112 400
rect 35504 0 35560 400
rect 35952 0 36008 400
rect 36400 0 36456 400
rect 36848 0 36904 400
rect 37296 0 37352 400
rect 37744 0 37800 400
rect 38192 0 38248 400
rect 38640 0 38696 400
rect 39088 0 39144 400
rect 39536 0 39592 400
rect 39984 0 40040 400
rect 40432 0 40488 400
rect 40880 0 40936 400
rect 41328 0 41384 400
rect 41776 0 41832 400
rect 42224 0 42280 400
rect 42672 0 42728 400
rect 43120 0 43176 400
rect 43568 0 43624 400
rect 44016 0 44072 400
rect 44464 0 44520 400
rect 44912 0 44968 400
rect 45360 0 45416 400
rect 45808 0 45864 400
rect 46256 0 46312 400
rect 46704 0 46760 400
rect 47152 0 47208 400
rect 47600 0 47656 400
rect 48048 0 48104 400
rect 48496 0 48552 400
rect 48944 0 49000 400
rect 49392 0 49448 400
rect 49840 0 49896 400
rect 50288 0 50344 400
rect 50736 0 50792 400
rect 51184 0 51240 400
rect 51632 0 51688 400
rect 52080 0 52136 400
rect 52528 0 52584 400
rect 52976 0 53032 400
rect 53424 0 53480 400
rect 53872 0 53928 400
rect 54320 0 54376 400
rect 54768 0 54824 400
rect 55216 0 55272 400
rect 55664 0 55720 400
rect 56112 0 56168 400
rect 56560 0 56616 400
rect 57008 0 57064 400
rect 57456 0 57512 400
rect 57904 0 57960 400
rect 58352 0 58408 400
rect 58800 0 58856 400
rect 59248 0 59304 400
rect 59696 0 59752 400
<< obsm2 >>
rect 126 49570 1986 49600
rect 2102 49570 2658 49600
rect 2774 49570 3330 49600
rect 3446 49570 4002 49600
rect 4118 49570 4674 49600
rect 4790 49570 5346 49600
rect 5462 49570 6018 49600
rect 6134 49570 6690 49600
rect 6806 49570 7362 49600
rect 7478 49570 8034 49600
rect 8150 49570 8706 49600
rect 8822 49570 9378 49600
rect 9494 49570 10050 49600
rect 10166 49570 10722 49600
rect 10838 49570 11394 49600
rect 11510 49570 12066 49600
rect 12182 49570 12738 49600
rect 12854 49570 13410 49600
rect 13526 49570 14082 49600
rect 14198 49570 14754 49600
rect 14870 49570 15426 49600
rect 15542 49570 16098 49600
rect 16214 49570 16770 49600
rect 16886 49570 17442 49600
rect 17558 49570 18114 49600
rect 18230 49570 18786 49600
rect 18902 49570 19458 49600
rect 19574 49570 20130 49600
rect 20246 49570 20802 49600
rect 20918 49570 21474 49600
rect 21590 49570 22146 49600
rect 22262 49570 22818 49600
rect 22934 49570 23490 49600
rect 23606 49570 24162 49600
rect 24278 49570 24834 49600
rect 24950 49570 25506 49600
rect 25622 49570 26178 49600
rect 26294 49570 26850 49600
rect 26966 49570 27522 49600
rect 27638 49570 28194 49600
rect 28310 49570 28866 49600
rect 28982 49570 29538 49600
rect 29654 49570 30210 49600
rect 30326 49570 30882 49600
rect 30998 49570 31554 49600
rect 31670 49570 32226 49600
rect 32342 49570 32898 49600
rect 33014 49570 33570 49600
rect 33686 49570 34242 49600
rect 34358 49570 34914 49600
rect 35030 49570 35586 49600
rect 35702 49570 36258 49600
rect 36374 49570 36930 49600
rect 37046 49570 37602 49600
rect 37718 49570 38274 49600
rect 38390 49570 38946 49600
rect 39062 49570 39618 49600
rect 39734 49570 40290 49600
rect 40406 49570 40962 49600
rect 41078 49570 41634 49600
rect 41750 49570 42306 49600
rect 42422 49570 42978 49600
rect 43094 49570 43650 49600
rect 43766 49570 44322 49600
rect 44438 49570 44994 49600
rect 45110 49570 45666 49600
rect 45782 49570 46338 49600
rect 46454 49570 47010 49600
rect 47126 49570 47682 49600
rect 47798 49570 48354 49600
rect 48470 49570 49026 49600
rect 49142 49570 49698 49600
rect 49814 49570 50370 49600
rect 50486 49570 51042 49600
rect 51158 49570 51714 49600
rect 51830 49570 52386 49600
rect 52502 49570 53058 49600
rect 53174 49570 53730 49600
rect 53846 49570 54402 49600
rect 54518 49570 55074 49600
rect 55190 49570 55746 49600
rect 55862 49570 56418 49600
rect 56534 49570 57090 49600
rect 57206 49570 57762 49600
rect 57878 49570 59738 49600
rect 126 430 59738 49570
rect 198 345 530 430
rect 646 345 978 430
rect 1094 345 1426 430
rect 1542 345 1874 430
rect 1990 345 2322 430
rect 2438 345 2770 430
rect 2886 345 3218 430
rect 3334 345 3666 430
rect 3782 345 4114 430
rect 4230 345 4562 430
rect 4678 345 5010 430
rect 5126 345 5458 430
rect 5574 345 5906 430
rect 6022 345 6354 430
rect 6470 345 6802 430
rect 6918 345 7250 430
rect 7366 345 7698 430
rect 7814 345 8146 430
rect 8262 345 8594 430
rect 8710 345 9042 430
rect 9158 345 9490 430
rect 9606 345 9938 430
rect 10054 345 10386 430
rect 10502 345 10834 430
rect 10950 345 11282 430
rect 11398 345 11730 430
rect 11846 345 12178 430
rect 12294 345 12626 430
rect 12742 345 13074 430
rect 13190 345 13522 430
rect 13638 345 13970 430
rect 14086 345 14418 430
rect 14534 345 14866 430
rect 14982 345 15314 430
rect 15430 345 15762 430
rect 15878 345 16210 430
rect 16326 345 16658 430
rect 16774 345 17106 430
rect 17222 345 17554 430
rect 17670 345 18002 430
rect 18118 345 18450 430
rect 18566 345 18898 430
rect 19014 345 19346 430
rect 19462 345 19794 430
rect 19910 345 20242 430
rect 20358 345 20690 430
rect 20806 345 21138 430
rect 21254 345 21586 430
rect 21702 345 22034 430
rect 22150 345 22482 430
rect 22598 345 22930 430
rect 23046 345 23378 430
rect 23494 345 23826 430
rect 23942 345 24274 430
rect 24390 345 24722 430
rect 24838 345 25170 430
rect 25286 345 25618 430
rect 25734 345 26066 430
rect 26182 345 26514 430
rect 26630 345 26962 430
rect 27078 345 27410 430
rect 27526 345 27858 430
rect 27974 345 28306 430
rect 28422 345 28754 430
rect 28870 345 29202 430
rect 29318 345 29650 430
rect 29766 345 30098 430
rect 30214 345 30546 430
rect 30662 345 30994 430
rect 31110 345 31442 430
rect 31558 345 31890 430
rect 32006 345 32338 430
rect 32454 345 32786 430
rect 32902 345 33234 430
rect 33350 345 33682 430
rect 33798 345 34130 430
rect 34246 345 34578 430
rect 34694 345 35026 430
rect 35142 345 35474 430
rect 35590 345 35922 430
rect 36038 345 36370 430
rect 36486 345 36818 430
rect 36934 345 37266 430
rect 37382 345 37714 430
rect 37830 345 38162 430
rect 38278 345 38610 430
rect 38726 345 39058 430
rect 39174 345 39506 430
rect 39622 345 39954 430
rect 40070 345 40402 430
rect 40518 345 40850 430
rect 40966 345 41298 430
rect 41414 345 41746 430
rect 41862 345 42194 430
rect 42310 345 42642 430
rect 42758 345 43090 430
rect 43206 345 43538 430
rect 43654 345 43986 430
rect 44102 345 44434 430
rect 44550 345 44882 430
rect 44998 345 45330 430
rect 45446 345 45778 430
rect 45894 345 46226 430
rect 46342 345 46674 430
rect 46790 345 47122 430
rect 47238 345 47570 430
rect 47686 345 48018 430
rect 48134 345 48466 430
rect 48582 345 48914 430
rect 49030 345 49362 430
rect 49478 345 49810 430
rect 49926 345 50258 430
rect 50374 345 50706 430
rect 50822 345 51154 430
rect 51270 345 51602 430
rect 51718 345 52050 430
rect 52166 345 52498 430
rect 52614 345 52946 430
rect 53062 345 53394 430
rect 53510 345 53842 430
rect 53958 345 54290 430
rect 54406 345 54738 430
rect 54854 345 55186 430
rect 55302 345 55634 430
rect 55750 345 56082 430
rect 56198 345 56530 430
rect 56646 345 56978 430
rect 57094 345 57426 430
rect 57542 345 57874 430
rect 57990 345 58322 430
rect 58438 345 58770 430
rect 58886 345 59218 430
rect 59334 345 59666 430
<< metal3 >>
rect 0 48832 400 48888
rect 0 48048 400 48104
rect 0 47264 400 47320
rect 0 46480 400 46536
rect 0 45696 400 45752
rect 0 44912 400 44968
rect 59600 44464 60000 44520
rect 0 44128 400 44184
rect 59600 44128 60000 44184
rect 59600 43792 60000 43848
rect 59600 43456 60000 43512
rect 0 43344 400 43400
rect 59600 43120 60000 43176
rect 59600 42784 60000 42840
rect 0 42560 400 42616
rect 59600 42448 60000 42504
rect 59600 42112 60000 42168
rect 0 41776 400 41832
rect 59600 41776 60000 41832
rect 59600 41440 60000 41496
rect 59600 41104 60000 41160
rect 0 40992 400 41048
rect 59600 40768 60000 40824
rect 59600 40432 60000 40488
rect 0 40208 400 40264
rect 59600 40096 60000 40152
rect 59600 39760 60000 39816
rect 0 39424 400 39480
rect 59600 39424 60000 39480
rect 59600 39088 60000 39144
rect 59600 38752 60000 38808
rect 0 38640 400 38696
rect 59600 38416 60000 38472
rect 59600 38080 60000 38136
rect 0 37856 400 37912
rect 59600 37744 60000 37800
rect 59600 37408 60000 37464
rect 0 37072 400 37128
rect 59600 37072 60000 37128
rect 59600 36736 60000 36792
rect 59600 36400 60000 36456
rect 0 36288 400 36344
rect 59600 36064 60000 36120
rect 59600 35728 60000 35784
rect 0 35504 400 35560
rect 59600 35392 60000 35448
rect 59600 35056 60000 35112
rect 0 34720 400 34776
rect 59600 34720 60000 34776
rect 59600 34384 60000 34440
rect 59600 34048 60000 34104
rect 0 33936 400 33992
rect 59600 33712 60000 33768
rect 59600 33376 60000 33432
rect 0 33152 400 33208
rect 59600 33040 60000 33096
rect 59600 32704 60000 32760
rect 0 32368 400 32424
rect 59600 32368 60000 32424
rect 59600 32032 60000 32088
rect 59600 31696 60000 31752
rect 0 31584 400 31640
rect 59600 31360 60000 31416
rect 59600 31024 60000 31080
rect 0 30800 400 30856
rect 59600 30688 60000 30744
rect 59600 30352 60000 30408
rect 0 30016 400 30072
rect 59600 30016 60000 30072
rect 59600 29680 60000 29736
rect 59600 29344 60000 29400
rect 0 29232 400 29288
rect 59600 29008 60000 29064
rect 59600 28672 60000 28728
rect 0 28448 400 28504
rect 59600 28336 60000 28392
rect 59600 28000 60000 28056
rect 0 27664 400 27720
rect 59600 27664 60000 27720
rect 59600 27328 60000 27384
rect 59600 26992 60000 27048
rect 0 26880 400 26936
rect 59600 26656 60000 26712
rect 59600 26320 60000 26376
rect 0 26096 400 26152
rect 59600 25984 60000 26040
rect 59600 25648 60000 25704
rect 0 25312 400 25368
rect 59600 25312 60000 25368
rect 59600 24976 60000 25032
rect 59600 24640 60000 24696
rect 0 24528 400 24584
rect 59600 24304 60000 24360
rect 59600 23968 60000 24024
rect 0 23744 400 23800
rect 59600 23632 60000 23688
rect 59600 23296 60000 23352
rect 0 22960 400 23016
rect 59600 22960 60000 23016
rect 59600 22624 60000 22680
rect 59600 22288 60000 22344
rect 0 22176 400 22232
rect 59600 21952 60000 22008
rect 59600 21616 60000 21672
rect 0 21392 400 21448
rect 59600 21280 60000 21336
rect 59600 20944 60000 21000
rect 0 20608 400 20664
rect 59600 20608 60000 20664
rect 59600 20272 60000 20328
rect 59600 19936 60000 19992
rect 0 19824 400 19880
rect 59600 19600 60000 19656
rect 59600 19264 60000 19320
rect 0 19040 400 19096
rect 59600 18928 60000 18984
rect 59600 18592 60000 18648
rect 0 18256 400 18312
rect 59600 18256 60000 18312
rect 59600 17920 60000 17976
rect 59600 17584 60000 17640
rect 0 17472 400 17528
rect 59600 17248 60000 17304
rect 59600 16912 60000 16968
rect 0 16688 400 16744
rect 59600 16576 60000 16632
rect 59600 16240 60000 16296
rect 0 15904 400 15960
rect 59600 15904 60000 15960
rect 59600 15568 60000 15624
rect 59600 15232 60000 15288
rect 0 15120 400 15176
rect 59600 14896 60000 14952
rect 59600 14560 60000 14616
rect 0 14336 400 14392
rect 59600 14224 60000 14280
rect 59600 13888 60000 13944
rect 0 13552 400 13608
rect 59600 13552 60000 13608
rect 59600 13216 60000 13272
rect 59600 12880 60000 12936
rect 0 12768 400 12824
rect 59600 12544 60000 12600
rect 59600 12208 60000 12264
rect 0 11984 400 12040
rect 59600 11872 60000 11928
rect 59600 11536 60000 11592
rect 0 11200 400 11256
rect 59600 11200 60000 11256
rect 59600 10864 60000 10920
rect 59600 10528 60000 10584
rect 0 10416 400 10472
rect 59600 10192 60000 10248
rect 59600 9856 60000 9912
rect 0 9632 400 9688
rect 59600 9520 60000 9576
rect 59600 9184 60000 9240
rect 0 8848 400 8904
rect 59600 8848 60000 8904
rect 59600 8512 60000 8568
rect 59600 8176 60000 8232
rect 0 8064 400 8120
rect 59600 7840 60000 7896
rect 59600 7504 60000 7560
rect 0 7280 400 7336
rect 59600 7168 60000 7224
rect 59600 6832 60000 6888
rect 0 6496 400 6552
rect 59600 6496 60000 6552
rect 59600 6160 60000 6216
rect 59600 5824 60000 5880
rect 0 5712 400 5768
rect 59600 5488 60000 5544
rect 0 4928 400 4984
rect 0 4144 400 4200
rect 0 3360 400 3416
rect 0 2576 400 2632
rect 0 1792 400 1848
rect 0 1008 400 1064
<< obsm3 >>
rect 430 48802 59743 48874
rect 121 48134 59743 48802
rect 430 48018 59743 48134
rect 121 47350 59743 48018
rect 430 47234 59743 47350
rect 121 46566 59743 47234
rect 430 46450 59743 46566
rect 121 45782 59743 46450
rect 430 45666 59743 45782
rect 121 44998 59743 45666
rect 430 44882 59743 44998
rect 121 44550 59743 44882
rect 121 44434 59570 44550
rect 121 44214 59743 44434
rect 430 44098 59570 44214
rect 121 43878 59743 44098
rect 121 43762 59570 43878
rect 121 43542 59743 43762
rect 121 43430 59570 43542
rect 430 43426 59570 43430
rect 430 43314 59743 43426
rect 121 43206 59743 43314
rect 121 43090 59570 43206
rect 121 42870 59743 43090
rect 121 42754 59570 42870
rect 121 42646 59743 42754
rect 430 42534 59743 42646
rect 430 42530 59570 42534
rect 121 42418 59570 42530
rect 121 42198 59743 42418
rect 121 42082 59570 42198
rect 121 41862 59743 42082
rect 430 41746 59570 41862
rect 121 41526 59743 41746
rect 121 41410 59570 41526
rect 121 41190 59743 41410
rect 121 41078 59570 41190
rect 430 41074 59570 41078
rect 430 40962 59743 41074
rect 121 40854 59743 40962
rect 121 40738 59570 40854
rect 121 40518 59743 40738
rect 121 40402 59570 40518
rect 121 40294 59743 40402
rect 430 40182 59743 40294
rect 430 40178 59570 40182
rect 121 40066 59570 40178
rect 121 39846 59743 40066
rect 121 39730 59570 39846
rect 121 39510 59743 39730
rect 430 39394 59570 39510
rect 121 39174 59743 39394
rect 121 39058 59570 39174
rect 121 38838 59743 39058
rect 121 38726 59570 38838
rect 430 38722 59570 38726
rect 430 38610 59743 38722
rect 121 38502 59743 38610
rect 121 38386 59570 38502
rect 121 38166 59743 38386
rect 121 38050 59570 38166
rect 121 37942 59743 38050
rect 430 37830 59743 37942
rect 430 37826 59570 37830
rect 121 37714 59570 37826
rect 121 37494 59743 37714
rect 121 37378 59570 37494
rect 121 37158 59743 37378
rect 430 37042 59570 37158
rect 121 36822 59743 37042
rect 121 36706 59570 36822
rect 121 36486 59743 36706
rect 121 36374 59570 36486
rect 430 36370 59570 36374
rect 430 36258 59743 36370
rect 121 36150 59743 36258
rect 121 36034 59570 36150
rect 121 35814 59743 36034
rect 121 35698 59570 35814
rect 121 35590 59743 35698
rect 430 35478 59743 35590
rect 430 35474 59570 35478
rect 121 35362 59570 35474
rect 121 35142 59743 35362
rect 121 35026 59570 35142
rect 121 34806 59743 35026
rect 430 34690 59570 34806
rect 121 34470 59743 34690
rect 121 34354 59570 34470
rect 121 34134 59743 34354
rect 121 34022 59570 34134
rect 430 34018 59570 34022
rect 430 33906 59743 34018
rect 121 33798 59743 33906
rect 121 33682 59570 33798
rect 121 33462 59743 33682
rect 121 33346 59570 33462
rect 121 33238 59743 33346
rect 430 33126 59743 33238
rect 430 33122 59570 33126
rect 121 33010 59570 33122
rect 121 32790 59743 33010
rect 121 32674 59570 32790
rect 121 32454 59743 32674
rect 430 32338 59570 32454
rect 121 32118 59743 32338
rect 121 32002 59570 32118
rect 121 31782 59743 32002
rect 121 31670 59570 31782
rect 430 31666 59570 31670
rect 430 31554 59743 31666
rect 121 31446 59743 31554
rect 121 31330 59570 31446
rect 121 31110 59743 31330
rect 121 30994 59570 31110
rect 121 30886 59743 30994
rect 430 30774 59743 30886
rect 430 30770 59570 30774
rect 121 30658 59570 30770
rect 121 30438 59743 30658
rect 121 30322 59570 30438
rect 121 30102 59743 30322
rect 430 29986 59570 30102
rect 121 29766 59743 29986
rect 121 29650 59570 29766
rect 121 29430 59743 29650
rect 121 29318 59570 29430
rect 430 29314 59570 29318
rect 430 29202 59743 29314
rect 121 29094 59743 29202
rect 121 28978 59570 29094
rect 121 28758 59743 28978
rect 121 28642 59570 28758
rect 121 28534 59743 28642
rect 430 28422 59743 28534
rect 430 28418 59570 28422
rect 121 28306 59570 28418
rect 121 28086 59743 28306
rect 121 27970 59570 28086
rect 121 27750 59743 27970
rect 430 27634 59570 27750
rect 121 27414 59743 27634
rect 121 27298 59570 27414
rect 121 27078 59743 27298
rect 121 26966 59570 27078
rect 430 26962 59570 26966
rect 430 26850 59743 26962
rect 121 26742 59743 26850
rect 121 26626 59570 26742
rect 121 26406 59743 26626
rect 121 26290 59570 26406
rect 121 26182 59743 26290
rect 430 26070 59743 26182
rect 430 26066 59570 26070
rect 121 25954 59570 26066
rect 121 25734 59743 25954
rect 121 25618 59570 25734
rect 121 25398 59743 25618
rect 430 25282 59570 25398
rect 121 25062 59743 25282
rect 121 24946 59570 25062
rect 121 24726 59743 24946
rect 121 24614 59570 24726
rect 430 24610 59570 24614
rect 430 24498 59743 24610
rect 121 24390 59743 24498
rect 121 24274 59570 24390
rect 121 24054 59743 24274
rect 121 23938 59570 24054
rect 121 23830 59743 23938
rect 430 23718 59743 23830
rect 430 23714 59570 23718
rect 121 23602 59570 23714
rect 121 23382 59743 23602
rect 121 23266 59570 23382
rect 121 23046 59743 23266
rect 430 22930 59570 23046
rect 121 22710 59743 22930
rect 121 22594 59570 22710
rect 121 22374 59743 22594
rect 121 22262 59570 22374
rect 430 22258 59570 22262
rect 430 22146 59743 22258
rect 121 22038 59743 22146
rect 121 21922 59570 22038
rect 121 21702 59743 21922
rect 121 21586 59570 21702
rect 121 21478 59743 21586
rect 430 21366 59743 21478
rect 430 21362 59570 21366
rect 121 21250 59570 21362
rect 121 21030 59743 21250
rect 121 20914 59570 21030
rect 121 20694 59743 20914
rect 430 20578 59570 20694
rect 121 20358 59743 20578
rect 121 20242 59570 20358
rect 121 20022 59743 20242
rect 121 19910 59570 20022
rect 430 19906 59570 19910
rect 430 19794 59743 19906
rect 121 19686 59743 19794
rect 121 19570 59570 19686
rect 121 19350 59743 19570
rect 121 19234 59570 19350
rect 121 19126 59743 19234
rect 430 19014 59743 19126
rect 430 19010 59570 19014
rect 121 18898 59570 19010
rect 121 18678 59743 18898
rect 121 18562 59570 18678
rect 121 18342 59743 18562
rect 430 18226 59570 18342
rect 121 18006 59743 18226
rect 121 17890 59570 18006
rect 121 17670 59743 17890
rect 121 17558 59570 17670
rect 430 17554 59570 17558
rect 430 17442 59743 17554
rect 121 17334 59743 17442
rect 121 17218 59570 17334
rect 121 16998 59743 17218
rect 121 16882 59570 16998
rect 121 16774 59743 16882
rect 430 16662 59743 16774
rect 430 16658 59570 16662
rect 121 16546 59570 16658
rect 121 16326 59743 16546
rect 121 16210 59570 16326
rect 121 15990 59743 16210
rect 430 15874 59570 15990
rect 121 15654 59743 15874
rect 121 15538 59570 15654
rect 121 15318 59743 15538
rect 121 15206 59570 15318
rect 430 15202 59570 15206
rect 430 15090 59743 15202
rect 121 14982 59743 15090
rect 121 14866 59570 14982
rect 121 14646 59743 14866
rect 121 14530 59570 14646
rect 121 14422 59743 14530
rect 430 14310 59743 14422
rect 430 14306 59570 14310
rect 121 14194 59570 14306
rect 121 13974 59743 14194
rect 121 13858 59570 13974
rect 121 13638 59743 13858
rect 430 13522 59570 13638
rect 121 13302 59743 13522
rect 121 13186 59570 13302
rect 121 12966 59743 13186
rect 121 12854 59570 12966
rect 430 12850 59570 12854
rect 430 12738 59743 12850
rect 121 12630 59743 12738
rect 121 12514 59570 12630
rect 121 12294 59743 12514
rect 121 12178 59570 12294
rect 121 12070 59743 12178
rect 430 11958 59743 12070
rect 430 11954 59570 11958
rect 121 11842 59570 11954
rect 121 11622 59743 11842
rect 121 11506 59570 11622
rect 121 11286 59743 11506
rect 430 11170 59570 11286
rect 121 10950 59743 11170
rect 121 10834 59570 10950
rect 121 10614 59743 10834
rect 121 10502 59570 10614
rect 430 10498 59570 10502
rect 430 10386 59743 10498
rect 121 10278 59743 10386
rect 121 10162 59570 10278
rect 121 9942 59743 10162
rect 121 9826 59570 9942
rect 121 9718 59743 9826
rect 430 9606 59743 9718
rect 430 9602 59570 9606
rect 121 9490 59570 9602
rect 121 9270 59743 9490
rect 121 9154 59570 9270
rect 121 8934 59743 9154
rect 430 8818 59570 8934
rect 121 8598 59743 8818
rect 121 8482 59570 8598
rect 121 8262 59743 8482
rect 121 8150 59570 8262
rect 430 8146 59570 8150
rect 430 8034 59743 8146
rect 121 7926 59743 8034
rect 121 7810 59570 7926
rect 121 7590 59743 7810
rect 121 7474 59570 7590
rect 121 7366 59743 7474
rect 430 7254 59743 7366
rect 430 7250 59570 7254
rect 121 7138 59570 7250
rect 121 6918 59743 7138
rect 121 6802 59570 6918
rect 121 6582 59743 6802
rect 430 6466 59570 6582
rect 121 6246 59743 6466
rect 121 6130 59570 6246
rect 121 5910 59743 6130
rect 121 5798 59570 5910
rect 430 5794 59570 5798
rect 430 5682 59743 5794
rect 121 5574 59743 5682
rect 121 5458 59570 5574
rect 121 5014 59743 5458
rect 430 4898 59743 5014
rect 121 4230 59743 4898
rect 430 4114 59743 4230
rect 121 3446 59743 4114
rect 430 3330 59743 3446
rect 121 2662 59743 3330
rect 430 2546 59743 2662
rect 121 1878 59743 2546
rect 430 1762 59743 1878
rect 121 1094 59743 1762
rect 430 978 59743 1094
rect 121 350 59743 978
<< metal4 >>
rect 2224 1538 2384 48246
rect 9904 1538 10064 48246
rect 17584 1538 17744 48246
rect 25264 1538 25424 48246
rect 32944 1538 33104 48246
rect 40624 1538 40784 48246
rect 48304 1538 48464 48246
rect 55984 1538 56144 48246
<< obsm4 >>
rect 7182 1508 9874 47871
rect 10094 1508 17554 47871
rect 17774 1508 25234 47871
rect 25454 1508 32914 47871
rect 33134 1508 40594 47871
rect 40814 1508 48274 47871
rect 48494 1508 55954 47871
rect 56174 1508 59178 47871
rect 7182 1241 59178 1508
<< labels >>
rlabel metal2 s 55776 49600 55832 50000 6 blinker_do[0]
port 1 nsew signal input
rlabel metal2 s 56448 49600 56504 50000 6 blinker_do[1]
port 2 nsew signal input
rlabel metal2 s 57120 49600 57176 50000 6 blinker_do[2]
port 3 nsew signal input
rlabel metal3 s 59600 17584 60000 17640 6 custom_settings[0]
port 4 nsew signal output
rlabel metal3 s 59600 20944 60000 21000 6 custom_settings[10]
port 5 nsew signal output
rlabel metal3 s 59600 21280 60000 21336 6 custom_settings[11]
port 6 nsew signal output
rlabel metal3 s 59600 21616 60000 21672 6 custom_settings[12]
port 7 nsew signal output
rlabel metal3 s 59600 21952 60000 22008 6 custom_settings[13]
port 8 nsew signal output
rlabel metal3 s 59600 22288 60000 22344 6 custom_settings[14]
port 9 nsew signal output
rlabel metal3 s 59600 22624 60000 22680 6 custom_settings[15]
port 10 nsew signal output
rlabel metal3 s 59600 22960 60000 23016 6 custom_settings[16]
port 11 nsew signal output
rlabel metal3 s 59600 23296 60000 23352 6 custom_settings[17]
port 12 nsew signal output
rlabel metal3 s 59600 23632 60000 23688 6 custom_settings[18]
port 13 nsew signal output
rlabel metal3 s 59600 23968 60000 24024 6 custom_settings[19]
port 14 nsew signal output
rlabel metal3 s 59600 17920 60000 17976 6 custom_settings[1]
port 15 nsew signal output
rlabel metal3 s 59600 24304 60000 24360 6 custom_settings[20]
port 16 nsew signal output
rlabel metal3 s 59600 24640 60000 24696 6 custom_settings[21]
port 17 nsew signal output
rlabel metal3 s 59600 24976 60000 25032 6 custom_settings[22]
port 18 nsew signal output
rlabel metal3 s 59600 25312 60000 25368 6 custom_settings[23]
port 19 nsew signal output
rlabel metal3 s 59600 25648 60000 25704 6 custom_settings[24]
port 20 nsew signal output
rlabel metal3 s 59600 25984 60000 26040 6 custom_settings[25]
port 21 nsew signal output
rlabel metal3 s 59600 26320 60000 26376 6 custom_settings[26]
port 22 nsew signal output
rlabel metal3 s 59600 26656 60000 26712 6 custom_settings[27]
port 23 nsew signal output
rlabel metal3 s 59600 26992 60000 27048 6 custom_settings[28]
port 24 nsew signal output
rlabel metal3 s 59600 27328 60000 27384 6 custom_settings[29]
port 25 nsew signal output
rlabel metal3 s 59600 18256 60000 18312 6 custom_settings[2]
port 26 nsew signal output
rlabel metal3 s 59600 27664 60000 27720 6 custom_settings[30]
port 27 nsew signal output
rlabel metal3 s 59600 28000 60000 28056 6 custom_settings[31]
port 28 nsew signal output
rlabel metal3 s 59600 18592 60000 18648 6 custom_settings[3]
port 29 nsew signal output
rlabel metal3 s 59600 18928 60000 18984 6 custom_settings[4]
port 30 nsew signal output
rlabel metal3 s 59600 19264 60000 19320 6 custom_settings[5]
port 31 nsew signal output
rlabel metal3 s 59600 19600 60000 19656 6 custom_settings[6]
port 32 nsew signal output
rlabel metal3 s 59600 19936 60000 19992 6 custom_settings[7]
port 33 nsew signal output
rlabel metal3 s 59600 20272 60000 20328 6 custom_settings[8]
port 34 nsew signal output
rlabel metal3 s 59600 20608 60000 20664 6 custom_settings[9]
port 35 nsew signal output
rlabel metal2 s 2016 49600 2072 50000 6 io_in[0]
port 36 nsew signal input
rlabel metal2 s 8736 49600 8792 50000 6 io_in[10]
port 37 nsew signal input
rlabel metal2 s 9408 49600 9464 50000 6 io_in[11]
port 38 nsew signal input
rlabel metal2 s 10080 49600 10136 50000 6 io_in[12]
port 39 nsew signal input
rlabel metal2 s 10752 49600 10808 50000 6 io_in[13]
port 40 nsew signal input
rlabel metal2 s 11424 49600 11480 50000 6 io_in[14]
port 41 nsew signal input
rlabel metal2 s 12096 49600 12152 50000 6 io_in[15]
port 42 nsew signal input
rlabel metal2 s 12768 49600 12824 50000 6 io_in[16]
port 43 nsew signal input
rlabel metal2 s 13440 49600 13496 50000 6 io_in[17]
port 44 nsew signal input
rlabel metal2 s 14112 49600 14168 50000 6 io_in[18]
port 45 nsew signal input
rlabel metal2 s 14784 49600 14840 50000 6 io_in[19]
port 46 nsew signal input
rlabel metal2 s 2688 49600 2744 50000 6 io_in[1]
port 47 nsew signal input
rlabel metal2 s 15456 49600 15512 50000 6 io_in[20]
port 48 nsew signal input
rlabel metal2 s 16128 49600 16184 50000 6 io_in[21]
port 49 nsew signal input
rlabel metal2 s 16800 49600 16856 50000 6 io_in[22]
port 50 nsew signal input
rlabel metal2 s 17472 49600 17528 50000 6 io_in[23]
port 51 nsew signal input
rlabel metal2 s 18144 49600 18200 50000 6 io_in[24]
port 52 nsew signal input
rlabel metal2 s 18816 49600 18872 50000 6 io_in[25]
port 53 nsew signal input
rlabel metal2 s 19488 49600 19544 50000 6 io_in[26]
port 54 nsew signal input
rlabel metal2 s 20160 49600 20216 50000 6 io_in[27]
port 55 nsew signal input
rlabel metal2 s 20832 49600 20888 50000 6 io_in[28]
port 56 nsew signal input
rlabel metal2 s 21504 49600 21560 50000 6 io_in[29]
port 57 nsew signal input
rlabel metal2 s 3360 49600 3416 50000 6 io_in[2]
port 58 nsew signal input
rlabel metal2 s 22176 49600 22232 50000 6 io_in[30]
port 59 nsew signal input
rlabel metal2 s 22848 49600 22904 50000 6 io_in[31]
port 60 nsew signal input
rlabel metal2 s 23520 49600 23576 50000 6 io_in[32]
port 61 nsew signal input
rlabel metal2 s 24192 49600 24248 50000 6 io_in[33]
port 62 nsew signal input
rlabel metal2 s 24864 49600 24920 50000 6 io_in[34]
port 63 nsew signal input
rlabel metal2 s 25536 49600 25592 50000 6 io_in[35]
port 64 nsew signal input
rlabel metal2 s 26208 49600 26264 50000 6 io_in[36]
port 65 nsew signal input
rlabel metal2 s 26880 49600 26936 50000 6 io_in[37]
port 66 nsew signal input
rlabel metal2 s 4032 49600 4088 50000 6 io_in[3]
port 67 nsew signal input
rlabel metal2 s 4704 49600 4760 50000 6 io_in[4]
port 68 nsew signal input
rlabel metal2 s 5376 49600 5432 50000 6 io_in[5]
port 69 nsew signal input
rlabel metal2 s 6048 49600 6104 50000 6 io_in[6]
port 70 nsew signal input
rlabel metal2 s 6720 49600 6776 50000 6 io_in[7]
port 71 nsew signal input
rlabel metal2 s 7392 49600 7448 50000 6 io_in[8]
port 72 nsew signal input
rlabel metal2 s 8064 49600 8120 50000 6 io_in[9]
port 73 nsew signal input
rlabel metal3 s 0 1008 400 1064 6 io_oeb[0]
port 74 nsew signal output
rlabel metal3 s 0 8848 400 8904 6 io_oeb[10]
port 75 nsew signal output
rlabel metal3 s 0 9632 400 9688 6 io_oeb[11]
port 76 nsew signal output
rlabel metal3 s 0 10416 400 10472 6 io_oeb[12]
port 77 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 io_oeb[13]
port 78 nsew signal output
rlabel metal3 s 0 11984 400 12040 6 io_oeb[14]
port 79 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 io_oeb[15]
port 80 nsew signal output
rlabel metal3 s 0 13552 400 13608 6 io_oeb[16]
port 81 nsew signal output
rlabel metal3 s 0 14336 400 14392 6 io_oeb[17]
port 82 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 io_oeb[18]
port 83 nsew signal output
rlabel metal3 s 0 15904 400 15960 6 io_oeb[19]
port 84 nsew signal output
rlabel metal3 s 0 1792 400 1848 6 io_oeb[1]
port 85 nsew signal output
rlabel metal3 s 0 16688 400 16744 6 io_oeb[20]
port 86 nsew signal output
rlabel metal3 s 0 17472 400 17528 6 io_oeb[21]
port 87 nsew signal output
rlabel metal3 s 0 18256 400 18312 6 io_oeb[22]
port 88 nsew signal output
rlabel metal3 s 0 19040 400 19096 6 io_oeb[23]
port 89 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 io_oeb[24]
port 90 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 io_oeb[25]
port 91 nsew signal output
rlabel metal3 s 0 21392 400 21448 6 io_oeb[26]
port 92 nsew signal output
rlabel metal3 s 0 22176 400 22232 6 io_oeb[27]
port 93 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 io_oeb[28]
port 94 nsew signal output
rlabel metal3 s 0 23744 400 23800 6 io_oeb[29]
port 95 nsew signal output
rlabel metal3 s 0 2576 400 2632 6 io_oeb[2]
port 96 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 io_oeb[30]
port 97 nsew signal output
rlabel metal3 s 0 25312 400 25368 6 io_oeb[31]
port 98 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 io_oeb[32]
port 99 nsew signal output
rlabel metal3 s 0 26880 400 26936 6 io_oeb[33]
port 100 nsew signal output
rlabel metal3 s 0 27664 400 27720 6 io_oeb[34]
port 101 nsew signal output
rlabel metal3 s 0 28448 400 28504 6 io_oeb[35]
port 102 nsew signal output
rlabel metal3 s 0 29232 400 29288 6 io_oeb[36]
port 103 nsew signal output
rlabel metal3 s 0 30016 400 30072 6 io_oeb[37]
port 104 nsew signal output
rlabel metal3 s 0 3360 400 3416 6 io_oeb[3]
port 105 nsew signal output
rlabel metal3 s 0 4144 400 4200 6 io_oeb[4]
port 106 nsew signal output
rlabel metal3 s 0 4928 400 4984 6 io_oeb[5]
port 107 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 io_oeb[6]
port 108 nsew signal output
rlabel metal3 s 0 6496 400 6552 6 io_oeb[7]
port 109 nsew signal output
rlabel metal3 s 0 7280 400 7336 6 io_oeb[8]
port 110 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 io_oeb[9]
port 111 nsew signal output
rlabel metal2 s 27552 49600 27608 50000 6 io_out[0]
port 112 nsew signal output
rlabel metal2 s 34272 49600 34328 50000 6 io_out[10]
port 113 nsew signal output
rlabel metal2 s 34944 49600 35000 50000 6 io_out[11]
port 114 nsew signal output
rlabel metal2 s 35616 49600 35672 50000 6 io_out[12]
port 115 nsew signal output
rlabel metal2 s 36288 49600 36344 50000 6 io_out[13]
port 116 nsew signal output
rlabel metal2 s 36960 49600 37016 50000 6 io_out[14]
port 117 nsew signal output
rlabel metal2 s 37632 49600 37688 50000 6 io_out[15]
port 118 nsew signal output
rlabel metal2 s 38304 49600 38360 50000 6 io_out[16]
port 119 nsew signal output
rlabel metal2 s 38976 49600 39032 50000 6 io_out[17]
port 120 nsew signal output
rlabel metal2 s 39648 49600 39704 50000 6 io_out[18]
port 121 nsew signal output
rlabel metal2 s 40320 49600 40376 50000 6 io_out[19]
port 122 nsew signal output
rlabel metal2 s 28224 49600 28280 50000 6 io_out[1]
port 123 nsew signal output
rlabel metal2 s 40992 49600 41048 50000 6 io_out[20]
port 124 nsew signal output
rlabel metal2 s 41664 49600 41720 50000 6 io_out[21]
port 125 nsew signal output
rlabel metal2 s 42336 49600 42392 50000 6 io_out[22]
port 126 nsew signal output
rlabel metal2 s 43008 49600 43064 50000 6 io_out[23]
port 127 nsew signal output
rlabel metal2 s 43680 49600 43736 50000 6 io_out[24]
port 128 nsew signal output
rlabel metal2 s 44352 49600 44408 50000 6 io_out[25]
port 129 nsew signal output
rlabel metal2 s 45024 49600 45080 50000 6 io_out[26]
port 130 nsew signal output
rlabel metal2 s 45696 49600 45752 50000 6 io_out[27]
port 131 nsew signal output
rlabel metal2 s 46368 49600 46424 50000 6 io_out[28]
port 132 nsew signal output
rlabel metal2 s 47040 49600 47096 50000 6 io_out[29]
port 133 nsew signal output
rlabel metal2 s 28896 49600 28952 50000 6 io_out[2]
port 134 nsew signal output
rlabel metal2 s 47712 49600 47768 50000 6 io_out[30]
port 135 nsew signal output
rlabel metal2 s 48384 49600 48440 50000 6 io_out[31]
port 136 nsew signal output
rlabel metal2 s 49056 49600 49112 50000 6 io_out[32]
port 137 nsew signal output
rlabel metal2 s 49728 49600 49784 50000 6 io_out[33]
port 138 nsew signal output
rlabel metal2 s 50400 49600 50456 50000 6 io_out[34]
port 139 nsew signal output
rlabel metal2 s 51072 49600 51128 50000 6 io_out[35]
port 140 nsew signal output
rlabel metal2 s 51744 49600 51800 50000 6 io_out[36]
port 141 nsew signal output
rlabel metal2 s 52416 49600 52472 50000 6 io_out[37]
port 142 nsew signal output
rlabel metal2 s 29568 49600 29624 50000 6 io_out[3]
port 143 nsew signal output
rlabel metal2 s 30240 49600 30296 50000 6 io_out[4]
port 144 nsew signal output
rlabel metal2 s 30912 49600 30968 50000 6 io_out[5]
port 145 nsew signal output
rlabel metal2 s 31584 49600 31640 50000 6 io_out[6]
port 146 nsew signal output
rlabel metal2 s 32256 49600 32312 50000 6 io_out[7]
port 147 nsew signal output
rlabel metal2 s 32928 49600 32984 50000 6 io_out[8]
port 148 nsew signal output
rlabel metal2 s 33600 49600 33656 50000 6 io_out[9]
port 149 nsew signal output
rlabel metal2 s 53088 49600 53144 50000 6 irq[0]
port 150 nsew signal output
rlabel metal2 s 53760 49600 53816 50000 6 irq[1]
port 151 nsew signal output
rlabel metal2 s 54432 49600 54488 50000 6 irq[2]
port 152 nsew signal output
rlabel metal2 s 42224 0 42280 400 6 qcpu_do[0]
port 153 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 qcpu_do[10]
port 154 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 qcpu_do[11]
port 155 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 qcpu_do[12]
port 156 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 qcpu_do[13]
port 157 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 qcpu_do[14]
port 158 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 qcpu_do[15]
port 159 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 qcpu_do[16]
port 160 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 qcpu_do[17]
port 161 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 qcpu_do[18]
port 162 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 qcpu_do[19]
port 163 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 qcpu_do[1]
port 164 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 qcpu_do[20]
port 165 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 qcpu_do[21]
port 166 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 qcpu_do[22]
port 167 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 qcpu_do[23]
port 168 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 qcpu_do[24]
port 169 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 qcpu_do[25]
port 170 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 qcpu_do[26]
port 171 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 qcpu_do[27]
port 172 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 qcpu_do[28]
port 173 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 qcpu_do[29]
port 174 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 qcpu_do[2]
port 175 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 qcpu_do[30]
port 176 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 qcpu_do[31]
port 177 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 qcpu_do[32]
port 178 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 qcpu_do[3]
port 179 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 qcpu_do[4]
port 180 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 qcpu_do[5]
port 181 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 qcpu_do[6]
port 182 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 qcpu_do[7]
port 183 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 qcpu_do[8]
port 184 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 qcpu_do[9]
port 185 nsew signal input
rlabel metal3 s 59600 28336 60000 28392 6 qcpu_oeb[0]
port 186 nsew signal input
rlabel metal3 s 59600 31696 60000 31752 6 qcpu_oeb[10]
port 187 nsew signal input
rlabel metal3 s 59600 32032 60000 32088 6 qcpu_oeb[11]
port 188 nsew signal input
rlabel metal3 s 59600 32368 60000 32424 6 qcpu_oeb[12]
port 189 nsew signal input
rlabel metal3 s 59600 32704 60000 32760 6 qcpu_oeb[13]
port 190 nsew signal input
rlabel metal3 s 59600 33040 60000 33096 6 qcpu_oeb[14]
port 191 nsew signal input
rlabel metal3 s 59600 33376 60000 33432 6 qcpu_oeb[15]
port 192 nsew signal input
rlabel metal3 s 59600 33712 60000 33768 6 qcpu_oeb[16]
port 193 nsew signal input
rlabel metal3 s 59600 34048 60000 34104 6 qcpu_oeb[17]
port 194 nsew signal input
rlabel metal3 s 59600 34384 60000 34440 6 qcpu_oeb[18]
port 195 nsew signal input
rlabel metal3 s 59600 34720 60000 34776 6 qcpu_oeb[19]
port 196 nsew signal input
rlabel metal3 s 59600 28672 60000 28728 6 qcpu_oeb[1]
port 197 nsew signal input
rlabel metal3 s 59600 35056 60000 35112 6 qcpu_oeb[20]
port 198 nsew signal input
rlabel metal3 s 59600 35392 60000 35448 6 qcpu_oeb[21]
port 199 nsew signal input
rlabel metal3 s 59600 35728 60000 35784 6 qcpu_oeb[22]
port 200 nsew signal input
rlabel metal3 s 59600 36064 60000 36120 6 qcpu_oeb[23]
port 201 nsew signal input
rlabel metal3 s 59600 36400 60000 36456 6 qcpu_oeb[24]
port 202 nsew signal input
rlabel metal3 s 59600 36736 60000 36792 6 qcpu_oeb[25]
port 203 nsew signal input
rlabel metal3 s 59600 37072 60000 37128 6 qcpu_oeb[26]
port 204 nsew signal input
rlabel metal3 s 59600 37408 60000 37464 6 qcpu_oeb[27]
port 205 nsew signal input
rlabel metal3 s 59600 37744 60000 37800 6 qcpu_oeb[28]
port 206 nsew signal input
rlabel metal3 s 59600 38080 60000 38136 6 qcpu_oeb[29]
port 207 nsew signal input
rlabel metal3 s 59600 29008 60000 29064 6 qcpu_oeb[2]
port 208 nsew signal input
rlabel metal3 s 59600 38416 60000 38472 6 qcpu_oeb[30]
port 209 nsew signal input
rlabel metal3 s 59600 38752 60000 38808 6 qcpu_oeb[31]
port 210 nsew signal input
rlabel metal3 s 59600 39088 60000 39144 6 qcpu_oeb[32]
port 211 nsew signal input
rlabel metal3 s 59600 29344 60000 29400 6 qcpu_oeb[3]
port 212 nsew signal input
rlabel metal3 s 59600 29680 60000 29736 6 qcpu_oeb[4]
port 213 nsew signal input
rlabel metal3 s 59600 30016 60000 30072 6 qcpu_oeb[5]
port 214 nsew signal input
rlabel metal3 s 59600 30352 60000 30408 6 qcpu_oeb[6]
port 215 nsew signal input
rlabel metal3 s 59600 30688 60000 30744 6 qcpu_oeb[7]
port 216 nsew signal input
rlabel metal3 s 59600 31024 60000 31080 6 qcpu_oeb[8]
port 217 nsew signal input
rlabel metal3 s 59600 31360 60000 31416 6 qcpu_oeb[9]
port 218 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 qcpu_sram_addr[0]
port 219 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 qcpu_sram_addr[1]
port 220 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 qcpu_sram_addr[2]
port 221 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 qcpu_sram_addr[3]
port 222 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 qcpu_sram_addr[4]
port 223 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 qcpu_sram_addr[5]
port 224 nsew signal input
rlabel metal2 s 59696 0 59752 400 6 qcpu_sram_gwe
port 225 nsew signal input
rlabel metal3 s 59600 39424 60000 39480 6 qcpu_sram_in[0]
port 226 nsew signal input
rlabel metal3 s 59600 39760 60000 39816 6 qcpu_sram_in[1]
port 227 nsew signal input
rlabel metal3 s 59600 40096 60000 40152 6 qcpu_sram_in[2]
port 228 nsew signal input
rlabel metal3 s 59600 40432 60000 40488 6 qcpu_sram_in[3]
port 229 nsew signal input
rlabel metal3 s 59600 40768 60000 40824 6 qcpu_sram_in[4]
port 230 nsew signal input
rlabel metal3 s 59600 41104 60000 41160 6 qcpu_sram_in[5]
port 231 nsew signal input
rlabel metal3 s 59600 41440 60000 41496 6 qcpu_sram_in[6]
port 232 nsew signal input
rlabel metal3 s 59600 41776 60000 41832 6 qcpu_sram_in[7]
port 233 nsew signal input
rlabel metal3 s 59600 42112 60000 42168 6 qcpu_sram_out[0]
port 234 nsew signal output
rlabel metal3 s 59600 42448 60000 42504 6 qcpu_sram_out[1]
port 235 nsew signal output
rlabel metal3 s 59600 42784 60000 42840 6 qcpu_sram_out[2]
port 236 nsew signal output
rlabel metal3 s 59600 43120 60000 43176 6 qcpu_sram_out[3]
port 237 nsew signal output
rlabel metal3 s 59600 43456 60000 43512 6 qcpu_sram_out[4]
port 238 nsew signal output
rlabel metal3 s 59600 43792 60000 43848 6 qcpu_sram_out[5]
port 239 nsew signal output
rlabel metal3 s 59600 44128 60000 44184 6 qcpu_sram_out[6]
port 240 nsew signal output
rlabel metal3 s 59600 44464 60000 44520 6 qcpu_sram_out[7]
port 241 nsew signal output
rlabel metal2 s 55104 49600 55160 50000 6 rst_blinker
port 242 nsew signal output
rlabel metal3 s 0 48832 400 48888 6 rst_qcpu
port 243 nsew signal output
rlabel metal3 s 0 30800 400 30856 6 rst_sid
port 244 nsew signal output
rlabel metal2 s 57792 49600 57848 50000 6 rst_sn76489
port 245 nsew signal output
rlabel metal3 s 0 31584 400 31640 6 sid_do[0]
port 246 nsew signal input
rlabel metal3 s 0 39424 400 39480 6 sid_do[10]
port 247 nsew signal input
rlabel metal3 s 0 40208 400 40264 6 sid_do[11]
port 248 nsew signal input
rlabel metal3 s 0 40992 400 41048 6 sid_do[12]
port 249 nsew signal input
rlabel metal3 s 0 41776 400 41832 6 sid_do[13]
port 250 nsew signal input
rlabel metal3 s 0 42560 400 42616 6 sid_do[14]
port 251 nsew signal input
rlabel metal3 s 0 43344 400 43400 6 sid_do[15]
port 252 nsew signal input
rlabel metal3 s 0 44128 400 44184 6 sid_do[16]
port 253 nsew signal input
rlabel metal3 s 0 44912 400 44968 6 sid_do[17]
port 254 nsew signal input
rlabel metal3 s 0 45696 400 45752 6 sid_do[18]
port 255 nsew signal input
rlabel metal3 s 0 46480 400 46536 6 sid_do[19]
port 256 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 sid_do[1]
port 257 nsew signal input
rlabel metal3 s 0 47264 400 47320 6 sid_do[20]
port 258 nsew signal input
rlabel metal3 s 0 33152 400 33208 6 sid_do[2]
port 259 nsew signal input
rlabel metal3 s 0 33936 400 33992 6 sid_do[3]
port 260 nsew signal input
rlabel metal3 s 0 34720 400 34776 6 sid_do[4]
port 261 nsew signal input
rlabel metal3 s 0 35504 400 35560 6 sid_do[5]
port 262 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 sid_do[6]
port 263 nsew signal input
rlabel metal3 s 0 37072 400 37128 6 sid_do[7]
port 264 nsew signal input
rlabel metal3 s 0 37856 400 37912 6 sid_do[8]
port 265 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 sid_do[9]
port 266 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 sid_oeb
port 267 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 sn76489_do[0]
port 268 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 sn76489_do[10]
port 269 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 sn76489_do[11]
port 270 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 sn76489_do[12]
port 271 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 sn76489_do[13]
port 272 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 sn76489_do[14]
port 273 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 sn76489_do[15]
port 274 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 sn76489_do[16]
port 275 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 sn76489_do[17]
port 276 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 sn76489_do[18]
port 277 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 sn76489_do[19]
port 278 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 sn76489_do[1]
port 279 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 sn76489_do[20]
port 280 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 sn76489_do[21]
port 281 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 sn76489_do[22]
port 282 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 sn76489_do[23]
port 283 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 sn76489_do[24]
port 284 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 sn76489_do[25]
port 285 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 sn76489_do[26]
port 286 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 sn76489_do[27]
port 287 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 sn76489_do[2]
port 288 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 sn76489_do[3]
port 289 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 sn76489_do[4]
port 290 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 sn76489_do[5]
port 291 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 sn76489_do[6]
port 292 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 sn76489_do[7]
port 293 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 sn76489_do[8]
port 294 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 sn76489_do[9]
port 295 nsew signal input
rlabel metal4 s 2224 1538 2384 48246 6 vdd
port 296 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 48246 6 vdd
port 296 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 48246 6 vdd
port 296 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 48246 6 vdd
port 296 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 48246 6 vss
port 297 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 48246 6 vss
port 297 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 48246 6 vss
port 297 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 48246 6 vss
port 297 nsew ground bidirectional
rlabel metal2 s 112 0 168 400 6 wb_clk_i
port 298 nsew signal input
rlabel metal2 s 560 0 616 400 6 wb_rst_i
port 299 nsew signal input
rlabel metal3 s 59600 17248 60000 17304 6 wbs_ack_o
port 300 nsew signal output
rlabel metal2 s 1008 0 1064 400 6 wbs_adr_i[0]
port 301 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 wbs_adr_i[10]
port 302 nsew signal input
rlabel metal2 s 5936 0 5992 400 6 wbs_adr_i[11]
port 303 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wbs_adr_i[12]
port 304 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_adr_i[13]
port 305 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 wbs_adr_i[14]
port 306 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_adr_i[15]
port 307 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_adr_i[16]
port 308 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_adr_i[17]
port 309 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_adr_i[18]
port 310 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_adr_i[19]
port 311 nsew signal input
rlabel metal2 s 1456 0 1512 400 6 wbs_adr_i[1]
port 312 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[20]
port 313 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 wbs_adr_i[21]
port 314 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[22]
port 315 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_adr_i[23]
port 316 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_adr_i[24]
port 317 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[25]
port 318 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_adr_i[26]
port 319 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 wbs_adr_i[27]
port 320 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 wbs_adr_i[28]
port 321 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[29]
port 322 nsew signal input
rlabel metal2 s 1904 0 1960 400 6 wbs_adr_i[2]
port 323 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[30]
port 324 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_adr_i[31]
port 325 nsew signal input
rlabel metal2 s 2352 0 2408 400 6 wbs_adr_i[3]
port 326 nsew signal input
rlabel metal2 s 2800 0 2856 400 6 wbs_adr_i[4]
port 327 nsew signal input
rlabel metal2 s 3248 0 3304 400 6 wbs_adr_i[5]
port 328 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 wbs_adr_i[6]
port 329 nsew signal input
rlabel metal2 s 4144 0 4200 400 6 wbs_adr_i[7]
port 330 nsew signal input
rlabel metal2 s 4592 0 4648 400 6 wbs_adr_i[8]
port 331 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_adr_i[9]
port 332 nsew signal input
rlabel metal3 s 59600 16576 60000 16632 6 wbs_cyc_i
port 333 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_dat_i[0]
port 334 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_i[10]
port 335 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_dat_i[11]
port 336 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[12]
port 337 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_i[13]
port 338 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_dat_i[14]
port 339 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[15]
port 340 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_i[16]
port 341 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 wbs_dat_i[17]
port 342 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_i[18]
port 343 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_i[19]
port 344 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_dat_i[1]
port 345 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_dat_i[20]
port 346 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_i[21]
port 347 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 wbs_dat_i[22]
port 348 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_i[23]
port 349 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[24]
port 350 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_i[25]
port 351 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_i[26]
port 352 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_dat_i[27]
port 353 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_i[28]
port 354 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_dat_i[29]
port 355 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_i[2]
port 356 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[30]
port 357 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_i[31]
port 358 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_i[3]
port 359 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_dat_i[4]
port 360 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_i[5]
port 361 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_i[6]
port 362 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_i[7]
port 363 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_i[8]
port 364 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_i[9]
port 365 nsew signal input
rlabel metal3 s 59600 5488 60000 5544 6 wbs_dat_o[0]
port 366 nsew signal output
rlabel metal3 s 59600 8848 60000 8904 6 wbs_dat_o[10]
port 367 nsew signal output
rlabel metal3 s 59600 9184 60000 9240 6 wbs_dat_o[11]
port 368 nsew signal output
rlabel metal3 s 59600 9520 60000 9576 6 wbs_dat_o[12]
port 369 nsew signal output
rlabel metal3 s 59600 9856 60000 9912 6 wbs_dat_o[13]
port 370 nsew signal output
rlabel metal3 s 59600 10192 60000 10248 6 wbs_dat_o[14]
port 371 nsew signal output
rlabel metal3 s 59600 10528 60000 10584 6 wbs_dat_o[15]
port 372 nsew signal output
rlabel metal3 s 59600 10864 60000 10920 6 wbs_dat_o[16]
port 373 nsew signal output
rlabel metal3 s 59600 11200 60000 11256 6 wbs_dat_o[17]
port 374 nsew signal output
rlabel metal3 s 59600 11536 60000 11592 6 wbs_dat_o[18]
port 375 nsew signal output
rlabel metal3 s 59600 11872 60000 11928 6 wbs_dat_o[19]
port 376 nsew signal output
rlabel metal3 s 59600 5824 60000 5880 6 wbs_dat_o[1]
port 377 nsew signal output
rlabel metal3 s 59600 12208 60000 12264 6 wbs_dat_o[20]
port 378 nsew signal output
rlabel metal3 s 59600 12544 60000 12600 6 wbs_dat_o[21]
port 379 nsew signal output
rlabel metal3 s 59600 12880 60000 12936 6 wbs_dat_o[22]
port 380 nsew signal output
rlabel metal3 s 59600 13216 60000 13272 6 wbs_dat_o[23]
port 381 nsew signal output
rlabel metal3 s 59600 13552 60000 13608 6 wbs_dat_o[24]
port 382 nsew signal output
rlabel metal3 s 59600 13888 60000 13944 6 wbs_dat_o[25]
port 383 nsew signal output
rlabel metal3 s 59600 14224 60000 14280 6 wbs_dat_o[26]
port 384 nsew signal output
rlabel metal3 s 59600 14560 60000 14616 6 wbs_dat_o[27]
port 385 nsew signal output
rlabel metal3 s 59600 14896 60000 14952 6 wbs_dat_o[28]
port 386 nsew signal output
rlabel metal3 s 59600 15232 60000 15288 6 wbs_dat_o[29]
port 387 nsew signal output
rlabel metal3 s 59600 6160 60000 6216 6 wbs_dat_o[2]
port 388 nsew signal output
rlabel metal3 s 59600 15568 60000 15624 6 wbs_dat_o[30]
port 389 nsew signal output
rlabel metal3 s 59600 15904 60000 15960 6 wbs_dat_o[31]
port 390 nsew signal output
rlabel metal3 s 59600 6496 60000 6552 6 wbs_dat_o[3]
port 391 nsew signal output
rlabel metal3 s 59600 6832 60000 6888 6 wbs_dat_o[4]
port 392 nsew signal output
rlabel metal3 s 59600 7168 60000 7224 6 wbs_dat_o[5]
port 393 nsew signal output
rlabel metal3 s 59600 7504 60000 7560 6 wbs_dat_o[6]
port 394 nsew signal output
rlabel metal3 s 59600 7840 60000 7896 6 wbs_dat_o[7]
port 395 nsew signal output
rlabel metal3 s 59600 8176 60000 8232 6 wbs_dat_o[8]
port 396 nsew signal output
rlabel metal3 s 59600 8512 60000 8568 6 wbs_dat_o[9]
port 397 nsew signal output
rlabel metal3 s 59600 16912 60000 16968 6 wbs_stb_i
port 398 nsew signal input
rlabel metal3 s 59600 16240 60000 16296 6 wbs_we_i
port 399 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7898606
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1_group/openlane/Multiplexer/runs/23_11_02_21_18/results/signoff/multiplexer.magic.gds
string GDS_START 359086
<< end >>

