VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_mc14500
  CLASS BLOCK ;
  FOREIGN wrapped_mc14500 ;
  ORIGIN 0.000 0.000 ;
  SIZE 185.000 BY 185.000 ;
  PIN SDI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 145.600 185.000 146.160 ;
    END
  END SDI
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 11.200 185.000 11.760 ;
    END
  END clk_i
  PIN custom_setting
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 172.480 185.000 173.040 ;
    END
  END custom_setting
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 38.080 185.000 38.640 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 51.520 185.000 52.080 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 64.960 185.000 65.520 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 78.400 185.000 78.960 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 91.840 185.000 92.400 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 105.280 185.000 105.840 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 118.720 185.000 119.280 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 132.160 185.000 132.720 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 181.000 8.400 185.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 181.000 64.400 185.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 181.000 70.000 185.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 181.000 75.600 185.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 181.000 81.200 185.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 181.000 86.800 185.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 181.000 92.400 185.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 181.000 98.000 185.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 181.000 103.600 185.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 181.000 109.200 185.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 181.000 114.800 185.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 181.000 14.000 185.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 181.000 120.400 185.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 181.000 126.000 185.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 181.000 131.600 185.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 181.000 137.200 185.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 181.000 142.800 185.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 181.000 148.400 185.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 181.000 154.000 185.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 181.000 159.600 185.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 181.000 165.200 185.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 181.000 170.800 185.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 181.000 19.600 185.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 181.000 176.400 185.000 ;
    END
  END io_out[30]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 181.000 25.200 185.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 181.000 30.800 185.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 181.000 36.400 185.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 181.000 42.000 185.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 181.000 47.600 185.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 181.000 53.200 185.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 181.000 58.800 185.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 24.640 185.000 25.200 ;
    END
  END rst_n
  PIN sram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 8.960 0.000 9.520 4.000 ;
    END
  END sram_addr[0]
  PIN sram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END sram_addr[1]
  PIN sram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 24.640 0.000 25.200 4.000 ;
    END
  END sram_addr[2]
  PIN sram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END sram_addr[3]
  PIN sram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END sram_addr[4]
  PIN sram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 0.000 48.720 4.000 ;
    END
  END sram_addr[5]
  PIN sram_gwe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 181.000 159.040 185.000 159.600 ;
    END
  END sram_gwe
  PIN sram_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END sram_in[0]
  PIN sram_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END sram_in[1]
  PIN sram_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END sram_in[2]
  PIN sram_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END sram_in[3]
  PIN sram_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END sram_in[4]
  PIN sram_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END sram_in[5]
  PIN sram_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 4.000 ;
    END
  END sram_in[6]
  PIN sram_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END sram_in[7]
  PIN sram_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END sram_out[0]
  PIN sram_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END sram_out[1]
  PIN sram_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END sram_out[2]
  PIN sram_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 0.000 142.800 4.000 ;
    END
  END sram_out[3]
  PIN sram_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END sram_out[4]
  PIN sram_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END sram_out[5]
  PIN sram_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 0.000 166.320 4.000 ;
    END
  END sram_out[6]
  PIN sram_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END sram_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 27.340 15.380 28.940 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.180 15.380 71.780 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 113.020 15.380 114.620 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 155.860 15.380 157.460 168.860 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 48.760 15.380 50.360 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 91.600 15.380 93.200 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134.440 15.380 136.040 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.280 15.380 178.880 168.860 ;
    END
  END vss
  OBS
      LAYER Nwell ;
        RECT 6.290 166.525 178.510 168.990 ;
        RECT 6.290 166.400 69.825 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 178.510 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 34.545 162.880 ;
        RECT 6.290 158.685 178.510 162.755 ;
        RECT 6.290 158.560 46.865 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 178.510 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 26.145 155.040 ;
        RECT 6.290 150.845 178.510 154.915 ;
        RECT 6.290 150.720 124.705 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 178.510 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 23.345 147.200 ;
        RECT 6.290 142.880 178.510 147.075 ;
      LAYER Pwell ;
        RECT 6.290 139.360 178.510 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 21.665 139.360 ;
        RECT 6.290 135.165 178.510 139.235 ;
        RECT 6.290 135.040 46.910 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 178.510 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 22.225 131.520 ;
        RECT 6.290 127.325 178.510 131.395 ;
        RECT 6.290 127.200 121.345 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 178.510 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 130.305 123.680 ;
        RECT 6.290 119.485 178.510 123.555 ;
        RECT 6.290 119.360 165.585 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 178.510 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 23.905 115.840 ;
        RECT 6.290 111.645 178.510 115.715 ;
        RECT 6.290 111.520 41.265 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 178.510 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 22.225 108.000 ;
        RECT 6.290 103.805 178.510 107.875 ;
        RECT 6.290 103.680 53.585 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 178.510 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 28.945 100.160 ;
        RECT 6.290 95.965 178.510 100.035 ;
        RECT 6.290 95.840 32.305 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 178.510 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 73.745 92.320 ;
        RECT 6.290 88.125 178.510 92.195 ;
        RECT 6.290 88.000 40.705 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 178.510 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 63.665 84.480 ;
        RECT 6.290 80.285 178.510 84.355 ;
        RECT 6.290 80.160 54.145 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 178.510 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 93.505 76.640 ;
        RECT 6.290 72.445 178.510 76.515 ;
        RECT 6.290 72.320 72.625 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 178.510 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 51.905 68.800 ;
        RECT 6.290 64.605 178.510 68.675 ;
        RECT 6.290 64.480 132.760 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 178.510 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 33.640 60.960 ;
        RECT 6.290 56.765 178.510 60.835 ;
        RECT 6.290 56.640 37.560 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 178.510 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 65.905 53.120 ;
        RECT 6.290 48.925 178.510 52.995 ;
        RECT 6.290 48.800 39.025 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 178.510 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 30.280 45.280 ;
        RECT 6.290 41.085 178.510 45.155 ;
        RECT 6.290 40.960 58.280 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 178.510 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 64.785 37.440 ;
        RECT 6.290 33.245 178.510 37.315 ;
        RECT 6.290 33.120 84.600 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 178.510 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 62.545 29.600 ;
        RECT 6.290 25.405 178.510 29.475 ;
        RECT 6.290 25.280 34.545 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 178.510 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 33.425 21.760 ;
        RECT 6.290 17.440 178.510 21.635 ;
      LAYER Pwell ;
        RECT 6.290 15.250 178.510 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 178.880 168.860 ;
      LAYER Metal2 ;
        RECT 8.700 180.700 13.140 181.300 ;
        RECT 14.300 180.700 18.740 181.300 ;
        RECT 19.900 180.700 24.340 181.300 ;
        RECT 25.500 180.700 29.940 181.300 ;
        RECT 31.100 180.700 35.540 181.300 ;
        RECT 36.700 180.700 41.140 181.300 ;
        RECT 42.300 180.700 46.740 181.300 ;
        RECT 47.900 180.700 52.340 181.300 ;
        RECT 53.500 180.700 57.940 181.300 ;
        RECT 59.100 180.700 63.540 181.300 ;
        RECT 64.700 180.700 69.140 181.300 ;
        RECT 70.300 180.700 74.740 181.300 ;
        RECT 75.900 180.700 80.340 181.300 ;
        RECT 81.500 180.700 85.940 181.300 ;
        RECT 87.100 180.700 91.540 181.300 ;
        RECT 92.700 180.700 97.140 181.300 ;
        RECT 98.300 180.700 102.740 181.300 ;
        RECT 103.900 180.700 108.340 181.300 ;
        RECT 109.500 180.700 113.940 181.300 ;
        RECT 115.100 180.700 119.540 181.300 ;
        RECT 120.700 180.700 125.140 181.300 ;
        RECT 126.300 180.700 130.740 181.300 ;
        RECT 131.900 180.700 136.340 181.300 ;
        RECT 137.500 180.700 141.940 181.300 ;
        RECT 143.100 180.700 147.540 181.300 ;
        RECT 148.700 180.700 153.140 181.300 ;
        RECT 154.300 180.700 158.740 181.300 ;
        RECT 159.900 180.700 164.340 181.300 ;
        RECT 165.500 180.700 169.940 181.300 ;
        RECT 171.100 180.700 175.540 181.300 ;
        RECT 176.700 180.700 181.300 181.300 ;
        RECT 7.980 4.300 181.300 180.700 ;
        RECT 7.980 4.000 8.660 4.300 ;
        RECT 9.820 4.000 16.500 4.300 ;
        RECT 17.660 4.000 24.340 4.300 ;
        RECT 25.500 4.000 32.180 4.300 ;
        RECT 33.340 4.000 40.020 4.300 ;
        RECT 41.180 4.000 47.860 4.300 ;
        RECT 49.020 4.000 55.700 4.300 ;
        RECT 56.860 4.000 63.540 4.300 ;
        RECT 64.700 4.000 71.380 4.300 ;
        RECT 72.540 4.000 79.220 4.300 ;
        RECT 80.380 4.000 87.060 4.300 ;
        RECT 88.220 4.000 94.900 4.300 ;
        RECT 96.060 4.000 102.740 4.300 ;
        RECT 103.900 4.000 110.580 4.300 ;
        RECT 111.740 4.000 118.420 4.300 ;
        RECT 119.580 4.000 126.260 4.300 ;
        RECT 127.420 4.000 134.100 4.300 ;
        RECT 135.260 4.000 141.940 4.300 ;
        RECT 143.100 4.000 149.780 4.300 ;
        RECT 150.940 4.000 157.620 4.300 ;
        RECT 158.780 4.000 165.460 4.300 ;
        RECT 166.620 4.000 173.300 4.300 ;
        RECT 174.460 4.000 181.300 4.300 ;
      LAYER Metal3 ;
        RECT 18.010 172.180 180.700 172.900 ;
        RECT 18.010 159.900 181.350 172.180 ;
        RECT 18.010 158.740 180.700 159.900 ;
        RECT 18.010 146.460 181.350 158.740 ;
        RECT 18.010 145.300 180.700 146.460 ;
        RECT 18.010 133.020 181.350 145.300 ;
        RECT 18.010 131.860 180.700 133.020 ;
        RECT 18.010 119.580 181.350 131.860 ;
        RECT 18.010 118.420 180.700 119.580 ;
        RECT 18.010 106.140 181.350 118.420 ;
        RECT 18.010 104.980 180.700 106.140 ;
        RECT 18.010 92.700 181.350 104.980 ;
        RECT 18.010 91.540 180.700 92.700 ;
        RECT 18.010 79.260 181.350 91.540 ;
        RECT 18.010 78.100 180.700 79.260 ;
        RECT 18.010 65.820 181.350 78.100 ;
        RECT 18.010 64.660 180.700 65.820 ;
        RECT 18.010 52.380 181.350 64.660 ;
        RECT 18.010 51.220 180.700 52.380 ;
        RECT 18.010 38.940 181.350 51.220 ;
        RECT 18.010 37.780 180.700 38.940 ;
        RECT 18.010 25.500 181.350 37.780 ;
        RECT 18.010 24.340 180.700 25.500 ;
        RECT 18.010 12.060 181.350 24.340 ;
        RECT 18.010 11.340 180.700 12.060 ;
      LAYER Metal4 ;
        RECT 38.220 26.410 48.460 155.590 ;
        RECT 50.660 26.410 69.880 155.590 ;
        RECT 72.080 26.410 91.300 155.590 ;
        RECT 93.500 26.410 112.720 155.590 ;
        RECT 114.920 26.410 134.140 155.590 ;
        RECT 136.340 26.410 155.560 155.590 ;
        RECT 157.760 26.410 175.700 155.590 ;
  END
END wrapped_mc14500
END LIBRARY

