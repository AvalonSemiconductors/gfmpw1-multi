magic
tech gf180mcuD
magscale 1 10
timestamp 1753964058
<< metal1 >>
rect 6906 22878 6918 22930
rect 6970 22927 6982 22930
rect 7746 22927 7758 22930
rect 6970 22881 7758 22927
rect 6970 22878 6982 22881
rect 7746 22878 7758 22881
rect 7810 22878 7822 22930
rect 1344 22762 24640 22796
rect 1344 22710 4126 22762
rect 4178 22710 4230 22762
rect 4282 22710 4334 22762
rect 4386 22710 9950 22762
rect 10002 22710 10054 22762
rect 10106 22710 10158 22762
rect 10210 22710 15774 22762
rect 15826 22710 15878 22762
rect 15930 22710 15982 22762
rect 16034 22710 21598 22762
rect 21650 22710 21702 22762
rect 21754 22710 21806 22762
rect 21858 22710 24640 22762
rect 1344 22676 24640 22710
rect 22542 22594 22594 22606
rect 6906 22542 6918 22594
rect 6970 22542 6982 22594
rect 7858 22486 7870 22538
rect 7922 22486 7934 22538
rect 22542 22530 22594 22542
rect 12126 22482 12178 22494
rect 21186 22430 21198 22482
rect 21250 22430 21262 22482
rect 12126 22418 12178 22430
rect 7198 22370 7250 22382
rect 7198 22306 7250 22318
rect 7422 22370 7474 22382
rect 11454 22370 11506 22382
rect 11732 22370 11784 22382
rect 7746 22318 7758 22370
rect 7810 22318 7822 22370
rect 8082 22318 8094 22370
rect 8146 22318 8158 22370
rect 11554 22318 11566 22370
rect 11618 22318 11630 22370
rect 7422 22306 7474 22318
rect 11454 22306 11506 22318
rect 11732 22306 11784 22318
rect 13582 22370 13634 22382
rect 13582 22306 13634 22318
rect 13974 22370 14026 22382
rect 13974 22306 14026 22318
rect 19742 22370 19794 22382
rect 20738 22318 20750 22370
rect 20802 22318 20814 22370
rect 19742 22306 19794 22318
rect 21074 22274 21086 22326
rect 21138 22274 21150 22326
rect 21522 22290 21534 22342
rect 21586 22290 21598 22342
rect 19574 22258 19626 22270
rect 19574 22194 19626 22206
rect 8598 22146 8650 22158
rect 8598 22082 8650 22094
rect 13246 22146 13298 22158
rect 13246 22082 13298 22094
rect 20078 22146 20130 22158
rect 20078 22082 20130 22094
rect 1344 21978 24800 22012
rect 1344 21926 7038 21978
rect 7090 21926 7142 21978
rect 7194 21926 7246 21978
rect 7298 21926 12862 21978
rect 12914 21926 12966 21978
rect 13018 21926 13070 21978
rect 13122 21926 18686 21978
rect 18738 21926 18790 21978
rect 18842 21926 18894 21978
rect 18946 21926 24510 21978
rect 24562 21926 24614 21978
rect 24666 21926 24718 21978
rect 24770 21926 24800 21978
rect 1344 21892 24800 21926
rect 7422 21698 7474 21710
rect 7422 21634 7474 21646
rect 7814 21642 7866 21654
rect 4734 21586 4786 21598
rect 8418 21590 8430 21642
rect 8482 21590 8494 21642
rect 7814 21578 7866 21590
rect 10782 21586 10834 21598
rect 8194 21534 8206 21586
rect 8258 21534 8270 21586
rect 9893 21534 9905 21586
rect 9957 21534 9969 21586
rect 4734 21522 4786 21534
rect 10782 21522 10834 21534
rect 11678 21586 11730 21598
rect 11678 21522 11730 21534
rect 14702 21586 14754 21598
rect 15598 21586 15650 21598
rect 14914 21534 14926 21586
rect 14978 21534 14990 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 14702 21522 14754 21534
rect 15598 21522 15650 21534
rect 17278 21586 17330 21598
rect 17278 21522 17330 21534
rect 20862 21586 20914 21598
rect 20862 21522 20914 21534
rect 7982 21474 8034 21486
rect 5506 21422 5518 21474
rect 5570 21422 5582 21474
rect 7982 21410 8034 21422
rect 11342 21474 11394 21486
rect 24278 21474 24330 21486
rect 12002 21422 12014 21474
rect 12066 21422 12078 21474
rect 13906 21422 13918 21474
rect 13970 21422 13982 21474
rect 18050 21422 18062 21474
rect 18114 21422 18126 21474
rect 19954 21422 19966 21474
rect 20018 21422 20030 21474
rect 21634 21422 21646 21474
rect 21698 21422 21710 21474
rect 23538 21422 23550 21474
rect 23602 21422 23614 21474
rect 11342 21410 11394 21422
rect 9662 21362 9714 21374
rect 15250 21366 15262 21418
rect 15314 21366 15326 21418
rect 24278 21410 24330 21422
rect 9662 21298 9714 21310
rect 15934 21362 15986 21374
rect 15934 21298 15986 21310
rect 1344 21194 24640 21228
rect 1344 21142 4126 21194
rect 4178 21142 4230 21194
rect 4282 21142 4334 21194
rect 4386 21142 9950 21194
rect 10002 21142 10054 21194
rect 10106 21142 10158 21194
rect 10210 21142 15774 21194
rect 15826 21142 15878 21194
rect 15930 21142 15982 21194
rect 16034 21142 21598 21194
rect 21650 21142 21702 21194
rect 21754 21142 21806 21194
rect 21858 21142 24640 21194
rect 1344 21108 24640 21142
rect 10446 20970 10498 20982
rect 12126 20970 12178 20982
rect 8822 20914 8874 20926
rect 8822 20850 8874 20862
rect 9550 20914 9602 20926
rect 11442 20918 11454 20970
rect 11506 20918 11518 20970
rect 10446 20906 10498 20918
rect 12126 20906 12178 20918
rect 14926 20970 14978 20982
rect 21354 20974 21366 21026
rect 21418 20974 21430 21026
rect 14926 20906 14978 20918
rect 15922 20862 15934 20914
rect 15986 20862 15998 20914
rect 17826 20862 17838 20914
rect 17890 20862 17902 20914
rect 19282 20862 19294 20914
rect 19346 20862 19358 20914
rect 9550 20850 9602 20862
rect 5518 20802 5570 20814
rect 9886 20802 9938 20814
rect 15150 20802 15202 20814
rect 20302 20802 20354 20814
rect 6290 20750 6302 20802
rect 6354 20750 6366 20802
rect 9202 20750 9214 20802
rect 9266 20750 9278 20802
rect 9662 20763 9714 20775
rect 5518 20738 5570 20750
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 10882 20750 10894 20802
rect 10946 20750 10958 20802
rect 11330 20750 11342 20802
rect 11394 20750 11406 20802
rect 11666 20750 11678 20802
rect 11730 20750 11742 20802
rect 12226 20750 12238 20802
rect 12290 20750 12302 20802
rect 9886 20738 9938 20750
rect 12902 20712 12914 20764
rect 12966 20712 12978 20764
rect 14126 20712 14138 20764
rect 14190 20712 14202 20764
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 18946 20750 18958 20802
rect 19010 20750 19022 20802
rect 15150 20738 15202 20750
rect 8206 20690 8258 20702
rect 9662 20699 9714 20711
rect 19170 20706 19182 20758
rect 19234 20706 19246 20758
rect 19618 20750 19630 20802
rect 19682 20750 19694 20802
rect 19898 20694 19910 20746
rect 19962 20694 19974 20746
rect 20302 20738 20354 20750
rect 21646 20802 21698 20814
rect 21646 20738 21698 20750
rect 21870 20802 21922 20814
rect 21870 20738 21922 20750
rect 22206 20802 22258 20814
rect 24334 20802 24386 20814
rect 23070 20750 23082 20802
rect 23134 20750 23146 20802
rect 22206 20738 22258 20750
rect 24334 20738 24386 20750
rect 8206 20626 8258 20638
rect 23326 20690 23378 20702
rect 19730 20582 19742 20634
rect 19794 20582 19806 20634
rect 23326 20626 23378 20638
rect 23998 20578 24050 20590
rect 23998 20514 24050 20526
rect 1344 20410 24800 20444
rect 1344 20358 7038 20410
rect 7090 20358 7142 20410
rect 7194 20358 7246 20410
rect 7298 20358 12862 20410
rect 12914 20358 12966 20410
rect 13018 20358 13070 20410
rect 13122 20358 18686 20410
rect 18738 20358 18790 20410
rect 18842 20358 18894 20410
rect 18946 20358 24510 20410
rect 24562 20358 24614 20410
rect 24666 20358 24718 20410
rect 24770 20358 24800 20410
rect 1344 20324 24800 20358
rect 4678 20242 4730 20254
rect 4678 20178 4730 20190
rect 5854 20242 5906 20254
rect 18062 20242 18114 20254
rect 12226 20190 12238 20242
rect 12290 20239 12302 20242
rect 12674 20239 12686 20242
rect 12290 20193 12686 20239
rect 12290 20190 12302 20193
rect 12674 20190 12686 20193
rect 12738 20190 12750 20242
rect 5854 20178 5906 20190
rect 8194 20134 8206 20186
rect 8258 20134 8270 20186
rect 18062 20178 18114 20190
rect 22318 20242 22370 20254
rect 20526 20130 20578 20142
rect 21522 20134 21534 20186
rect 21586 20134 21598 20186
rect 22318 20178 22370 20190
rect 8542 20057 8594 20069
rect 6190 20018 6242 20030
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 15296 20056 15348 20068
rect 8542 19993 8594 20005
rect 8766 20018 8818 20030
rect 6190 19954 6242 19966
rect 8766 19954 8818 19966
rect 9662 20018 9714 20030
rect 9662 19954 9714 19966
rect 9886 20018 9938 20030
rect 9886 19954 9938 19966
rect 10446 20018 10498 20030
rect 10446 19954 10498 19966
rect 10670 20018 10722 20030
rect 10670 19954 10722 19966
rect 11230 20018 11282 20030
rect 11230 19954 11282 19966
rect 11454 20018 11506 20030
rect 11454 19954 11506 19966
rect 15038 20018 15090 20030
rect 15138 19966 15150 20018
rect 15202 19966 15214 20018
rect 15296 19992 15348 20004
rect 18398 20018 18450 20030
rect 15038 19954 15090 19966
rect 18398 19954 18450 19966
rect 19406 20018 19458 20030
rect 19406 19954 19458 19966
rect 19742 20018 19794 20030
rect 19742 19954 19794 19966
rect 20190 20018 20242 20030
rect 20346 20022 20358 20074
rect 20410 20022 20422 20074
rect 20526 20066 20578 20078
rect 21590 20047 21642 20059
rect 20190 19954 20242 19966
rect 20638 20018 20690 20030
rect 21298 19966 21310 20018
rect 21362 19966 21374 20018
rect 21590 19983 21642 19995
rect 22878 20018 22930 20030
rect 23742 20022 23754 20074
rect 23806 20022 23818 20074
rect 20638 19954 20690 19966
rect 22654 19962 22706 19974
rect 15710 19906 15762 19918
rect 11722 19854 11734 19906
rect 11786 19854 11798 19906
rect 15710 19842 15762 19854
rect 18790 19906 18842 19918
rect 18790 19842 18842 19854
rect 19238 19906 19290 19918
rect 22878 19954 22930 19966
rect 22654 19898 22706 19910
rect 19238 19842 19290 19854
rect 5014 19794 5066 19806
rect 20918 19794 20970 19806
rect 10154 19742 10166 19794
rect 10218 19742 10230 19794
rect 10938 19742 10950 19794
rect 11002 19742 11014 19794
rect 5014 19730 5066 19742
rect 20918 19730 20970 19742
rect 23998 19794 24050 19806
rect 23998 19730 24050 19742
rect 1344 19626 24640 19660
rect 1344 19574 4126 19626
rect 4178 19574 4230 19626
rect 4282 19574 4334 19626
rect 4386 19574 9950 19626
rect 10002 19574 10054 19626
rect 10106 19574 10158 19626
rect 10210 19574 15774 19626
rect 15826 19574 15878 19626
rect 15930 19574 15982 19626
rect 16034 19574 21598 19626
rect 21650 19574 21702 19626
rect 21754 19574 21806 19626
rect 21858 19574 24640 19626
rect 1344 19540 24640 19574
rect 7982 19458 8034 19470
rect 7982 19394 8034 19406
rect 9494 19402 9546 19414
rect 20346 19406 20358 19458
rect 20410 19406 20422 19458
rect 9494 19338 9546 19350
rect 22598 19346 22650 19358
rect 9874 19294 9886 19346
rect 9938 19294 9950 19346
rect 12070 19290 12122 19302
rect 13570 19294 13582 19346
rect 13634 19294 13646 19346
rect 21298 19294 21310 19346
rect 21362 19294 21374 19346
rect 2046 19234 2098 19246
rect 8318 19234 8370 19246
rect 2818 19182 2830 19234
rect 2882 19182 2894 19234
rect 5506 19182 5518 19234
rect 5570 19182 5582 19234
rect 2046 19170 2098 19182
rect 8318 19170 8370 19182
rect 8654 19234 8706 19246
rect 10670 19234 10722 19246
rect 9650 19182 9662 19234
rect 9714 19182 9726 19234
rect 8654 19170 8706 19182
rect 9986 19138 9998 19190
rect 10050 19138 10062 19190
rect 10210 19182 10222 19234
rect 10274 19182 10286 19234
rect 10670 19170 10722 19182
rect 10838 19234 10890 19246
rect 10838 19170 10890 19182
rect 11118 19234 11170 19246
rect 11118 19170 11170 19182
rect 11398 19234 11450 19246
rect 11398 19170 11450 19182
rect 11902 19234 11954 19246
rect 22598 19282 22650 19294
rect 12070 19226 12122 19238
rect 12350 19234 12402 19246
rect 16270 19234 16322 19246
rect 11902 19170 11954 19182
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 12350 19170 12402 19182
rect 16270 19170 16322 19182
rect 16830 19234 16882 19246
rect 20638 19234 20690 19246
rect 17602 19182 17614 19234
rect 17666 19182 17678 19234
rect 16830 19170 16882 19182
rect 20638 19170 20690 19182
rect 20862 19234 20914 19246
rect 24110 19234 24162 19246
rect 20862 19170 20914 19182
rect 21410 19138 21422 19190
rect 21474 19138 21486 19190
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 23221 19182 23233 19234
rect 23285 19182 23297 19234
rect 24110 19170 24162 19182
rect 4734 19122 4786 19134
rect 4734 19058 4786 19070
rect 8990 19122 9042 19134
rect 8990 19058 9042 19070
rect 11006 19122 11058 19134
rect 11006 19058 11058 19070
rect 12238 19122 12290 19134
rect 12238 19058 12290 19070
rect 12630 19122 12682 19134
rect 12630 19058 12682 19070
rect 19518 19122 19570 19134
rect 19518 19058 19570 19070
rect 22990 19122 23042 19134
rect 22990 19058 23042 19070
rect 5686 19010 5738 19022
rect 5686 18946 5738 18958
rect 6246 19010 6298 19022
rect 6246 18946 6298 18958
rect 1344 18842 24800 18876
rect 1344 18790 7038 18842
rect 7090 18790 7142 18842
rect 7194 18790 7246 18842
rect 7298 18790 12862 18842
rect 12914 18790 12966 18842
rect 13018 18790 13070 18842
rect 13122 18790 18686 18842
rect 18738 18790 18790 18842
rect 18842 18790 18894 18842
rect 18946 18790 24510 18842
rect 24562 18790 24614 18842
rect 24666 18790 24718 18842
rect 24770 18790 24800 18842
rect 1344 18756 24800 18790
rect 17838 18674 17890 18686
rect 17838 18610 17890 18622
rect 20178 18566 20190 18618
rect 20242 18566 20254 18618
rect 1598 18450 1650 18462
rect 1598 18386 1650 18398
rect 4286 18450 4338 18462
rect 4286 18386 4338 18398
rect 5070 18450 5122 18462
rect 5070 18386 5122 18398
rect 5294 18450 5346 18462
rect 5294 18386 5346 18398
rect 5854 18450 5906 18462
rect 7870 18450 7922 18462
rect 12910 18450 12962 18462
rect 6718 18398 6730 18450
rect 6782 18398 6794 18450
rect 10994 18398 11006 18450
rect 11058 18398 11070 18450
rect 11330 18398 11342 18450
rect 11394 18398 11406 18450
rect 12002 18398 12014 18450
rect 12066 18398 12078 18450
rect 5854 18386 5906 18398
rect 7870 18386 7922 18398
rect 12910 18386 12962 18398
rect 13358 18450 13410 18462
rect 13358 18386 13410 18398
rect 13694 18450 13746 18462
rect 13694 18386 13746 18398
rect 15150 18450 15202 18462
rect 15150 18386 15202 18398
rect 18174 18450 18226 18462
rect 20402 18454 20414 18506
rect 20466 18454 20478 18506
rect 20638 18450 20690 18462
rect 19954 18398 19966 18450
rect 20018 18398 20030 18450
rect 18174 18386 18226 18398
rect 20638 18386 20690 18398
rect 22766 18450 22818 18462
rect 23426 18454 23438 18506
rect 23490 18454 23502 18506
rect 23662 18450 23714 18462
rect 22978 18398 22990 18450
rect 23042 18398 23054 18450
rect 22766 18386 22818 18398
rect 23662 18386 23714 18398
rect 23998 18450 24050 18462
rect 23998 18386 24050 18398
rect 22038 18338 22090 18350
rect 2370 18286 2382 18338
rect 2434 18286 2446 18338
rect 6974 18226 7026 18238
rect 4778 18174 4790 18226
rect 4842 18174 4854 18226
rect 6974 18162 7026 18174
rect 7534 18226 7586 18238
rect 11106 18230 11118 18282
rect 11170 18230 11182 18282
rect 22038 18274 22090 18286
rect 23326 18338 23378 18350
rect 23326 18274 23378 18286
rect 7534 18162 7586 18174
rect 11846 18226 11898 18238
rect 11846 18162 11898 18174
rect 12574 18226 12626 18238
rect 12574 18162 12626 18174
rect 15486 18226 15538 18238
rect 15486 18162 15538 18174
rect 22430 18226 22482 18238
rect 22430 18162 22482 18174
rect 1344 18058 24640 18092
rect 1344 18006 4126 18058
rect 4178 18006 4230 18058
rect 4282 18006 4334 18058
rect 4386 18006 9950 18058
rect 10002 18006 10054 18058
rect 10106 18006 10158 18058
rect 10210 18006 15774 18058
rect 15826 18006 15878 18058
rect 15930 18006 15982 18058
rect 16034 18006 21598 18058
rect 21650 18006 21702 18058
rect 21754 18006 21806 18058
rect 21858 18006 24640 18058
rect 1344 17972 24640 18006
rect 11566 17890 11618 17902
rect 4286 17834 4338 17846
rect 11566 17826 11618 17838
rect 13694 17890 13746 17902
rect 4286 17770 4338 17782
rect 5742 17778 5794 17790
rect 12226 17782 12238 17834
rect 12290 17782 12302 17834
rect 13694 17826 13746 17838
rect 14578 17726 14590 17778
rect 14642 17726 14654 17778
rect 16482 17726 16494 17778
rect 16546 17726 16558 17778
rect 5742 17714 5794 17726
rect 4958 17666 5010 17678
rect 3938 17614 3950 17666
rect 4002 17614 4014 17666
rect 4162 17614 4174 17666
rect 4226 17614 4238 17666
rect 4666 17614 4678 17666
rect 4730 17614 4742 17666
rect 4958 17602 5010 17614
rect 5182 17666 5234 17678
rect 5182 17602 5234 17614
rect 6134 17666 6186 17678
rect 6414 17666 6466 17678
rect 6290 17614 6302 17666
rect 6354 17614 6366 17666
rect 6134 17602 6186 17614
rect 6414 17602 6466 17614
rect 6750 17666 6802 17678
rect 7926 17666 7978 17678
rect 7410 17614 7422 17666
rect 7474 17614 7486 17666
rect 6750 17602 6802 17614
rect 7926 17602 7978 17614
rect 8206 17666 8258 17678
rect 8486 17666 8538 17678
rect 8306 17614 8318 17666
rect 8370 17614 8382 17666
rect 8206 17602 8258 17614
rect 8486 17602 8538 17614
rect 8654 17666 8706 17678
rect 8654 17602 8706 17614
rect 8878 17666 8930 17678
rect 8878 17602 8930 17614
rect 11118 17666 11170 17678
rect 11118 17602 11170 17614
rect 11902 17666 11954 17678
rect 13358 17666 13410 17678
rect 12226 17614 12238 17666
rect 12290 17614 12302 17666
rect 12450 17614 12462 17666
rect 12514 17614 12526 17666
rect 11902 17602 11954 17614
rect 13358 17602 13410 17614
rect 17278 17666 17330 17678
rect 17278 17602 17330 17614
rect 17390 17666 17442 17678
rect 22094 17666 22146 17678
rect 18162 17614 18174 17666
rect 18226 17614 18238 17666
rect 17390 17602 17442 17614
rect 22094 17602 22146 17614
rect 24334 17666 24386 17678
rect 20078 17554 20130 17566
rect 22958 17558 22970 17610
rect 23022 17558 23034 17610
rect 24334 17602 24386 17614
rect 7522 17446 7534 17498
rect 7586 17446 7598 17498
rect 20078 17490 20130 17502
rect 23214 17554 23266 17566
rect 23214 17490 23266 17502
rect 9214 17442 9266 17454
rect 9214 17378 9266 17390
rect 10782 17442 10834 17454
rect 10782 17378 10834 17390
rect 23998 17442 24050 17454
rect 23998 17378 24050 17390
rect 1344 17274 24800 17308
rect 1344 17222 7038 17274
rect 7090 17222 7142 17274
rect 7194 17222 7246 17274
rect 7298 17222 12862 17274
rect 12914 17222 12966 17274
rect 13018 17222 13070 17274
rect 13122 17222 18686 17274
rect 18738 17222 18790 17274
rect 18842 17222 18894 17274
rect 18946 17222 24510 17274
rect 24562 17222 24614 17274
rect 24666 17222 24718 17274
rect 24770 17222 24800 17274
rect 1344 17188 24800 17222
rect 18174 17106 18226 17118
rect 3266 16998 3278 17050
rect 3330 16998 3342 17050
rect 6190 16994 6242 17006
rect 4062 16938 4114 16950
rect 3726 16882 3778 16894
rect 3042 16830 3054 16882
rect 3106 16830 3118 16882
rect 4162 16886 4174 16938
rect 4226 16886 4238 16938
rect 4386 16886 4398 16938
rect 4450 16886 4462 16938
rect 4610 16886 4622 16938
rect 4674 16886 4686 16938
rect 4062 16874 4114 16886
rect 5854 16882 5906 16894
rect 6010 16886 6022 16938
rect 6074 16886 6086 16938
rect 6190 16930 6242 16942
rect 6582 16994 6634 17006
rect 12562 16998 12574 17050
rect 12626 16998 12638 17050
rect 18174 17042 18226 17054
rect 6582 16930 6634 16942
rect 15430 16994 15482 17006
rect 20178 16998 20190 17050
rect 20242 16998 20254 17050
rect 21522 16998 21534 17050
rect 21586 16998 21598 17050
rect 23090 16998 23102 17050
rect 23154 16998 23166 17050
rect 8504 16920 8556 16932
rect 3726 16818 3778 16830
rect 5854 16818 5906 16830
rect 6302 16882 6354 16894
rect 7926 16882 7978 16894
rect 6850 16830 6862 16882
rect 6914 16830 6926 16882
rect 6302 16818 6354 16830
rect 7926 16818 7978 16830
rect 8206 16882 8258 16894
rect 8306 16830 8318 16882
rect 8370 16830 8382 16882
rect 9874 16886 9886 16938
rect 9938 16886 9950 16938
rect 14590 16917 14642 16929
rect 10222 16882 10274 16894
rect 8504 16856 8556 16868
rect 9538 16830 9550 16882
rect 9602 16830 9614 16882
rect 8206 16818 8258 16830
rect 10222 16818 10274 16830
rect 10558 16882 10610 16894
rect 10558 16818 10610 16830
rect 11790 16882 11842 16894
rect 12910 16882 12962 16894
rect 12338 16830 12350 16882
rect 12402 16830 12414 16882
rect 11790 16818 11842 16830
rect 12910 16818 12962 16830
rect 13134 16882 13186 16894
rect 13402 16830 13414 16882
rect 13466 16830 13478 16882
rect 14590 16853 14642 16865
rect 14702 16910 14754 16922
rect 14702 16846 14754 16858
rect 14926 16910 14978 16922
rect 15138 16886 15150 16938
rect 15202 16886 15214 16938
rect 15430 16930 15482 16942
rect 14926 16846 14978 16858
rect 18510 16882 18562 16894
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 19618 16845 19630 16897
rect 19682 16845 19694 16897
rect 20066 16830 20078 16882
rect 20130 16830 20142 16882
rect 20402 16857 20414 16909
rect 20466 16857 20478 16909
rect 20750 16882 20802 16894
rect 22318 16882 22370 16894
rect 23314 16886 23326 16938
rect 23378 16886 23390 16938
rect 23662 16882 23714 16894
rect 21746 16830 21758 16882
rect 21810 16830 21822 16882
rect 22978 16830 22990 16882
rect 23042 16830 23054 16882
rect 13134 16818 13186 16830
rect 18510 16818 18562 16830
rect 20750 16818 20802 16830
rect 22318 16818 22370 16830
rect 23662 16818 23714 16830
rect 9762 16718 9774 16770
rect 9826 16718 9838 16770
rect 19730 16718 19742 16770
rect 19794 16718 19806 16770
rect 4902 16658 4954 16670
rect 4902 16594 4954 16606
rect 8878 16658 8930 16670
rect 8878 16594 8930 16606
rect 1344 16490 24640 16524
rect 1344 16438 4126 16490
rect 4178 16438 4230 16490
rect 4282 16438 4334 16490
rect 4386 16438 9950 16490
rect 10002 16438 10054 16490
rect 10106 16438 10158 16490
rect 10210 16438 15774 16490
rect 15826 16438 15878 16490
rect 15930 16438 15982 16490
rect 16034 16438 21598 16490
rect 21650 16438 21702 16490
rect 21754 16438 21806 16490
rect 21858 16438 24640 16490
rect 1344 16404 24640 16438
rect 8654 16322 8706 16334
rect 8654 16258 8706 16270
rect 14534 16322 14586 16334
rect 14534 16258 14586 16270
rect 17390 16322 17442 16334
rect 17390 16258 17442 16270
rect 4958 16210 5010 16222
rect 3154 16158 3166 16210
rect 3218 16158 3230 16210
rect 3882 16158 3894 16210
rect 3946 16158 3958 16210
rect 4958 16146 5010 16158
rect 6526 16210 6578 16222
rect 6526 16146 6578 16158
rect 3502 16098 3554 16110
rect 2818 16046 2830 16098
rect 2882 16046 2894 16098
rect 3042 16031 3054 16083
rect 3106 16031 3118 16083
rect 3502 16034 3554 16046
rect 3614 16098 3666 16110
rect 3614 16034 3666 16046
rect 4286 16098 4338 16110
rect 6862 16098 6914 16110
rect 4386 16046 4398 16098
rect 4450 16046 4462 16098
rect 6290 16046 6302 16098
rect 6354 16046 6366 16098
rect 4286 16034 4338 16046
rect 4552 15990 4564 16042
rect 4616 15990 4628 16042
rect 6626 15990 6638 16042
rect 6690 15990 6702 16042
rect 6862 16034 6914 16046
rect 7198 16098 7250 16110
rect 7198 16034 7250 16046
rect 7646 16098 7698 16110
rect 7646 16034 7698 16046
rect 7982 16098 8034 16110
rect 7982 16034 8034 16046
rect 8990 16098 9042 16110
rect 8990 16034 9042 16046
rect 9326 16098 9378 16110
rect 9326 16034 9378 16046
rect 11230 16098 11282 16110
rect 11230 16034 11282 16046
rect 11454 16098 11506 16110
rect 11454 16034 11506 16046
rect 12014 16098 12066 16110
rect 12014 16034 12066 16046
rect 12238 16098 12290 16110
rect 19294 16098 19346 16110
rect 12506 16046 12518 16098
rect 12570 16046 12582 16098
rect 14354 16046 14366 16098
rect 14418 16046 14430 16098
rect 12238 16034 12290 16046
rect 16706 16018 16718 16070
rect 16770 16018 16782 16070
rect 19294 16034 19346 16046
rect 19630 16098 19682 16110
rect 19630 16034 19682 16046
rect 20078 16098 20130 16110
rect 23662 16098 23714 16110
rect 20626 16046 20638 16098
rect 20690 16046 20702 16098
rect 22773 16046 22785 16098
rect 22837 16046 22849 16098
rect 20078 16034 20130 16046
rect 20402 15990 20414 16042
rect 20466 15990 20478 16042
rect 23662 16034 23714 16046
rect 22542 15986 22594 15998
rect 11722 15934 11734 15986
rect 11786 15934 11798 15986
rect 9662 15874 9714 15886
rect 20066 15878 20078 15930
rect 20130 15878 20142 15930
rect 22542 15922 22594 15934
rect 24278 15986 24330 15998
rect 24278 15922 24330 15934
rect 9662 15810 9714 15822
rect 1344 15706 24800 15740
rect 1344 15654 7038 15706
rect 7090 15654 7142 15706
rect 7194 15654 7246 15706
rect 7298 15654 12862 15706
rect 12914 15654 12966 15706
rect 13018 15654 13070 15706
rect 13122 15654 18686 15706
rect 18738 15654 18790 15706
rect 18842 15654 18894 15706
rect 18946 15654 24510 15706
rect 24562 15654 24614 15706
rect 24666 15654 24718 15706
rect 24770 15654 24800 15706
rect 1344 15620 24800 15654
rect 8710 15538 8762 15550
rect 8710 15474 8762 15486
rect 12350 15538 12402 15550
rect 12350 15474 12402 15486
rect 21242 15374 21254 15426
rect 21306 15374 21318 15426
rect 3826 15318 3838 15370
rect 3890 15318 3902 15370
rect 4498 15318 4510 15370
rect 4562 15318 4574 15370
rect 5618 15318 5630 15370
rect 5682 15318 5694 15370
rect 6290 15318 6302 15370
rect 6354 15318 6366 15370
rect 7256 15314 7308 15326
rect 7534 15314 7586 15326
rect 7410 15262 7422 15314
rect 7474 15262 7486 15314
rect 7256 15250 7308 15262
rect 7534 15250 7586 15262
rect 7758 15314 7810 15326
rect 7758 15250 7810 15262
rect 7982 15314 8034 15326
rect 10054 15314 10106 15326
rect 10334 15314 10386 15326
rect 8866 15262 8878 15314
rect 8930 15262 8942 15314
rect 10210 15262 10222 15314
rect 10274 15262 10286 15314
rect 7982 15250 8034 15262
rect 10054 15250 10106 15262
rect 10334 15250 10386 15262
rect 10558 15314 10610 15326
rect 10558 15250 10610 15262
rect 12014 15314 12066 15326
rect 14298 15278 14310 15330
rect 14362 15278 14374 15330
rect 14466 15318 14478 15370
rect 14530 15318 14542 15370
rect 14690 15318 14702 15370
rect 14754 15318 14766 15370
rect 14952 15278 14964 15330
rect 15016 15278 15028 15330
rect 15206 15314 15258 15326
rect 12014 15250 12066 15262
rect 15206 15250 15258 15262
rect 15486 15314 15538 15326
rect 15486 15250 15538 15262
rect 17278 15314 17330 15326
rect 17278 15250 17330 15262
rect 19966 15314 20018 15326
rect 20514 15277 20526 15329
rect 20578 15277 20590 15329
rect 21534 15314 21586 15326
rect 20850 15262 20862 15314
rect 20914 15262 20926 15314
rect 19966 15250 20018 15262
rect 21534 15250 21586 15262
rect 21758 15314 21810 15326
rect 23146 15318 23158 15370
rect 23210 15318 23222 15370
rect 23550 15314 23602 15326
rect 22866 15262 22878 15314
rect 22930 15262 22942 15314
rect 21758 15250 21810 15262
rect 23550 15250 23602 15262
rect 23886 15314 23938 15326
rect 23886 15250 23938 15262
rect 9662 15202 9714 15214
rect 3938 15094 3950 15146
rect 4002 15094 4014 15146
rect 9662 15138 9714 15150
rect 10894 15202 10946 15214
rect 18050 15150 18062 15202
rect 18114 15150 18126 15202
rect 20402 15150 20414 15202
rect 20466 15150 20478 15202
rect 22978 15150 22990 15202
rect 23042 15150 23054 15202
rect 10894 15138 10946 15150
rect 6862 15090 6914 15102
rect 15822 15090 15874 15102
rect 8250 15038 8262 15090
rect 8314 15038 8326 15090
rect 6862 15026 6914 15038
rect 15822 15026 15874 15038
rect 1344 14922 24640 14956
rect 1344 14870 4126 14922
rect 4178 14870 4230 14922
rect 4282 14870 4334 14922
rect 4386 14870 9950 14922
rect 10002 14870 10054 14922
rect 10106 14870 10158 14922
rect 10210 14870 15774 14922
rect 15826 14870 15878 14922
rect 15930 14870 15982 14922
rect 16034 14870 21598 14922
rect 21650 14870 21702 14922
rect 21754 14870 21806 14922
rect 21858 14870 24640 14922
rect 1344 14836 24640 14870
rect 18174 14754 18226 14766
rect 23102 14754 23154 14766
rect 20346 14702 20358 14754
rect 20410 14702 20422 14754
rect 18174 14690 18226 14702
rect 23102 14690 23154 14702
rect 9438 14642 9490 14654
rect 4274 14590 4286 14642
rect 4338 14590 4350 14642
rect 9438 14578 9490 14590
rect 13638 14586 13690 14598
rect 17042 14590 17054 14642
rect 17106 14590 17118 14642
rect 1598 14530 1650 14542
rect 5798 14530 5850 14542
rect 9774 14530 9826 14542
rect 2370 14478 2382 14530
rect 2434 14478 2446 14530
rect 4722 14478 4734 14530
rect 4786 14478 4798 14530
rect 6514 14478 6526 14530
rect 6578 14478 6590 14530
rect 1598 14466 1650 14478
rect 5798 14466 5850 14478
rect 8754 14450 8766 14502
rect 8818 14450 8830 14502
rect 9090 14478 9102 14530
rect 9154 14478 9166 14530
rect 9550 14491 9602 14503
rect 9774 14466 9826 14478
rect 10110 14530 10162 14542
rect 10110 14466 10162 14478
rect 13022 14530 13074 14542
rect 13638 14522 13690 14534
rect 14142 14530 14194 14542
rect 13022 14466 13074 14478
rect 14142 14466 14194 14478
rect 14384 14530 14436 14542
rect 14384 14466 14436 14478
rect 17838 14530 17890 14542
rect 17838 14466 17890 14478
rect 18510 14530 18562 14542
rect 18510 14466 18562 14478
rect 20638 14530 20690 14542
rect 20638 14466 20690 14478
rect 20862 14530 20914 14542
rect 21982 14530 22034 14542
rect 21298 14478 21310 14530
rect 21362 14478 21374 14530
rect 20862 14466 20914 14478
rect 9550 14427 9602 14439
rect 13470 14418 13522 14430
rect 13470 14354 13522 14366
rect 15150 14418 15202 14430
rect 21578 14422 21590 14474
rect 21642 14422 21654 14474
rect 21982 14466 22034 14478
rect 24222 14530 24274 14542
rect 23333 14422 23345 14474
rect 23397 14422 23409 14474
rect 24222 14466 24274 14478
rect 15150 14354 15202 14366
rect 4902 14306 4954 14318
rect 4902 14242 4954 14254
rect 12686 14306 12738 14318
rect 21410 14310 21422 14362
rect 21474 14310 21486 14362
rect 12686 14242 12738 14254
rect 1344 14138 24800 14172
rect 1344 14086 7038 14138
rect 7090 14086 7142 14138
rect 7194 14086 7246 14138
rect 7298 14086 12862 14138
rect 12914 14086 12966 14138
rect 13018 14086 13070 14138
rect 13122 14086 18686 14138
rect 18738 14086 18790 14138
rect 18842 14086 18894 14138
rect 18946 14086 24510 14138
rect 24562 14086 24614 14138
rect 24666 14086 24718 14138
rect 24770 14086 24800 14138
rect 1344 14052 24800 14086
rect 2662 13970 2714 13982
rect 2662 13906 2714 13918
rect 14926 13970 14978 13982
rect 14926 13906 14978 13918
rect 23606 13970 23658 13982
rect 23606 13906 23658 13918
rect 24110 13970 24162 13982
rect 24110 13906 24162 13918
rect 14254 13858 14306 13870
rect 4510 13746 4562 13758
rect 2818 13694 2830 13746
rect 2882 13694 2894 13746
rect 4510 13682 4562 13694
rect 4846 13746 4898 13758
rect 4846 13682 4898 13694
rect 6862 13746 6914 13758
rect 7242 13750 7254 13802
rect 7306 13750 7318 13802
rect 8128 13784 8180 13796
rect 14254 13794 14306 13806
rect 7870 13746 7922 13758
rect 7410 13694 7422 13746
rect 7474 13694 7486 13746
rect 7970 13694 7982 13746
rect 8034 13694 8046 13746
rect 8128 13720 8180 13732
rect 11398 13746 11450 13758
rect 6862 13682 6914 13694
rect 7870 13682 7922 13694
rect 11398 13682 11450 13694
rect 11566 13746 11618 13758
rect 14590 13746 14642 13758
rect 12338 13694 12350 13746
rect 12402 13694 12414 13746
rect 11566 13682 11618 13694
rect 14590 13682 14642 13694
rect 18174 13746 18226 13758
rect 18174 13682 18226 13694
rect 20862 13746 20914 13758
rect 21298 13694 21310 13746
rect 21362 13694 21374 13746
rect 21634 13709 21646 13761
rect 21698 13709 21710 13761
rect 22430 13746 22482 13758
rect 22642 13750 22654 13802
rect 22706 13750 22718 13802
rect 23774 13746 23826 13758
rect 23090 13694 23102 13746
rect 23154 13694 23166 13746
rect 20862 13682 20914 13694
rect 22430 13682 22482 13694
rect 23774 13682 23826 13694
rect 7198 13634 7250 13646
rect 7198 13570 7250 13582
rect 10950 13634 11002 13646
rect 22766 13634 22818 13646
rect 18946 13582 18958 13634
rect 19010 13582 19022 13634
rect 21746 13582 21758 13634
rect 21810 13582 21822 13634
rect 10950 13570 11002 13582
rect 22766 13570 22818 13582
rect 8542 13522 8594 13534
rect 8542 13458 8594 13470
rect 1344 13354 24640 13388
rect 1344 13302 4126 13354
rect 4178 13302 4230 13354
rect 4282 13302 4334 13354
rect 4386 13302 9950 13354
rect 10002 13302 10054 13354
rect 10106 13302 10158 13354
rect 10210 13302 15774 13354
rect 15826 13302 15878 13354
rect 15930 13302 15982 13354
rect 16034 13302 21598 13354
rect 21650 13302 21702 13354
rect 21754 13302 21806 13354
rect 21858 13302 24640 13354
rect 1344 13268 24640 13302
rect 19070 13186 19122 13198
rect 5630 13130 5682 13142
rect 4902 13074 4954 13086
rect 4274 13022 4286 13074
rect 4338 13022 4350 13074
rect 19070 13122 19122 13134
rect 22318 13186 22370 13198
rect 22318 13122 22370 13134
rect 5630 13066 5682 13078
rect 9046 13074 9098 13086
rect 4902 13010 4954 13022
rect 15362 13022 15374 13074
rect 15426 13022 15438 13074
rect 9046 13010 9098 13022
rect 1598 12962 1650 12974
rect 6862 12962 6914 12974
rect 2370 12910 2382 12962
rect 2434 12910 2446 12962
rect 5730 12910 5742 12962
rect 5794 12910 5806 12962
rect 5954 12910 5966 12962
rect 6018 12910 6030 12962
rect 1598 12898 1650 12910
rect 6862 12898 6914 12910
rect 7086 12962 7138 12974
rect 7086 12898 7138 12910
rect 7254 12962 7306 12974
rect 7534 12962 7586 12974
rect 7410 12910 7422 12962
rect 7474 12910 7486 12962
rect 7254 12898 7306 12910
rect 7534 12898 7586 12910
rect 8654 12962 8706 12974
rect 8654 12898 8706 12910
rect 9214 12962 9266 12974
rect 14590 12962 14642 12974
rect 18062 12962 18114 12974
rect 9986 12910 9998 12962
rect 10050 12910 10062 12962
rect 17266 12910 17278 12962
rect 17330 12910 17342 12962
rect 9214 12898 9266 12910
rect 7814 12850 7866 12862
rect 7814 12786 7866 12798
rect 11902 12850 11954 12862
rect 11902 12786 11954 12798
rect 13918 12850 13970 12862
rect 14074 12854 14086 12906
rect 14138 12854 14150 12906
rect 14590 12898 14642 12910
rect 18062 12898 18114 12910
rect 19406 12962 19458 12974
rect 19406 12898 19458 12910
rect 23438 12962 23490 12974
rect 13918 12786 13970 12798
rect 14832 12850 14884 12862
rect 22549 12854 22561 12906
rect 22613 12854 22625 12906
rect 23438 12898 23490 12910
rect 23998 12962 24050 12974
rect 23998 12898 24050 12910
rect 24334 12962 24386 12974
rect 24334 12898 24386 12910
rect 14832 12786 14884 12798
rect 6526 12738 6578 12750
rect 6526 12674 6578 12686
rect 8318 12738 8370 12750
rect 8318 12674 8370 12686
rect 1344 12570 24800 12604
rect 1344 12518 7038 12570
rect 7090 12518 7142 12570
rect 7194 12518 7246 12570
rect 7298 12518 12862 12570
rect 12914 12518 12966 12570
rect 13018 12518 13070 12570
rect 13122 12518 18686 12570
rect 18738 12518 18790 12570
rect 18842 12518 18894 12570
rect 18946 12518 24510 12570
rect 24562 12518 24614 12570
rect 24666 12518 24718 12570
rect 24770 12518 24800 12570
rect 1344 12484 24800 12518
rect 3838 12402 3890 12414
rect 3838 12338 3890 12350
rect 13358 12402 13410 12414
rect 13358 12338 13410 12350
rect 15934 12402 15986 12414
rect 15934 12338 15986 12350
rect 24054 12346 24106 12358
rect 7646 12290 7698 12302
rect 6784 12216 6836 12228
rect 7646 12226 7698 12238
rect 21086 12290 21138 12302
rect 22082 12294 22094 12346
rect 22146 12294 22158 12346
rect 22866 12294 22878 12346
rect 22930 12294 22942 12346
rect 24054 12282 24106 12294
rect 4174 12178 4226 12190
rect 4318 12164 4330 12216
rect 4382 12164 4394 12216
rect 5406 12178 5458 12190
rect 5058 12126 5070 12178
rect 5122 12126 5134 12178
rect 4174 12114 4226 12126
rect 5406 12114 5458 12126
rect 5630 12178 5682 12190
rect 5630 12114 5682 12126
rect 6526 12178 6578 12190
rect 6626 12126 6638 12178
rect 6690 12126 6702 12178
rect 7802 12182 7814 12234
rect 7866 12182 7878 12234
rect 6784 12152 6836 12164
rect 8318 12178 8370 12190
rect 6526 12114 6578 12126
rect 8318 12114 8370 12126
rect 8560 12178 8612 12190
rect 8560 12114 8612 12126
rect 9438 12178 9490 12190
rect 9438 12114 9490 12126
rect 9662 12178 9714 12190
rect 9662 12114 9714 12126
rect 10334 12178 10386 12190
rect 10490 12182 10502 12234
rect 10554 12182 10566 12234
rect 21086 12226 21138 12238
rect 10334 12114 10386 12126
rect 11006 12178 11058 12190
rect 11778 12153 11790 12205
rect 11842 12153 11854 12205
rect 14366 12178 14418 12190
rect 11006 12114 11058 12126
rect 14366 12114 14418 12126
rect 15598 12178 15650 12190
rect 15598 12114 15650 12126
rect 18398 12178 18450 12190
rect 21970 12182 21982 12234
rect 22034 12182 22046 12234
rect 22206 12178 22258 12190
rect 23202 12182 23214 12234
rect 23266 12182 23278 12234
rect 23438 12178 23490 12190
rect 21522 12126 21534 12178
rect 21586 12126 21598 12178
rect 22866 12126 22878 12178
rect 22930 12126 22942 12178
rect 23874 12126 23886 12178
rect 23938 12126 23950 12178
rect 18398 12114 18450 12126
rect 22206 12114 22258 12126
rect 23438 12114 23490 12126
rect 7198 12066 7250 12078
rect 5182 12010 5234 12022
rect 19170 12014 19182 12066
rect 19234 12014 19246 12066
rect 7198 12002 7250 12014
rect 5182 11946 5234 11958
rect 11248 11954 11300 11966
rect 5898 11902 5910 11954
rect 5962 11902 5974 11954
rect 9930 11902 9942 11954
rect 9994 11902 10006 11954
rect 11248 11890 11300 11902
rect 14702 11954 14754 11966
rect 14702 11890 14754 11902
rect 1344 11786 24640 11820
rect 1344 11734 4126 11786
rect 4178 11734 4230 11786
rect 4282 11734 4334 11786
rect 4386 11734 9950 11786
rect 10002 11734 10054 11786
rect 10106 11734 10158 11786
rect 10210 11734 15774 11786
rect 15826 11734 15878 11786
rect 15930 11734 15982 11786
rect 16034 11734 21598 11786
rect 21650 11734 21702 11786
rect 21754 11734 21806 11786
rect 21858 11734 24640 11786
rect 1344 11700 24640 11734
rect 19518 11618 19570 11630
rect 7522 11510 7534 11562
rect 7586 11510 7598 11562
rect 19518 11554 19570 11566
rect 24278 11506 24330 11518
rect 5798 11450 5850 11462
rect 22530 11454 22542 11506
rect 22594 11454 22606 11506
rect 23314 11454 23326 11506
rect 23378 11454 23390 11506
rect 5630 11394 5682 11406
rect 3938 11309 3950 11361
rect 4002 11309 4014 11361
rect 4274 11305 4286 11357
rect 4338 11305 4350 11357
rect 4610 11286 4622 11338
rect 4674 11286 4686 11338
rect 4920 11309 4932 11361
rect 4984 11309 4996 11361
rect 24278 11442 24330 11454
rect 5798 11386 5850 11398
rect 6078 11394 6130 11406
rect 9662 11394 9714 11406
rect 5954 11342 5966 11394
rect 6018 11342 6030 11394
rect 7410 11342 7422 11394
rect 7474 11342 7486 11394
rect 7746 11342 7758 11394
rect 7810 11342 7822 11394
rect 5630 11330 5682 11342
rect 6078 11330 6130 11342
rect 9662 11330 9714 11342
rect 9998 11394 10050 11406
rect 9998 11330 10050 11342
rect 10110 11394 10162 11406
rect 15262 11394 15314 11406
rect 18734 11394 18786 11406
rect 10882 11342 10894 11394
rect 10946 11342 10958 11394
rect 17938 11342 17950 11394
rect 18002 11342 18014 11394
rect 10110 11330 10162 11342
rect 5070 11282 5122 11294
rect 5070 11218 5122 11230
rect 6358 11282 6410 11294
rect 6358 11218 6410 11230
rect 12798 11282 12850 11294
rect 14746 11286 14758 11338
rect 14810 11286 14822 11338
rect 15262 11330 15314 11342
rect 18734 11330 18786 11342
rect 19854 11394 19906 11406
rect 21982 11394 22034 11406
rect 21298 11342 21310 11394
rect 21362 11342 21374 11394
rect 21758 11355 21810 11367
rect 19854 11330 19906 11342
rect 21982 11330 22034 11342
rect 22642 11327 22654 11379
rect 22706 11327 22718 11379
rect 22866 11342 22878 11394
rect 22930 11342 22942 11394
rect 12798 11218 12850 11230
rect 15504 11282 15556 11294
rect 14914 11174 14926 11226
rect 14978 11174 14990 11226
rect 15504 11218 15556 11230
rect 16046 11282 16098 11294
rect 21758 11291 21810 11303
rect 23426 11298 23438 11350
rect 23490 11298 23502 11350
rect 23650 11342 23662 11394
rect 23714 11342 23726 11394
rect 16046 11218 16098 11230
rect 21522 11174 21534 11226
rect 21586 11174 21598 11226
rect 1344 11002 24800 11036
rect 1344 10950 7038 11002
rect 7090 10950 7142 11002
rect 7194 10950 7246 11002
rect 7298 10950 12862 11002
rect 12914 10950 12966 11002
rect 13018 10950 13070 11002
rect 13122 10950 18686 11002
rect 18738 10950 18790 11002
rect 18842 10950 18894 11002
rect 18946 10950 24510 11002
rect 24562 10950 24614 11002
rect 24666 10950 24718 11002
rect 24770 10950 24800 11002
rect 1344 10916 24800 10950
rect 16270 10834 16322 10846
rect 16270 10770 16322 10782
rect 18734 10834 18786 10846
rect 18734 10770 18786 10782
rect 23382 10834 23434 10846
rect 23382 10770 23434 10782
rect 13470 10722 13522 10734
rect 4734 10666 4786 10678
rect 3558 10639 3610 10651
rect 3266 10558 3278 10610
rect 3330 10558 3342 10610
rect 3558 10575 3610 10587
rect 4050 10558 4062 10610
rect 4114 10558 4126 10610
rect 4274 10558 4286 10610
rect 4338 10558 4350 10610
rect 4734 10602 4786 10614
rect 4846 10638 4898 10650
rect 5058 10614 5070 10666
rect 5122 10614 5134 10666
rect 5294 10638 5346 10650
rect 4846 10574 4898 10586
rect 5886 10596 5898 10648
rect 5950 10596 5962 10648
rect 6694 10610 6746 10622
rect 8206 10610 8258 10622
rect 8418 10614 8430 10666
rect 8482 10614 8494 10666
rect 13470 10658 13522 10670
rect 14384 10722 14436 10734
rect 22586 10670 22598 10722
rect 22650 10670 22662 10722
rect 9662 10610 9714 10622
rect 13626 10614 13638 10666
rect 13690 10614 13702 10666
rect 14384 10658 14436 10670
rect 5294 10574 5346 10586
rect 7186 10558 7198 10610
rect 7250 10558 7262 10610
rect 7522 10558 7534 10610
rect 7586 10558 7598 10610
rect 8866 10558 8878 10610
rect 8930 10558 8942 10610
rect 6694 10546 6746 10558
rect 8206 10546 8258 10558
rect 9662 10546 9714 10558
rect 14142 10610 14194 10622
rect 14142 10546 14194 10558
rect 15934 10610 15986 10622
rect 17714 10585 17726 10637
rect 17778 10585 17790 10637
rect 21758 10610 21810 10622
rect 15934 10546 15986 10558
rect 21758 10546 21810 10558
rect 22878 10610 22930 10622
rect 22878 10546 22930 10558
rect 23102 10610 23154 10622
rect 23774 10610 23826 10622
rect 23538 10558 23550 10610
rect 23602 10558 23614 10610
rect 23102 10546 23154 10558
rect 23774 10546 23826 10558
rect 22262 10498 22314 10510
rect 3602 10446 3614 10498
rect 3666 10446 3678 10498
rect 4398 10442 4450 10454
rect 7646 10442 7698 10454
rect 8642 10446 8654 10498
rect 8706 10446 8718 10498
rect 10434 10446 10446 10498
rect 10498 10446 10510 10498
rect 12338 10446 12350 10498
rect 12402 10446 12414 10498
rect 4398 10378 4450 10390
rect 5574 10386 5626 10398
rect 6402 10390 6414 10442
rect 6466 10390 6478 10442
rect 22262 10434 22314 10446
rect 7646 10378 7698 10390
rect 21422 10386 21474 10398
rect 5574 10322 5626 10334
rect 21422 10322 21474 10334
rect 24110 10386 24162 10398
rect 24110 10322 24162 10334
rect 1344 10218 24640 10252
rect 1344 10166 4126 10218
rect 4178 10166 4230 10218
rect 4282 10166 4334 10218
rect 4386 10166 9950 10218
rect 10002 10166 10054 10218
rect 10106 10166 10158 10218
rect 10210 10166 15774 10218
rect 15826 10166 15878 10218
rect 15930 10166 15982 10218
rect 16034 10166 21598 10218
rect 21650 10166 21702 10218
rect 21754 10166 21806 10218
rect 21858 10166 24640 10218
rect 1344 10132 24640 10166
rect 14384 10050 14436 10062
rect 6682 9998 6694 10050
rect 6746 9998 6758 10050
rect 14384 9986 14436 9998
rect 9650 9886 9662 9938
rect 9714 9886 9726 9938
rect 13638 9882 13690 9894
rect 21970 9886 21982 9938
rect 22034 9886 22046 9938
rect 6974 9826 7026 9838
rect 6974 9762 7026 9774
rect 7198 9826 7250 9838
rect 7198 9762 7250 9774
rect 7310 9826 7362 9838
rect 7310 9762 7362 9774
rect 7534 9826 7586 9838
rect 11902 9826 11954 9838
rect 7534 9762 7586 9774
rect 10658 9746 10670 9798
rect 10722 9746 10734 9798
rect 11902 9762 11954 9774
rect 13470 9826 13522 9838
rect 13638 9818 13690 9830
rect 14142 9826 14194 9838
rect 13470 9762 13522 9774
rect 14142 9762 14194 9774
rect 15486 9826 15538 9838
rect 14814 9714 14866 9726
rect 14970 9718 14982 9770
rect 15034 9718 15046 9770
rect 15486 9762 15538 9774
rect 16494 9826 16546 9838
rect 19182 9826 19234 9838
rect 18386 9774 18398 9826
rect 18450 9774 18462 9826
rect 16494 9762 16546 9774
rect 19182 9762 19234 9774
rect 19854 9826 19906 9838
rect 19854 9762 19906 9774
rect 21198 9826 21250 9838
rect 21198 9762 21250 9774
rect 7802 9662 7814 9714
rect 7866 9662 7878 9714
rect 14814 9650 14866 9662
rect 15728 9714 15780 9726
rect 15728 9650 15780 9662
rect 23886 9714 23938 9726
rect 23886 9650 23938 9662
rect 12238 9602 12290 9614
rect 12238 9538 12290 9550
rect 19518 9602 19570 9614
rect 19518 9538 19570 9550
rect 1344 9434 24800 9468
rect 1344 9382 7038 9434
rect 7090 9382 7142 9434
rect 7194 9382 7246 9434
rect 7298 9382 12862 9434
rect 12914 9382 12966 9434
rect 13018 9382 13070 9434
rect 13122 9382 18686 9434
rect 18738 9382 18790 9434
rect 18842 9382 18894 9434
rect 18946 9382 24510 9434
rect 24562 9382 24614 9434
rect 24666 9382 24718 9434
rect 24770 9382 24800 9434
rect 1344 9348 24800 9382
rect 16606 9266 16658 9278
rect 16606 9202 16658 9214
rect 19126 9266 19178 9278
rect 19126 9202 19178 9214
rect 12910 9154 12962 9166
rect 4958 9042 5010 9054
rect 10222 9042 10274 9054
rect 8082 8990 8094 9042
rect 8146 8990 8158 9042
rect 9538 8990 9550 9042
rect 9602 8990 9614 9042
rect 9874 8990 9886 9042
rect 9938 8990 9950 9042
rect 4958 8978 5010 8990
rect 10222 8978 10274 8990
rect 11678 9042 11730 9054
rect 11678 8978 11730 8990
rect 11996 9042 12048 9054
rect 11996 8978 12048 8990
rect 12238 9042 12290 9054
rect 12730 9046 12742 9098
rect 12794 9046 12806 9098
rect 12910 9090 12962 9102
rect 14496 9154 14548 9166
rect 14496 9090 14548 9102
rect 12238 8978 12290 8990
rect 13582 9042 13634 9054
rect 14254 9042 14306 9054
rect 13582 8978 13634 8990
rect 13750 8986 13802 8998
rect 14254 8978 14306 8990
rect 16270 9042 16322 9054
rect 23333 9046 23345 9098
rect 23397 9046 23409 9098
rect 16270 8978 16322 8990
rect 24222 9042 24274 9054
rect 24222 8978 24274 8990
rect 5730 8878 5742 8930
rect 5794 8878 5806 8930
rect 7634 8878 7646 8930
rect 7698 8878 7710 8930
rect 13750 8922 13802 8934
rect 22710 8930 22762 8942
rect 9998 8874 10050 8886
rect 22710 8866 22762 8878
rect 9998 8810 10050 8822
rect 10558 8818 10610 8830
rect 10558 8754 10610 8766
rect 11342 8818 11394 8830
rect 11342 8754 11394 8766
rect 23102 8818 23154 8830
rect 23102 8754 23154 8766
rect 1344 8650 24640 8684
rect 1344 8598 4126 8650
rect 4178 8598 4230 8650
rect 4282 8598 4334 8650
rect 4386 8598 9950 8650
rect 10002 8598 10054 8650
rect 10106 8598 10158 8650
rect 10210 8598 15774 8650
rect 15826 8598 15878 8650
rect 15930 8598 15982 8650
rect 16034 8598 21598 8650
rect 21650 8598 21702 8650
rect 21754 8598 21806 8650
rect 21858 8598 24640 8650
rect 1344 8564 24640 8598
rect 5854 8482 5906 8494
rect 5854 8418 5906 8430
rect 22094 8426 22146 8438
rect 7634 8318 7646 8370
rect 7698 8318 7710 8370
rect 10658 8318 10670 8370
rect 10722 8318 10734 8370
rect 15698 8318 15710 8370
rect 15762 8318 15774 8370
rect 22094 8362 22146 8374
rect 23102 8370 23154 8382
rect 23102 8306 23154 8318
rect 5518 8258 5570 8270
rect 5518 8194 5570 8206
rect 6190 8258 6242 8270
rect 6190 8194 6242 8206
rect 6862 8258 6914 8270
rect 6862 8194 6914 8206
rect 9886 8258 9938 8270
rect 9886 8194 9938 8206
rect 14254 8258 14306 8270
rect 14254 8194 14306 8206
rect 14926 8258 14978 8270
rect 18398 8258 18450 8270
rect 24222 8258 24274 8270
rect 17602 8206 17614 8258
rect 17666 8206 17678 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 9550 8146 9602 8158
rect 9550 8082 9602 8094
rect 12574 8146 12626 8158
rect 14410 8150 14422 8202
rect 14474 8150 14486 8202
rect 14926 8194 14978 8206
rect 18398 8194 18450 8206
rect 19954 8191 19966 8243
rect 20018 8191 20030 8243
rect 22194 8206 22206 8258
rect 22258 8206 22270 8258
rect 22530 8206 22542 8258
rect 22594 8206 22606 8258
rect 12574 8082 12626 8094
rect 15168 8146 15220 8158
rect 23333 8150 23345 8202
rect 23397 8150 23409 8202
rect 24222 8194 24274 8206
rect 15168 8082 15220 8094
rect 6526 8034 6578 8046
rect 19730 8038 19742 8090
rect 19794 8038 19806 8090
rect 6526 7970 6578 7982
rect 1344 7866 24800 7900
rect 1344 7814 7038 7866
rect 7090 7814 7142 7866
rect 7194 7814 7246 7866
rect 7298 7814 12862 7866
rect 12914 7814 12966 7866
rect 13018 7814 13070 7866
rect 13122 7814 18686 7866
rect 18738 7814 18790 7866
rect 18842 7814 18894 7866
rect 18946 7814 24510 7866
rect 24562 7814 24614 7866
rect 24666 7814 24718 7866
rect 24770 7814 24800 7866
rect 1344 7780 24800 7814
rect 16158 7698 16210 7710
rect 16158 7634 16210 7646
rect 24110 7698 24162 7710
rect 24110 7634 24162 7646
rect 11118 7586 11170 7598
rect 11118 7522 11170 7534
rect 13470 7586 13522 7598
rect 13470 7522 13522 7534
rect 14384 7586 14436 7598
rect 5182 7474 5234 7486
rect 8206 7474 8258 7486
rect 5954 7422 5966 7474
rect 6018 7422 6030 7474
rect 11790 7474 11842 7486
rect 13626 7478 13638 7530
rect 13690 7478 13702 7530
rect 14384 7522 14436 7534
rect 21646 7586 21698 7598
rect 21646 7522 21698 7534
rect 5182 7410 5234 7422
rect 8206 7410 8258 7422
rect 11286 7418 11338 7430
rect 11790 7410 11842 7422
rect 14142 7474 14194 7486
rect 14142 7410 14194 7422
rect 15822 7474 15874 7486
rect 18386 7437 18398 7489
rect 18450 7437 18462 7489
rect 18958 7474 19010 7486
rect 22418 7478 22430 7530
rect 22482 7478 22494 7530
rect 22766 7474 22818 7486
rect 18722 7422 18734 7474
rect 18786 7422 18798 7474
rect 19730 7422 19742 7474
rect 19794 7422 19806 7474
rect 22194 7422 22206 7474
rect 22258 7422 22270 7474
rect 15822 7410 15874 7422
rect 18958 7410 19010 7422
rect 22766 7410 22818 7422
rect 23102 7474 23154 7486
rect 23102 7410 23154 7422
rect 23774 7474 23826 7486
rect 23774 7410 23826 7422
rect 7858 7310 7870 7362
rect 7922 7310 7934 7362
rect 11286 7354 11338 7366
rect 22430 7362 22482 7374
rect 18274 7310 18286 7362
rect 18338 7310 18350 7362
rect 22430 7298 22482 7310
rect 8542 7250 8594 7262
rect 8542 7186 8594 7198
rect 12032 7250 12084 7262
rect 12032 7186 12084 7198
rect 1344 7082 24640 7116
rect 1344 7030 4126 7082
rect 4178 7030 4230 7082
rect 4282 7030 4334 7082
rect 4386 7030 9950 7082
rect 10002 7030 10054 7082
rect 10106 7030 10158 7082
rect 10210 7030 15774 7082
rect 15826 7030 15878 7082
rect 15930 7030 15982 7082
rect 16034 7030 21598 7082
rect 21650 7030 21702 7082
rect 21754 7030 21806 7082
rect 21858 7030 24640 7082
rect 1344 6996 24640 7030
rect 22374 6914 22426 6926
rect 22374 6850 22426 6862
rect 23606 6802 23658 6814
rect 8306 6750 8318 6802
rect 8370 6750 8382 6802
rect 13906 6750 13918 6802
rect 13970 6750 13982 6802
rect 15810 6750 15822 6802
rect 15874 6750 15886 6802
rect 17490 6750 17502 6802
rect 17554 6750 17566 6802
rect 23606 6738 23658 6750
rect 7534 6690 7586 6702
rect 7534 6626 7586 6638
rect 10222 6690 10274 6702
rect 10222 6626 10274 6638
rect 11678 6690 11730 6702
rect 11678 6626 11730 6638
rect 11846 6690 11898 6702
rect 11846 6626 11898 6638
rect 12350 6690 12402 6702
rect 12350 6626 12402 6638
rect 16606 6690 16658 6702
rect 16606 6626 16658 6638
rect 16718 6690 16770 6702
rect 20526 6690 20578 6702
rect 19954 6638 19966 6690
rect 20018 6638 20030 6690
rect 16718 6626 16770 6638
rect 12592 6578 12644 6590
rect 12592 6514 12644 6526
rect 19406 6578 19458 6590
rect 20290 6582 20302 6634
rect 20354 6582 20366 6634
rect 20526 6626 20578 6638
rect 21646 6690 21698 6702
rect 21646 6626 21698 6638
rect 22094 6690 22146 6702
rect 21802 6582 21814 6634
rect 21866 6582 21878 6634
rect 22094 6626 22146 6638
rect 23214 6690 23266 6702
rect 23214 6626 23266 6638
rect 24334 6690 24386 6702
rect 24334 6626 24386 6638
rect 19406 6514 19458 6526
rect 21982 6578 22034 6590
rect 19954 6470 19966 6522
rect 20018 6470 20030 6522
rect 21982 6514 22034 6526
rect 22878 6466 22930 6478
rect 22878 6402 22930 6414
rect 23998 6466 24050 6478
rect 23998 6402 24050 6414
rect 1344 6298 24800 6332
rect 1344 6246 7038 6298
rect 7090 6246 7142 6298
rect 7194 6246 7246 6298
rect 7298 6246 12862 6298
rect 12914 6246 12966 6298
rect 13018 6246 13070 6298
rect 13122 6246 18686 6298
rect 18738 6246 18790 6298
rect 18842 6246 18894 6298
rect 18946 6246 24510 6298
rect 24562 6246 24614 6298
rect 24666 6246 24718 6298
rect 24770 6246 24800 6298
rect 1344 6212 24800 6246
rect 14814 6130 14866 6142
rect 14814 6066 14866 6078
rect 12686 6018 12738 6030
rect 11230 5906 11282 5918
rect 11230 5842 11282 5854
rect 11772 5906 11824 5918
rect 11772 5842 11824 5854
rect 12014 5906 12066 5918
rect 12506 5910 12518 5962
rect 12570 5910 12582 5962
rect 12686 5954 12738 5966
rect 13246 6018 13298 6030
rect 13246 5954 13298 5966
rect 18510 6018 18562 6030
rect 20794 5966 20806 6018
rect 20858 5966 20870 6018
rect 13402 5910 13414 5962
rect 13466 5910 13478 5962
rect 18510 5954 18562 5966
rect 12014 5842 12066 5854
rect 13918 5906 13970 5918
rect 13918 5842 13970 5854
rect 14160 5906 14212 5918
rect 14160 5842 14212 5854
rect 14478 5906 14530 5918
rect 18741 5910 18753 5962
rect 18805 5910 18817 5962
rect 14478 5842 14530 5854
rect 19630 5906 19682 5918
rect 20066 5898 20078 5950
rect 20130 5898 20142 5950
rect 21086 5906 21138 5918
rect 20290 5854 20302 5906
rect 20354 5854 20366 5906
rect 19630 5842 19682 5854
rect 21086 5842 21138 5854
rect 21198 5906 21250 5918
rect 21198 5842 21250 5854
rect 21422 5906 21474 5918
rect 22549 5910 22561 5962
rect 22613 5910 22625 5962
rect 21422 5842 21474 5854
rect 23438 5906 23490 5918
rect 23438 5842 23490 5854
rect 24334 5906 24386 5918
rect 24334 5842 24386 5854
rect 21758 5794 21810 5806
rect 19954 5742 19966 5794
rect 20018 5742 20030 5794
rect 21758 5730 21810 5742
rect 10894 5682 10946 5694
rect 10894 5618 10946 5630
rect 22318 5682 22370 5694
rect 22318 5618 22370 5630
rect 23998 5682 24050 5694
rect 23998 5618 24050 5630
rect 1344 5514 24640 5548
rect 1344 5462 4126 5514
rect 4178 5462 4230 5514
rect 4282 5462 4334 5514
rect 4386 5462 9950 5514
rect 10002 5462 10054 5514
rect 10106 5462 10158 5514
rect 10210 5462 15774 5514
rect 15826 5462 15878 5514
rect 15930 5462 15982 5514
rect 16034 5462 21598 5514
rect 21650 5462 21702 5514
rect 21754 5462 21806 5514
rect 21858 5462 24640 5514
rect 1344 5428 24640 5462
rect 23326 5234 23378 5246
rect 10546 5182 10558 5234
rect 10610 5182 10622 5234
rect 12450 5182 12462 5234
rect 12514 5182 12526 5234
rect 20402 5182 20414 5234
rect 20466 5182 20478 5234
rect 23326 5170 23378 5182
rect 9774 5122 9826 5134
rect 9774 5058 9826 5070
rect 19742 5122 19794 5134
rect 21422 5122 21474 5134
rect 20066 5070 20078 5122
rect 20130 5070 20142 5122
rect 19742 5058 19794 5070
rect 20290 5055 20302 5107
rect 20354 5055 20366 5107
rect 21422 5058 21474 5070
rect 22542 5122 22594 5134
rect 23662 5122 23714 5134
rect 22978 5070 22990 5122
rect 23042 5070 23054 5122
rect 22286 5014 22298 5066
rect 22350 5014 22362 5066
rect 22542 5058 22594 5070
rect 23426 5014 23438 5066
rect 23490 5014 23502 5066
rect 23662 5058 23714 5070
rect 23998 5122 24050 5134
rect 23998 5058 24050 5070
rect 19406 4898 19458 4910
rect 19406 4834 19458 4846
rect 1344 4730 24800 4764
rect 1344 4678 7038 4730
rect 7090 4678 7142 4730
rect 7194 4678 7246 4730
rect 7298 4678 12862 4730
rect 12914 4678 12966 4730
rect 13018 4678 13070 4730
rect 13122 4678 18686 4730
rect 18738 4678 18790 4730
rect 18842 4678 18894 4730
rect 18946 4678 24510 4730
rect 24562 4678 24614 4730
rect 24666 4678 24718 4730
rect 24770 4678 24800 4730
rect 1344 4644 24800 4678
rect 20974 4450 21026 4462
rect 20974 4386 21026 4398
rect 23998 4450 24050 4462
rect 23998 4386 24050 4398
rect 18286 4338 18338 4350
rect 21310 4338 21362 4350
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 22082 4286 22094 4338
rect 22146 4286 22158 4338
rect 18286 4274 18338 4286
rect 21310 4274 21362 4286
rect 1344 3946 24640 3980
rect 1344 3894 4126 3946
rect 4178 3894 4230 3946
rect 4282 3894 4334 3946
rect 4386 3894 9950 3946
rect 10002 3894 10054 3946
rect 10106 3894 10158 3946
rect 10210 3894 15774 3946
rect 15826 3894 15878 3946
rect 15930 3894 15982 3946
rect 16034 3894 21598 3946
rect 21650 3894 21702 3946
rect 21754 3894 21806 3946
rect 21858 3894 24640 3946
rect 1344 3860 24640 3894
rect 21870 3778 21922 3790
rect 21870 3714 21922 3726
rect 23438 3778 23490 3790
rect 23438 3714 23490 3726
rect 24054 3666 24106 3678
rect 24054 3602 24106 3614
rect 21534 3554 21586 3566
rect 21534 3490 21586 3502
rect 22318 3554 22370 3566
rect 23182 3502 23194 3554
rect 23246 3502 23258 3554
rect 22318 3490 22370 3502
rect 21366 3442 21418 3454
rect 21366 3378 21418 3390
rect 1344 3162 24800 3196
rect 1344 3110 7038 3162
rect 7090 3110 7142 3162
rect 7194 3110 7246 3162
rect 7298 3110 12862 3162
rect 12914 3110 12966 3162
rect 13018 3110 13070 3162
rect 13122 3110 18686 3162
rect 18738 3110 18790 3162
rect 18842 3110 18894 3162
rect 18946 3110 24510 3162
rect 24562 3110 24614 3162
rect 24666 3110 24718 3162
rect 24770 3110 24800 3162
rect 1344 3076 24800 3110
<< via1 >>
rect 6918 22878 6970 22930
rect 7758 22878 7810 22930
rect 4126 22710 4178 22762
rect 4230 22710 4282 22762
rect 4334 22710 4386 22762
rect 9950 22710 10002 22762
rect 10054 22710 10106 22762
rect 10158 22710 10210 22762
rect 15774 22710 15826 22762
rect 15878 22710 15930 22762
rect 15982 22710 16034 22762
rect 21598 22710 21650 22762
rect 21702 22710 21754 22762
rect 21806 22710 21858 22762
rect 6918 22542 6970 22594
rect 22542 22542 22594 22594
rect 7870 22486 7922 22538
rect 12126 22430 12178 22482
rect 21198 22430 21250 22482
rect 7198 22318 7250 22370
rect 7422 22318 7474 22370
rect 7758 22318 7810 22370
rect 8094 22318 8146 22370
rect 11454 22318 11506 22370
rect 11566 22318 11618 22370
rect 11732 22318 11784 22370
rect 13582 22318 13634 22370
rect 13974 22318 14026 22370
rect 19742 22318 19794 22370
rect 20750 22318 20802 22370
rect 21086 22274 21138 22326
rect 21534 22290 21586 22342
rect 19574 22206 19626 22258
rect 8598 22094 8650 22146
rect 13246 22094 13298 22146
rect 20078 22094 20130 22146
rect 7038 21926 7090 21978
rect 7142 21926 7194 21978
rect 7246 21926 7298 21978
rect 12862 21926 12914 21978
rect 12966 21926 13018 21978
rect 13070 21926 13122 21978
rect 18686 21926 18738 21978
rect 18790 21926 18842 21978
rect 18894 21926 18946 21978
rect 24510 21926 24562 21978
rect 24614 21926 24666 21978
rect 24718 21926 24770 21978
rect 7422 21646 7474 21698
rect 4734 21534 4786 21586
rect 7814 21590 7866 21642
rect 8430 21590 8482 21642
rect 8206 21534 8258 21586
rect 9905 21534 9957 21586
rect 10782 21534 10834 21586
rect 11678 21534 11730 21586
rect 14702 21534 14754 21586
rect 14926 21534 14978 21586
rect 15262 21534 15314 21586
rect 15598 21534 15650 21586
rect 17278 21534 17330 21586
rect 20862 21534 20914 21586
rect 5518 21422 5570 21474
rect 7982 21422 8034 21474
rect 11342 21422 11394 21474
rect 12014 21422 12066 21474
rect 13918 21422 13970 21474
rect 18062 21422 18114 21474
rect 19966 21422 20018 21474
rect 21646 21422 21698 21474
rect 23550 21422 23602 21474
rect 24278 21422 24330 21474
rect 15262 21366 15314 21418
rect 9662 21310 9714 21362
rect 15934 21310 15986 21362
rect 4126 21142 4178 21194
rect 4230 21142 4282 21194
rect 4334 21142 4386 21194
rect 9950 21142 10002 21194
rect 10054 21142 10106 21194
rect 10158 21142 10210 21194
rect 15774 21142 15826 21194
rect 15878 21142 15930 21194
rect 15982 21142 16034 21194
rect 21598 21142 21650 21194
rect 21702 21142 21754 21194
rect 21806 21142 21858 21194
rect 8822 20862 8874 20914
rect 9550 20862 9602 20914
rect 10446 20918 10498 20970
rect 11454 20918 11506 20970
rect 12126 20918 12178 20970
rect 21366 20974 21418 21026
rect 14926 20918 14978 20970
rect 15934 20862 15986 20914
rect 17838 20862 17890 20914
rect 19294 20862 19346 20914
rect 5518 20750 5570 20802
rect 6302 20750 6354 20802
rect 9214 20750 9266 20802
rect 9662 20711 9714 20763
rect 9886 20750 9938 20802
rect 10558 20750 10610 20802
rect 10894 20750 10946 20802
rect 11342 20750 11394 20802
rect 11678 20750 11730 20802
rect 12238 20750 12290 20802
rect 12914 20712 12966 20764
rect 14138 20712 14190 20764
rect 14814 20750 14866 20802
rect 15150 20750 15202 20802
rect 18958 20750 19010 20802
rect 19182 20706 19234 20758
rect 19630 20750 19682 20802
rect 20302 20750 20354 20802
rect 19910 20694 19962 20746
rect 21646 20750 21698 20802
rect 21870 20750 21922 20802
rect 22206 20750 22258 20802
rect 23082 20750 23134 20802
rect 24334 20750 24386 20802
rect 8206 20638 8258 20690
rect 23326 20638 23378 20690
rect 19742 20582 19794 20634
rect 23998 20526 24050 20578
rect 7038 20358 7090 20410
rect 7142 20358 7194 20410
rect 7246 20358 7298 20410
rect 12862 20358 12914 20410
rect 12966 20358 13018 20410
rect 13070 20358 13122 20410
rect 18686 20358 18738 20410
rect 18790 20358 18842 20410
rect 18894 20358 18946 20410
rect 24510 20358 24562 20410
rect 24614 20358 24666 20410
rect 24718 20358 24770 20410
rect 4678 20190 4730 20242
rect 5854 20190 5906 20242
rect 12238 20190 12290 20242
rect 12686 20190 12738 20242
rect 18062 20190 18114 20242
rect 8206 20134 8258 20186
rect 22318 20190 22370 20242
rect 21534 20134 21586 20186
rect 20526 20078 20578 20130
rect 5182 19966 5234 20018
rect 6190 19966 6242 20018
rect 8094 19966 8146 20018
rect 8542 20005 8594 20057
rect 8766 19966 8818 20018
rect 9662 19966 9714 20018
rect 9886 19966 9938 20018
rect 10446 19966 10498 20018
rect 10670 19966 10722 20018
rect 11230 19966 11282 20018
rect 11454 19966 11506 20018
rect 15038 19966 15090 20018
rect 15150 19966 15202 20018
rect 15296 20004 15348 20056
rect 18398 19966 18450 20018
rect 19406 19966 19458 20018
rect 19742 19966 19794 20018
rect 20358 20022 20410 20074
rect 20190 19966 20242 20018
rect 20638 19966 20690 20018
rect 21310 19966 21362 20018
rect 21590 19995 21642 20047
rect 23754 20022 23806 20074
rect 11734 19854 11786 19906
rect 15710 19854 15762 19906
rect 18790 19854 18842 19906
rect 19238 19854 19290 19906
rect 22654 19910 22706 19962
rect 22878 19966 22930 20018
rect 5014 19742 5066 19794
rect 10166 19742 10218 19794
rect 10950 19742 11002 19794
rect 20918 19742 20970 19794
rect 23998 19742 24050 19794
rect 4126 19574 4178 19626
rect 4230 19574 4282 19626
rect 4334 19574 4386 19626
rect 9950 19574 10002 19626
rect 10054 19574 10106 19626
rect 10158 19574 10210 19626
rect 15774 19574 15826 19626
rect 15878 19574 15930 19626
rect 15982 19574 16034 19626
rect 21598 19574 21650 19626
rect 21702 19574 21754 19626
rect 21806 19574 21858 19626
rect 7982 19406 8034 19458
rect 20358 19406 20410 19458
rect 9494 19350 9546 19402
rect 9886 19294 9938 19346
rect 13582 19294 13634 19346
rect 21310 19294 21362 19346
rect 22598 19294 22650 19346
rect 2046 19182 2098 19234
rect 2830 19182 2882 19234
rect 5518 19182 5570 19234
rect 8318 19182 8370 19234
rect 8654 19182 8706 19234
rect 9662 19182 9714 19234
rect 9998 19138 10050 19190
rect 10222 19182 10274 19234
rect 10670 19182 10722 19234
rect 10838 19182 10890 19234
rect 11118 19182 11170 19234
rect 11398 19182 11450 19234
rect 11902 19182 11954 19234
rect 12070 19238 12122 19290
rect 12350 19182 12402 19234
rect 15486 19182 15538 19234
rect 16270 19182 16322 19234
rect 16830 19182 16882 19234
rect 17614 19182 17666 19234
rect 20638 19182 20690 19234
rect 20862 19182 20914 19234
rect 21422 19138 21474 19190
rect 21758 19182 21810 19234
rect 23233 19182 23285 19234
rect 24110 19182 24162 19234
rect 4734 19070 4786 19122
rect 8990 19070 9042 19122
rect 11006 19070 11058 19122
rect 12238 19070 12290 19122
rect 12630 19070 12682 19122
rect 19518 19070 19570 19122
rect 22990 19070 23042 19122
rect 5686 18958 5738 19010
rect 6246 18958 6298 19010
rect 7038 18790 7090 18842
rect 7142 18790 7194 18842
rect 7246 18790 7298 18842
rect 12862 18790 12914 18842
rect 12966 18790 13018 18842
rect 13070 18790 13122 18842
rect 18686 18790 18738 18842
rect 18790 18790 18842 18842
rect 18894 18790 18946 18842
rect 24510 18790 24562 18842
rect 24614 18790 24666 18842
rect 24718 18790 24770 18842
rect 17838 18622 17890 18674
rect 20190 18566 20242 18618
rect 1598 18398 1650 18450
rect 4286 18398 4338 18450
rect 5070 18398 5122 18450
rect 5294 18398 5346 18450
rect 5854 18398 5906 18450
rect 6730 18398 6782 18450
rect 7870 18398 7922 18450
rect 11006 18398 11058 18450
rect 11342 18398 11394 18450
rect 12014 18398 12066 18450
rect 12910 18398 12962 18450
rect 13358 18398 13410 18450
rect 13694 18398 13746 18450
rect 15150 18398 15202 18450
rect 20414 18454 20466 18506
rect 18174 18398 18226 18450
rect 19966 18398 20018 18450
rect 20638 18398 20690 18450
rect 23438 18454 23490 18506
rect 22766 18398 22818 18450
rect 22990 18398 23042 18450
rect 23662 18398 23714 18450
rect 23998 18398 24050 18450
rect 2382 18286 2434 18338
rect 22038 18286 22090 18338
rect 4790 18174 4842 18226
rect 6974 18174 7026 18226
rect 11118 18230 11170 18282
rect 23326 18286 23378 18338
rect 7534 18174 7586 18226
rect 11846 18174 11898 18226
rect 12574 18174 12626 18226
rect 15486 18174 15538 18226
rect 22430 18174 22482 18226
rect 4126 18006 4178 18058
rect 4230 18006 4282 18058
rect 4334 18006 4386 18058
rect 9950 18006 10002 18058
rect 10054 18006 10106 18058
rect 10158 18006 10210 18058
rect 15774 18006 15826 18058
rect 15878 18006 15930 18058
rect 15982 18006 16034 18058
rect 21598 18006 21650 18058
rect 21702 18006 21754 18058
rect 21806 18006 21858 18058
rect 4286 17782 4338 17834
rect 11566 17838 11618 17890
rect 13694 17838 13746 17890
rect 12238 17782 12290 17834
rect 5742 17726 5794 17778
rect 14590 17726 14642 17778
rect 16494 17726 16546 17778
rect 3950 17614 4002 17666
rect 4174 17614 4226 17666
rect 4678 17614 4730 17666
rect 4958 17614 5010 17666
rect 5182 17614 5234 17666
rect 6134 17614 6186 17666
rect 6302 17614 6354 17666
rect 6414 17614 6466 17666
rect 6750 17614 6802 17666
rect 7422 17614 7474 17666
rect 7926 17614 7978 17666
rect 8206 17614 8258 17666
rect 8318 17614 8370 17666
rect 8486 17614 8538 17666
rect 8654 17614 8706 17666
rect 8878 17614 8930 17666
rect 11118 17614 11170 17666
rect 11902 17614 11954 17666
rect 12238 17614 12290 17666
rect 12462 17614 12514 17666
rect 13358 17614 13410 17666
rect 17278 17614 17330 17666
rect 17390 17614 17442 17666
rect 18174 17614 18226 17666
rect 22094 17614 22146 17666
rect 24334 17614 24386 17666
rect 22970 17558 23022 17610
rect 20078 17502 20130 17554
rect 7534 17446 7586 17498
rect 23214 17502 23266 17554
rect 9214 17390 9266 17442
rect 10782 17390 10834 17442
rect 23998 17390 24050 17442
rect 7038 17222 7090 17274
rect 7142 17222 7194 17274
rect 7246 17222 7298 17274
rect 12862 17222 12914 17274
rect 12966 17222 13018 17274
rect 13070 17222 13122 17274
rect 18686 17222 18738 17274
rect 18790 17222 18842 17274
rect 18894 17222 18946 17274
rect 24510 17222 24562 17274
rect 24614 17222 24666 17274
rect 24718 17222 24770 17274
rect 18174 17054 18226 17106
rect 3278 16998 3330 17050
rect 6190 16942 6242 16994
rect 3054 16830 3106 16882
rect 3726 16830 3778 16882
rect 4062 16886 4114 16938
rect 4174 16886 4226 16938
rect 4398 16886 4450 16938
rect 4622 16886 4674 16938
rect 6022 16886 6074 16938
rect 12574 16998 12626 17050
rect 6582 16942 6634 16994
rect 20190 16998 20242 17050
rect 21534 16998 21586 17050
rect 23102 16998 23154 17050
rect 15430 16942 15482 16994
rect 5854 16830 5906 16882
rect 6302 16830 6354 16882
rect 6862 16830 6914 16882
rect 7926 16830 7978 16882
rect 8206 16830 8258 16882
rect 8318 16830 8370 16882
rect 8504 16868 8556 16920
rect 9886 16886 9938 16938
rect 9550 16830 9602 16882
rect 10222 16830 10274 16882
rect 10558 16830 10610 16882
rect 11790 16830 11842 16882
rect 12350 16830 12402 16882
rect 12910 16830 12962 16882
rect 13134 16830 13186 16882
rect 13414 16830 13466 16882
rect 14590 16865 14642 16917
rect 14702 16858 14754 16910
rect 14926 16858 14978 16910
rect 15150 16886 15202 16938
rect 18510 16830 18562 16882
rect 19406 16830 19458 16882
rect 19630 16845 19682 16897
rect 20078 16830 20130 16882
rect 20414 16857 20466 16909
rect 23326 16886 23378 16938
rect 20750 16830 20802 16882
rect 21758 16830 21810 16882
rect 22318 16830 22370 16882
rect 22990 16830 23042 16882
rect 23662 16830 23714 16882
rect 9774 16718 9826 16770
rect 19742 16718 19794 16770
rect 4902 16606 4954 16658
rect 8878 16606 8930 16658
rect 4126 16438 4178 16490
rect 4230 16438 4282 16490
rect 4334 16438 4386 16490
rect 9950 16438 10002 16490
rect 10054 16438 10106 16490
rect 10158 16438 10210 16490
rect 15774 16438 15826 16490
rect 15878 16438 15930 16490
rect 15982 16438 16034 16490
rect 21598 16438 21650 16490
rect 21702 16438 21754 16490
rect 21806 16438 21858 16490
rect 8654 16270 8706 16322
rect 14534 16270 14586 16322
rect 17390 16270 17442 16322
rect 3166 16158 3218 16210
rect 3894 16158 3946 16210
rect 4958 16158 5010 16210
rect 6526 16158 6578 16210
rect 2830 16046 2882 16098
rect 3054 16031 3106 16083
rect 3502 16046 3554 16098
rect 3614 16046 3666 16098
rect 4286 16046 4338 16098
rect 4398 16046 4450 16098
rect 6302 16046 6354 16098
rect 6862 16046 6914 16098
rect 4564 15990 4616 16042
rect 6638 15990 6690 16042
rect 7198 16046 7250 16098
rect 7646 16046 7698 16098
rect 7982 16046 8034 16098
rect 8990 16046 9042 16098
rect 9326 16046 9378 16098
rect 11230 16046 11282 16098
rect 11454 16046 11506 16098
rect 12014 16046 12066 16098
rect 12238 16046 12290 16098
rect 12518 16046 12570 16098
rect 14366 16046 14418 16098
rect 16718 16018 16770 16070
rect 19294 16046 19346 16098
rect 19630 16046 19682 16098
rect 20078 16046 20130 16098
rect 20638 16046 20690 16098
rect 22785 16046 22837 16098
rect 23662 16046 23714 16098
rect 20414 15990 20466 16042
rect 11734 15934 11786 15986
rect 22542 15934 22594 15986
rect 20078 15878 20130 15930
rect 24278 15934 24330 15986
rect 9662 15822 9714 15874
rect 7038 15654 7090 15706
rect 7142 15654 7194 15706
rect 7246 15654 7298 15706
rect 12862 15654 12914 15706
rect 12966 15654 13018 15706
rect 13070 15654 13122 15706
rect 18686 15654 18738 15706
rect 18790 15654 18842 15706
rect 18894 15654 18946 15706
rect 24510 15654 24562 15706
rect 24614 15654 24666 15706
rect 24718 15654 24770 15706
rect 8710 15486 8762 15538
rect 12350 15486 12402 15538
rect 21254 15374 21306 15426
rect 3838 15318 3890 15370
rect 4510 15318 4562 15370
rect 5630 15318 5682 15370
rect 6302 15318 6354 15370
rect 7256 15262 7308 15314
rect 7422 15262 7474 15314
rect 7534 15262 7586 15314
rect 7758 15262 7810 15314
rect 7982 15262 8034 15314
rect 8878 15262 8930 15314
rect 10054 15262 10106 15314
rect 10222 15262 10274 15314
rect 10334 15262 10386 15314
rect 10558 15262 10610 15314
rect 12014 15262 12066 15314
rect 14310 15278 14362 15330
rect 14478 15318 14530 15370
rect 14702 15318 14754 15370
rect 14964 15278 15016 15330
rect 15206 15262 15258 15314
rect 15486 15262 15538 15314
rect 17278 15262 17330 15314
rect 19966 15262 20018 15314
rect 20526 15277 20578 15329
rect 20862 15262 20914 15314
rect 21534 15262 21586 15314
rect 23158 15318 23210 15370
rect 21758 15262 21810 15314
rect 22878 15262 22930 15314
rect 23550 15262 23602 15314
rect 23886 15262 23938 15314
rect 9662 15150 9714 15202
rect 3950 15094 4002 15146
rect 10894 15150 10946 15202
rect 18062 15150 18114 15202
rect 20414 15150 20466 15202
rect 22990 15150 23042 15202
rect 6862 15038 6914 15090
rect 8262 15038 8314 15090
rect 15822 15038 15874 15090
rect 4126 14870 4178 14922
rect 4230 14870 4282 14922
rect 4334 14870 4386 14922
rect 9950 14870 10002 14922
rect 10054 14870 10106 14922
rect 10158 14870 10210 14922
rect 15774 14870 15826 14922
rect 15878 14870 15930 14922
rect 15982 14870 16034 14922
rect 21598 14870 21650 14922
rect 21702 14870 21754 14922
rect 21806 14870 21858 14922
rect 18174 14702 18226 14754
rect 20358 14702 20410 14754
rect 23102 14702 23154 14754
rect 4286 14590 4338 14642
rect 9438 14590 9490 14642
rect 17054 14590 17106 14642
rect 1598 14478 1650 14530
rect 2382 14478 2434 14530
rect 4734 14478 4786 14530
rect 5798 14478 5850 14530
rect 6526 14478 6578 14530
rect 8766 14450 8818 14502
rect 9102 14478 9154 14530
rect 9550 14439 9602 14491
rect 9774 14478 9826 14530
rect 10110 14478 10162 14530
rect 13022 14478 13074 14530
rect 13638 14534 13690 14586
rect 14142 14478 14194 14530
rect 14384 14478 14436 14530
rect 17838 14478 17890 14530
rect 18510 14478 18562 14530
rect 20638 14478 20690 14530
rect 20862 14478 20914 14530
rect 21310 14478 21362 14530
rect 21982 14478 22034 14530
rect 13470 14366 13522 14418
rect 21590 14422 21642 14474
rect 24222 14478 24274 14530
rect 23345 14422 23397 14474
rect 15150 14366 15202 14418
rect 4902 14254 4954 14306
rect 21422 14310 21474 14362
rect 12686 14254 12738 14306
rect 7038 14086 7090 14138
rect 7142 14086 7194 14138
rect 7246 14086 7298 14138
rect 12862 14086 12914 14138
rect 12966 14086 13018 14138
rect 13070 14086 13122 14138
rect 18686 14086 18738 14138
rect 18790 14086 18842 14138
rect 18894 14086 18946 14138
rect 24510 14086 24562 14138
rect 24614 14086 24666 14138
rect 24718 14086 24770 14138
rect 2662 13918 2714 13970
rect 14926 13918 14978 13970
rect 23606 13918 23658 13970
rect 24110 13918 24162 13970
rect 14254 13806 14306 13858
rect 2830 13694 2882 13746
rect 4510 13694 4562 13746
rect 4846 13694 4898 13746
rect 7254 13750 7306 13802
rect 6862 13694 6914 13746
rect 7422 13694 7474 13746
rect 7870 13694 7922 13746
rect 7982 13694 8034 13746
rect 8128 13732 8180 13784
rect 11398 13694 11450 13746
rect 11566 13694 11618 13746
rect 12350 13694 12402 13746
rect 14590 13694 14642 13746
rect 18174 13694 18226 13746
rect 20862 13694 20914 13746
rect 21310 13694 21362 13746
rect 21646 13709 21698 13761
rect 22654 13750 22706 13802
rect 22430 13694 22482 13746
rect 23102 13694 23154 13746
rect 23774 13694 23826 13746
rect 7198 13582 7250 13634
rect 10950 13582 11002 13634
rect 18958 13582 19010 13634
rect 21758 13582 21810 13634
rect 22766 13582 22818 13634
rect 8542 13470 8594 13522
rect 4126 13302 4178 13354
rect 4230 13302 4282 13354
rect 4334 13302 4386 13354
rect 9950 13302 10002 13354
rect 10054 13302 10106 13354
rect 10158 13302 10210 13354
rect 15774 13302 15826 13354
rect 15878 13302 15930 13354
rect 15982 13302 16034 13354
rect 21598 13302 21650 13354
rect 21702 13302 21754 13354
rect 21806 13302 21858 13354
rect 4286 13022 4338 13074
rect 4902 13022 4954 13074
rect 5630 13078 5682 13130
rect 19070 13134 19122 13186
rect 22318 13134 22370 13186
rect 9046 13022 9098 13074
rect 15374 13022 15426 13074
rect 1598 12910 1650 12962
rect 2382 12910 2434 12962
rect 5742 12910 5794 12962
rect 5966 12910 6018 12962
rect 6862 12910 6914 12962
rect 7086 12910 7138 12962
rect 7254 12910 7306 12962
rect 7422 12910 7474 12962
rect 7534 12910 7586 12962
rect 8654 12910 8706 12962
rect 9214 12910 9266 12962
rect 9998 12910 10050 12962
rect 14590 12910 14642 12962
rect 17278 12910 17330 12962
rect 18062 12910 18114 12962
rect 7814 12798 7866 12850
rect 11902 12798 11954 12850
rect 14086 12854 14138 12906
rect 19406 12910 19458 12962
rect 23438 12910 23490 12962
rect 13918 12798 13970 12850
rect 22561 12854 22613 12906
rect 23998 12910 24050 12962
rect 24334 12910 24386 12962
rect 14832 12798 14884 12850
rect 6526 12686 6578 12738
rect 8318 12686 8370 12738
rect 7038 12518 7090 12570
rect 7142 12518 7194 12570
rect 7246 12518 7298 12570
rect 12862 12518 12914 12570
rect 12966 12518 13018 12570
rect 13070 12518 13122 12570
rect 18686 12518 18738 12570
rect 18790 12518 18842 12570
rect 18894 12518 18946 12570
rect 24510 12518 24562 12570
rect 24614 12518 24666 12570
rect 24718 12518 24770 12570
rect 3838 12350 3890 12402
rect 13358 12350 13410 12402
rect 15934 12350 15986 12402
rect 7646 12238 7698 12290
rect 22094 12294 22146 12346
rect 22878 12294 22930 12346
rect 24054 12294 24106 12346
rect 21086 12238 21138 12290
rect 4174 12126 4226 12178
rect 4330 12164 4382 12216
rect 5070 12126 5122 12178
rect 5406 12126 5458 12178
rect 5630 12126 5682 12178
rect 6526 12126 6578 12178
rect 6638 12126 6690 12178
rect 6784 12164 6836 12216
rect 7814 12182 7866 12234
rect 8318 12126 8370 12178
rect 8560 12126 8612 12178
rect 9438 12126 9490 12178
rect 9662 12126 9714 12178
rect 10502 12182 10554 12234
rect 10334 12126 10386 12178
rect 11006 12126 11058 12178
rect 11790 12153 11842 12205
rect 14366 12126 14418 12178
rect 15598 12126 15650 12178
rect 21982 12182 22034 12234
rect 23214 12182 23266 12234
rect 18398 12126 18450 12178
rect 21534 12126 21586 12178
rect 22206 12126 22258 12178
rect 22878 12126 22930 12178
rect 23438 12126 23490 12178
rect 23886 12126 23938 12178
rect 5182 11958 5234 12010
rect 7198 12014 7250 12066
rect 19182 12014 19234 12066
rect 5910 11902 5962 11954
rect 9942 11902 9994 11954
rect 11248 11902 11300 11954
rect 14702 11902 14754 11954
rect 4126 11734 4178 11786
rect 4230 11734 4282 11786
rect 4334 11734 4386 11786
rect 9950 11734 10002 11786
rect 10054 11734 10106 11786
rect 10158 11734 10210 11786
rect 15774 11734 15826 11786
rect 15878 11734 15930 11786
rect 15982 11734 16034 11786
rect 21598 11734 21650 11786
rect 21702 11734 21754 11786
rect 21806 11734 21858 11786
rect 19518 11566 19570 11618
rect 7534 11510 7586 11562
rect 22542 11454 22594 11506
rect 23326 11454 23378 11506
rect 24278 11454 24330 11506
rect 3950 11309 4002 11361
rect 4286 11305 4338 11357
rect 4622 11286 4674 11338
rect 4932 11309 4984 11361
rect 5630 11342 5682 11394
rect 5798 11398 5850 11450
rect 5966 11342 6018 11394
rect 6078 11342 6130 11394
rect 7422 11342 7474 11394
rect 7758 11342 7810 11394
rect 9662 11342 9714 11394
rect 9998 11342 10050 11394
rect 10110 11342 10162 11394
rect 10894 11342 10946 11394
rect 15262 11342 15314 11394
rect 17950 11342 18002 11394
rect 18734 11342 18786 11394
rect 5070 11230 5122 11282
rect 6358 11230 6410 11282
rect 14758 11286 14810 11338
rect 19854 11342 19906 11394
rect 21310 11342 21362 11394
rect 21758 11303 21810 11355
rect 21982 11342 22034 11394
rect 22654 11327 22706 11379
rect 22878 11342 22930 11394
rect 12798 11230 12850 11282
rect 15504 11230 15556 11282
rect 14926 11174 14978 11226
rect 23438 11298 23490 11350
rect 23662 11342 23714 11394
rect 16046 11230 16098 11282
rect 21534 11174 21586 11226
rect 7038 10950 7090 11002
rect 7142 10950 7194 11002
rect 7246 10950 7298 11002
rect 12862 10950 12914 11002
rect 12966 10950 13018 11002
rect 13070 10950 13122 11002
rect 18686 10950 18738 11002
rect 18790 10950 18842 11002
rect 18894 10950 18946 11002
rect 24510 10950 24562 11002
rect 24614 10950 24666 11002
rect 24718 10950 24770 11002
rect 16270 10782 16322 10834
rect 18734 10782 18786 10834
rect 23382 10782 23434 10834
rect 13470 10670 13522 10722
rect 3278 10558 3330 10610
rect 3558 10587 3610 10639
rect 4734 10614 4786 10666
rect 4062 10558 4114 10610
rect 4286 10558 4338 10610
rect 4846 10586 4898 10638
rect 5070 10614 5122 10666
rect 5294 10586 5346 10638
rect 5898 10596 5950 10648
rect 8430 10614 8482 10666
rect 14384 10670 14436 10722
rect 22598 10670 22650 10722
rect 13638 10614 13690 10666
rect 6694 10558 6746 10610
rect 7198 10558 7250 10610
rect 7534 10558 7586 10610
rect 8206 10558 8258 10610
rect 8878 10558 8930 10610
rect 9662 10558 9714 10610
rect 14142 10558 14194 10610
rect 15934 10558 15986 10610
rect 17726 10585 17778 10637
rect 21758 10558 21810 10610
rect 22878 10558 22930 10610
rect 23102 10558 23154 10610
rect 23550 10558 23602 10610
rect 23774 10558 23826 10610
rect 3614 10446 3666 10498
rect 8654 10446 8706 10498
rect 10446 10446 10498 10498
rect 12350 10446 12402 10498
rect 22262 10446 22314 10498
rect 4398 10390 4450 10442
rect 6414 10390 6466 10442
rect 7646 10390 7698 10442
rect 5574 10334 5626 10386
rect 21422 10334 21474 10386
rect 24110 10334 24162 10386
rect 4126 10166 4178 10218
rect 4230 10166 4282 10218
rect 4334 10166 4386 10218
rect 9950 10166 10002 10218
rect 10054 10166 10106 10218
rect 10158 10166 10210 10218
rect 15774 10166 15826 10218
rect 15878 10166 15930 10218
rect 15982 10166 16034 10218
rect 21598 10166 21650 10218
rect 21702 10166 21754 10218
rect 21806 10166 21858 10218
rect 6694 9998 6746 10050
rect 14384 9998 14436 10050
rect 9662 9886 9714 9938
rect 21982 9886 22034 9938
rect 6974 9774 7026 9826
rect 7198 9774 7250 9826
rect 7310 9774 7362 9826
rect 7534 9774 7586 9826
rect 10670 9746 10722 9798
rect 11902 9774 11954 9826
rect 13470 9774 13522 9826
rect 13638 9830 13690 9882
rect 14142 9774 14194 9826
rect 15486 9774 15538 9826
rect 14982 9718 15034 9770
rect 16494 9774 16546 9826
rect 18398 9774 18450 9826
rect 19182 9774 19234 9826
rect 19854 9774 19906 9826
rect 21198 9774 21250 9826
rect 7814 9662 7866 9714
rect 14814 9662 14866 9714
rect 15728 9662 15780 9714
rect 23886 9662 23938 9714
rect 12238 9550 12290 9602
rect 19518 9550 19570 9602
rect 7038 9382 7090 9434
rect 7142 9382 7194 9434
rect 7246 9382 7298 9434
rect 12862 9382 12914 9434
rect 12966 9382 13018 9434
rect 13070 9382 13122 9434
rect 18686 9382 18738 9434
rect 18790 9382 18842 9434
rect 18894 9382 18946 9434
rect 24510 9382 24562 9434
rect 24614 9382 24666 9434
rect 24718 9382 24770 9434
rect 16606 9214 16658 9266
rect 19126 9214 19178 9266
rect 12910 9102 12962 9154
rect 4958 8990 5010 9042
rect 8094 8990 8146 9042
rect 9550 8990 9602 9042
rect 9886 8990 9938 9042
rect 10222 8990 10274 9042
rect 11678 8990 11730 9042
rect 11996 8990 12048 9042
rect 12742 9046 12794 9098
rect 14496 9102 14548 9154
rect 12238 8990 12290 9042
rect 13582 8990 13634 9042
rect 13750 8934 13802 8986
rect 14254 8990 14306 9042
rect 23345 9046 23397 9098
rect 16270 8990 16322 9042
rect 24222 8990 24274 9042
rect 5742 8878 5794 8930
rect 7646 8878 7698 8930
rect 9998 8822 10050 8874
rect 22710 8878 22762 8930
rect 10558 8766 10610 8818
rect 11342 8766 11394 8818
rect 23102 8766 23154 8818
rect 4126 8598 4178 8650
rect 4230 8598 4282 8650
rect 4334 8598 4386 8650
rect 9950 8598 10002 8650
rect 10054 8598 10106 8650
rect 10158 8598 10210 8650
rect 15774 8598 15826 8650
rect 15878 8598 15930 8650
rect 15982 8598 16034 8650
rect 21598 8598 21650 8650
rect 21702 8598 21754 8650
rect 21806 8598 21858 8650
rect 5854 8430 5906 8482
rect 22094 8374 22146 8426
rect 7646 8318 7698 8370
rect 10670 8318 10722 8370
rect 15710 8318 15762 8370
rect 23102 8318 23154 8370
rect 5518 8206 5570 8258
rect 6190 8206 6242 8258
rect 6862 8206 6914 8258
rect 9886 8206 9938 8258
rect 14254 8206 14306 8258
rect 14926 8206 14978 8258
rect 17614 8206 17666 8258
rect 18398 8206 18450 8258
rect 19742 8206 19794 8258
rect 9550 8094 9602 8146
rect 14422 8150 14474 8202
rect 19966 8191 20018 8243
rect 22206 8206 22258 8258
rect 22542 8206 22594 8258
rect 24222 8206 24274 8258
rect 12574 8094 12626 8146
rect 23345 8150 23397 8202
rect 15168 8094 15220 8146
rect 19742 8038 19794 8090
rect 6526 7982 6578 8034
rect 7038 7814 7090 7866
rect 7142 7814 7194 7866
rect 7246 7814 7298 7866
rect 12862 7814 12914 7866
rect 12966 7814 13018 7866
rect 13070 7814 13122 7866
rect 18686 7814 18738 7866
rect 18790 7814 18842 7866
rect 18894 7814 18946 7866
rect 24510 7814 24562 7866
rect 24614 7814 24666 7866
rect 24718 7814 24770 7866
rect 16158 7646 16210 7698
rect 24110 7646 24162 7698
rect 11118 7534 11170 7586
rect 13470 7534 13522 7586
rect 14384 7534 14436 7586
rect 5182 7422 5234 7474
rect 5966 7422 6018 7474
rect 8206 7422 8258 7474
rect 13638 7478 13690 7530
rect 21646 7534 21698 7586
rect 11286 7366 11338 7418
rect 11790 7422 11842 7474
rect 14142 7422 14194 7474
rect 15822 7422 15874 7474
rect 18398 7437 18450 7489
rect 22430 7478 22482 7530
rect 18734 7422 18786 7474
rect 18958 7422 19010 7474
rect 19742 7422 19794 7474
rect 22206 7422 22258 7474
rect 22766 7422 22818 7474
rect 23102 7422 23154 7474
rect 23774 7422 23826 7474
rect 7870 7310 7922 7362
rect 18286 7310 18338 7362
rect 22430 7310 22482 7362
rect 8542 7198 8594 7250
rect 12032 7198 12084 7250
rect 4126 7030 4178 7082
rect 4230 7030 4282 7082
rect 4334 7030 4386 7082
rect 9950 7030 10002 7082
rect 10054 7030 10106 7082
rect 10158 7030 10210 7082
rect 15774 7030 15826 7082
rect 15878 7030 15930 7082
rect 15982 7030 16034 7082
rect 21598 7030 21650 7082
rect 21702 7030 21754 7082
rect 21806 7030 21858 7082
rect 22374 6862 22426 6914
rect 8318 6750 8370 6802
rect 13918 6750 13970 6802
rect 15822 6750 15874 6802
rect 17502 6750 17554 6802
rect 23606 6750 23658 6802
rect 7534 6638 7586 6690
rect 10222 6638 10274 6690
rect 11678 6638 11730 6690
rect 11846 6638 11898 6690
rect 12350 6638 12402 6690
rect 16606 6638 16658 6690
rect 16718 6638 16770 6690
rect 19966 6638 20018 6690
rect 20526 6638 20578 6690
rect 12592 6526 12644 6578
rect 20302 6582 20354 6634
rect 21646 6638 21698 6690
rect 22094 6638 22146 6690
rect 21814 6582 21866 6634
rect 23214 6638 23266 6690
rect 24334 6638 24386 6690
rect 19406 6526 19458 6578
rect 21982 6526 22034 6578
rect 19966 6470 20018 6522
rect 22878 6414 22930 6466
rect 23998 6414 24050 6466
rect 7038 6246 7090 6298
rect 7142 6246 7194 6298
rect 7246 6246 7298 6298
rect 12862 6246 12914 6298
rect 12966 6246 13018 6298
rect 13070 6246 13122 6298
rect 18686 6246 18738 6298
rect 18790 6246 18842 6298
rect 18894 6246 18946 6298
rect 24510 6246 24562 6298
rect 24614 6246 24666 6298
rect 24718 6246 24770 6298
rect 14814 6078 14866 6130
rect 12686 5966 12738 6018
rect 11230 5854 11282 5906
rect 11772 5854 11824 5906
rect 12518 5910 12570 5962
rect 13246 5966 13298 6018
rect 18510 5966 18562 6018
rect 20806 5966 20858 6018
rect 13414 5910 13466 5962
rect 12014 5854 12066 5906
rect 13918 5854 13970 5906
rect 14160 5854 14212 5906
rect 18753 5910 18805 5962
rect 14478 5854 14530 5906
rect 19630 5854 19682 5906
rect 20078 5898 20130 5950
rect 20302 5854 20354 5906
rect 21086 5854 21138 5906
rect 21198 5854 21250 5906
rect 22561 5910 22613 5962
rect 21422 5854 21474 5906
rect 23438 5854 23490 5906
rect 24334 5854 24386 5906
rect 19966 5742 20018 5794
rect 21758 5742 21810 5794
rect 10894 5630 10946 5682
rect 22318 5630 22370 5682
rect 23998 5630 24050 5682
rect 4126 5462 4178 5514
rect 4230 5462 4282 5514
rect 4334 5462 4386 5514
rect 9950 5462 10002 5514
rect 10054 5462 10106 5514
rect 10158 5462 10210 5514
rect 15774 5462 15826 5514
rect 15878 5462 15930 5514
rect 15982 5462 16034 5514
rect 21598 5462 21650 5514
rect 21702 5462 21754 5514
rect 21806 5462 21858 5514
rect 10558 5182 10610 5234
rect 12462 5182 12514 5234
rect 20414 5182 20466 5234
rect 23326 5182 23378 5234
rect 9774 5070 9826 5122
rect 19742 5070 19794 5122
rect 20078 5070 20130 5122
rect 20302 5055 20354 5107
rect 21422 5070 21474 5122
rect 22542 5070 22594 5122
rect 22990 5070 23042 5122
rect 23662 5070 23714 5122
rect 22298 5014 22350 5066
rect 23438 5014 23490 5066
rect 23998 5070 24050 5122
rect 19406 4846 19458 4898
rect 7038 4678 7090 4730
rect 7142 4678 7194 4730
rect 7246 4678 7298 4730
rect 12862 4678 12914 4730
rect 12966 4678 13018 4730
rect 13070 4678 13122 4730
rect 18686 4678 18738 4730
rect 18790 4678 18842 4730
rect 18894 4678 18946 4730
rect 24510 4678 24562 4730
rect 24614 4678 24666 4730
rect 24718 4678 24770 4730
rect 20974 4398 21026 4450
rect 23998 4398 24050 4450
rect 18286 4286 18338 4338
rect 19070 4286 19122 4338
rect 21310 4286 21362 4338
rect 22094 4286 22146 4338
rect 4126 3894 4178 3946
rect 4230 3894 4282 3946
rect 4334 3894 4386 3946
rect 9950 3894 10002 3946
rect 10054 3894 10106 3946
rect 10158 3894 10210 3946
rect 15774 3894 15826 3946
rect 15878 3894 15930 3946
rect 15982 3894 16034 3946
rect 21598 3894 21650 3946
rect 21702 3894 21754 3946
rect 21806 3894 21858 3946
rect 21870 3726 21922 3778
rect 23438 3726 23490 3778
rect 24054 3614 24106 3666
rect 21534 3502 21586 3554
rect 22318 3502 22370 3554
rect 23194 3502 23246 3554
rect 21366 3390 21418 3442
rect 7038 3110 7090 3162
rect 7142 3110 7194 3162
rect 7246 3110 7298 3162
rect 12862 3110 12914 3162
rect 12966 3110 13018 3162
rect 13070 3110 13122 3162
rect 18686 3110 18738 3162
rect 18790 3110 18842 3162
rect 18894 3110 18946 3162
rect 24510 3110 24562 3162
rect 24614 3110 24666 3162
rect 24718 3110 24770 3162
<< metal2 >>
rect 4256 25200 4368 26000
rect 12768 25200 12880 26000
rect 21280 25200 21392 26000
rect 4284 22932 4340 25200
rect 4284 22876 4564 22932
rect 4124 22764 4388 22774
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4124 22698 4388 22708
rect 4124 21196 4388 21206
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4124 21130 4388 21140
rect 4124 19628 4388 19638
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4124 19562 4388 19572
rect 2044 19234 2100 19246
rect 2044 19182 2046 19234
rect 2098 19182 2100 19234
rect 2044 18564 2100 19182
rect 2828 19234 2884 19246
rect 2828 19182 2830 19234
rect 2882 19182 2884 19234
rect 2828 18676 2884 19182
rect 2828 18610 2884 18620
rect 1596 18508 2100 18564
rect 1596 18450 1652 18508
rect 1596 18398 1598 18450
rect 1650 18398 1652 18450
rect 1596 14530 1652 18398
rect 4284 18452 4340 18462
rect 4284 18358 4340 18396
rect 2380 18338 2436 18350
rect 2380 18286 2382 18338
rect 2434 18286 2436 18338
rect 2380 16884 2436 18286
rect 4124 18060 4388 18070
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4124 17994 4388 18004
rect 4284 17834 4340 17846
rect 4284 17782 4286 17834
rect 4338 17782 4340 17834
rect 3948 17666 4004 17678
rect 3948 17614 3950 17666
rect 4002 17614 4004 17666
rect 3724 17108 3780 17118
rect 3276 17050 3332 17062
rect 3276 16998 3278 17050
rect 3330 16998 3332 17050
rect 3276 16996 3332 16998
rect 3276 16930 3332 16940
rect 3052 16884 3108 16894
rect 2380 16818 2436 16828
rect 2940 16882 3108 16884
rect 2940 16830 3054 16882
rect 3106 16830 3108 16882
rect 2940 16828 3108 16830
rect 2828 16100 2884 16110
rect 2940 16100 2996 16828
rect 3052 16818 3108 16828
rect 3388 16884 3444 16894
rect 2884 16044 2996 16100
rect 3052 16212 3108 16222
rect 3052 16083 3108 16156
rect 2828 16006 2884 16044
rect 3052 16031 3054 16083
rect 3106 16031 3108 16083
rect 3052 16019 3108 16031
rect 3164 16210 3220 16222
rect 3164 16158 3166 16210
rect 3218 16158 3220 16210
rect 3164 15764 3220 16158
rect 3164 15698 3220 15708
rect 3388 14868 3444 16828
rect 3724 16882 3780 17052
rect 3948 16996 4004 17614
rect 4172 17668 4228 17678
rect 4060 16996 4116 17006
rect 3948 16940 4060 16996
rect 3724 16830 3726 16882
rect 3778 16830 3780 16882
rect 4060 16938 4116 16940
rect 4060 16886 4062 16938
rect 4114 16886 4116 16938
rect 4060 16874 4116 16886
rect 4172 16938 4228 17612
rect 4284 17332 4340 17782
rect 4284 17266 4340 17276
rect 4172 16886 4174 16938
rect 4226 16886 4228 16938
rect 4172 16874 4228 16886
rect 4396 16996 4452 17006
rect 4396 16938 4452 16940
rect 4396 16886 4398 16938
rect 4450 16886 4452 16938
rect 3612 16772 3668 16782
rect 3612 16212 3668 16716
rect 3500 16100 3556 16110
rect 3500 16006 3556 16044
rect 3612 16098 3668 16156
rect 3612 16046 3614 16098
rect 3666 16046 3668 16098
rect 3612 16034 3668 16046
rect 3388 14812 3556 14868
rect 1596 14478 1598 14530
rect 1650 14478 1652 14530
rect 1596 13524 1652 14478
rect 2380 14532 2436 14542
rect 2380 14530 2716 14532
rect 2380 14478 2382 14530
rect 2434 14478 2716 14530
rect 2380 14476 2716 14478
rect 2380 14466 2436 14476
rect 2660 13970 2716 14476
rect 3500 14308 3556 14812
rect 3500 14242 3556 14252
rect 2660 13918 2662 13970
rect 2714 13918 2716 13970
rect 2660 13906 2716 13918
rect 2828 13748 2884 13758
rect 2828 13654 2884 13692
rect 1596 12962 1652 13468
rect 3724 13076 3780 16830
rect 4396 16660 4452 16886
rect 4508 16772 4564 22876
rect 6916 22930 6972 22942
rect 6916 22878 6918 22930
rect 6970 22878 6972 22930
rect 6916 22594 6972 22878
rect 6916 22542 6918 22594
rect 6970 22542 6972 22594
rect 6916 22530 6972 22542
rect 7756 22930 7812 22942
rect 7756 22878 7758 22930
rect 7810 22878 7812 22930
rect 7196 22370 7252 22382
rect 7196 22318 7198 22370
rect 7250 22318 7252 22370
rect 7196 22148 7252 22318
rect 7196 22082 7252 22092
rect 7420 22370 7476 22382
rect 7420 22318 7422 22370
rect 7474 22318 7476 22370
rect 7036 21980 7300 21990
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7036 21914 7300 21924
rect 7420 21698 7476 22318
rect 7756 22370 7812 22878
rect 9948 22764 10212 22774
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 9948 22698 10212 22708
rect 7756 22318 7758 22370
rect 7810 22318 7812 22370
rect 7756 22306 7812 22318
rect 7868 22538 7924 22550
rect 7868 22486 7870 22538
rect 7922 22486 7924 22538
rect 7420 21646 7422 21698
rect 7474 21646 7476 21698
rect 7868 21654 7924 22486
rect 11340 22540 11786 22596
rect 4732 21586 4788 21598
rect 4732 21534 4734 21586
rect 4786 21534 4788 21586
rect 4732 20282 4788 21534
rect 7420 21588 7476 21646
rect 7812 21642 7924 21654
rect 7812 21590 7814 21642
rect 7866 21590 7924 21642
rect 7812 21588 7924 21590
rect 8092 22370 8148 22382
rect 8092 22318 8094 22370
rect 8146 22318 8148 22370
rect 7812 21578 7868 21588
rect 7420 21522 7476 21532
rect 5516 21476 5572 21486
rect 5516 21382 5572 21420
rect 7980 21476 8036 21486
rect 7980 21382 8036 21420
rect 8092 21140 8148 22318
rect 10108 22372 10164 22382
rect 8428 22148 8484 22158
rect 8428 21642 8484 22092
rect 8596 22148 8652 22158
rect 9324 22148 9380 22158
rect 8596 22146 8820 22148
rect 8596 22094 8598 22146
rect 8650 22094 8820 22146
rect 8596 22092 8820 22094
rect 8596 22082 8652 22092
rect 7980 21084 8148 21140
rect 8204 21588 8260 21598
rect 8428 21590 8430 21642
rect 8482 21590 8484 21642
rect 8428 21578 8484 21590
rect 7980 20916 8036 21084
rect 8204 20916 8260 21532
rect 4676 20244 4788 20282
rect 4732 20188 4788 20244
rect 5516 20802 5572 20814
rect 6300 20804 6356 20814
rect 5516 20750 5518 20802
rect 5570 20750 5572 20802
rect 5516 20244 5572 20750
rect 4676 20178 4732 20188
rect 5516 20178 5572 20188
rect 5852 20802 6356 20804
rect 5852 20750 6302 20802
rect 6354 20750 6356 20802
rect 5852 20748 6356 20750
rect 5852 20242 5908 20748
rect 6300 20738 6356 20748
rect 7036 20412 7300 20422
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7036 20346 7300 20356
rect 5852 20190 5854 20242
rect 5906 20190 5908 20242
rect 5852 20178 5908 20190
rect 6300 20244 6356 20254
rect 5180 20018 5236 20030
rect 5180 19966 5182 20018
rect 5234 19966 5236 20018
rect 5012 19794 5068 19806
rect 5012 19742 5014 19794
rect 5066 19742 5068 19794
rect 4732 19122 4788 19134
rect 5012 19124 5068 19742
rect 4732 19070 4734 19122
rect 4786 19070 4788 19122
rect 4732 18900 4788 19070
rect 4732 18834 4788 18844
rect 4956 19068 5068 19124
rect 4788 18228 4844 18238
rect 4788 18226 4900 18228
rect 4788 18174 4790 18226
rect 4842 18174 4900 18226
rect 4788 18162 4900 18174
rect 4676 17668 4732 17678
rect 4676 17574 4732 17612
rect 4620 17108 4676 17118
rect 4620 16938 4676 17052
rect 4620 16886 4622 16938
rect 4674 16886 4676 16938
rect 4620 16874 4676 16886
rect 4844 16884 4900 18162
rect 4956 17666 5012 19068
rect 5068 18900 5124 18910
rect 5180 18900 5236 19966
rect 6188 20018 6244 20030
rect 6188 19966 6190 20018
rect 6242 19966 6244 20018
rect 6188 19908 6244 19966
rect 6188 19842 6244 19852
rect 5516 19236 5572 19246
rect 5124 18844 5236 18900
rect 5292 19234 5572 19236
rect 5292 19182 5518 19234
rect 5570 19182 5572 19234
rect 5292 19180 5572 19182
rect 5068 18450 5124 18844
rect 5068 18398 5070 18450
rect 5122 18398 5124 18450
rect 5068 18340 5124 18398
rect 5068 18274 5124 18284
rect 5292 18452 5348 19180
rect 5516 19170 5572 19180
rect 6300 19022 6356 20188
rect 7980 19458 8036 20860
rect 8092 20860 8260 20916
rect 8764 20926 8820 22092
rect 8764 20914 8876 20926
rect 8764 20862 8822 20914
rect 8874 20862 8876 20914
rect 8092 20804 8148 20860
rect 8092 20018 8148 20748
rect 8764 20850 8876 20862
rect 8204 20692 8260 20702
rect 8204 20690 8372 20692
rect 8204 20638 8206 20690
rect 8258 20638 8372 20690
rect 8204 20636 8372 20638
rect 8204 20626 8260 20636
rect 8092 19966 8094 20018
rect 8146 19966 8148 20018
rect 8092 19954 8148 19966
rect 8204 20186 8260 20198
rect 8204 20134 8206 20186
rect 8258 20134 8260 20186
rect 8204 19908 8260 20134
rect 8316 20132 8372 20636
rect 8764 20244 8820 20850
rect 9212 20804 9268 20814
rect 9212 20710 9268 20748
rect 8764 20178 8820 20188
rect 8988 20580 9044 20590
rect 8316 20076 8596 20132
rect 8540 20057 8596 20076
rect 8540 20005 8542 20057
rect 8594 20005 8596 20057
rect 8204 19852 8484 19908
rect 7980 19406 7982 19458
rect 8034 19406 8036 19458
rect 7980 19394 8036 19406
rect 8316 19236 8372 19246
rect 5684 19012 5740 19022
rect 5684 19010 5908 19012
rect 5684 18958 5686 19010
rect 5738 18958 5908 19010
rect 5684 18956 5908 18958
rect 5684 18946 5740 18956
rect 5852 18452 5908 18956
rect 6244 19010 6356 19022
rect 6244 18958 6246 19010
rect 6298 18958 6356 19010
rect 6244 18956 6356 18958
rect 8092 19234 8372 19236
rect 8092 19182 8318 19234
rect 8370 19182 8372 19234
rect 8092 19180 8372 19182
rect 6244 18788 6300 18956
rect 7036 18844 7300 18854
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 6244 18732 6580 18788
rect 7036 18778 7300 18788
rect 6524 18676 6580 18732
rect 6524 18620 6916 18676
rect 4956 17614 4958 17666
rect 5010 17614 5012 17666
rect 4956 17556 5012 17614
rect 5180 17668 5236 17678
rect 5292 17668 5348 18396
rect 5628 18450 5908 18452
rect 5628 18398 5854 18450
rect 5906 18398 5908 18450
rect 5628 18396 5908 18398
rect 5628 18004 5684 18396
rect 5852 18386 5908 18396
rect 6728 18450 6784 18462
rect 6728 18398 6730 18450
rect 6782 18398 6784 18450
rect 6728 18340 6784 18398
rect 6728 18274 6784 18284
rect 6524 18004 6580 18014
rect 5628 17948 6188 18004
rect 5180 17666 5348 17668
rect 5180 17614 5182 17666
rect 5234 17614 5348 17666
rect 5180 17612 5348 17614
rect 5740 17778 5796 17790
rect 5740 17726 5742 17778
rect 5794 17726 5796 17778
rect 5180 17602 5236 17612
rect 4956 17490 5012 17500
rect 5068 17108 5124 17118
rect 4956 16884 5012 16894
rect 4844 16828 4956 16884
rect 4956 16818 5012 16828
rect 4508 16716 4788 16772
rect 3948 16604 4452 16660
rect 3948 16222 4004 16604
rect 4124 16492 4388 16502
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4124 16426 4388 16436
rect 3892 16210 4004 16222
rect 3892 16158 3894 16210
rect 3946 16158 4004 16210
rect 3892 16146 4004 16158
rect 3836 15764 3892 15774
rect 3836 15370 3892 15708
rect 3836 15318 3838 15370
rect 3890 15318 3892 15370
rect 3948 15428 4004 16146
rect 4396 16212 4452 16222
rect 4284 16098 4340 16110
rect 4284 16046 4286 16098
rect 4338 16046 4340 16098
rect 4284 15876 4340 16046
rect 4396 16098 4452 16156
rect 4396 16046 4398 16098
rect 4450 16046 4452 16098
rect 4396 16034 4452 16046
rect 4562 16100 4618 16120
rect 4562 16042 4618 16044
rect 4562 15990 4564 16042
rect 4616 15990 4618 16042
rect 4562 15988 4618 15990
rect 4508 15932 4618 15988
rect 4508 15876 4564 15932
rect 4732 15876 4788 16716
rect 4900 16660 4956 16670
rect 5068 16660 5124 17052
rect 4900 16658 5124 16660
rect 4900 16606 4902 16658
rect 4954 16606 5124 16658
rect 4900 16604 5124 16606
rect 4900 16594 4956 16604
rect 4284 15810 4340 15820
rect 4396 15820 4564 15876
rect 4620 15820 4788 15876
rect 4956 16210 5012 16222
rect 4956 16158 4958 16210
rect 5010 16158 5012 16210
rect 3948 15362 4004 15372
rect 3836 15306 3892 15318
rect 4396 15204 4452 15820
rect 4508 15428 4564 15438
rect 4508 15370 4564 15372
rect 4508 15318 4510 15370
rect 4562 15318 4564 15370
rect 4508 15306 4564 15318
rect 3724 13010 3780 13020
rect 3948 15146 4004 15158
rect 4396 15148 4564 15204
rect 3948 15094 3950 15146
rect 4002 15094 4004 15146
rect 1596 12910 1598 12962
rect 1650 12910 1652 12962
rect 1596 12898 1652 12910
rect 2380 12964 2436 12974
rect 2380 12870 2436 12908
rect 3836 12964 3892 12974
rect 3836 12402 3892 12908
rect 3948 12740 4004 15094
rect 4124 14924 4388 14934
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4124 14858 4388 14868
rect 4284 14644 4340 14654
rect 4508 14644 4564 15148
rect 4284 14642 4564 14644
rect 4284 14590 4286 14642
rect 4338 14590 4564 14642
rect 4284 14588 4564 14590
rect 4284 14578 4340 14588
rect 4508 13748 4564 13758
rect 4124 13356 4388 13366
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4124 13290 4388 13300
rect 4284 13076 4340 13086
rect 4284 12982 4340 13020
rect 4284 12740 4340 12750
rect 3948 12684 4284 12740
rect 4340 12684 4384 12740
rect 4284 12646 4384 12684
rect 3836 12350 3838 12402
rect 3890 12350 3892 12402
rect 3276 12292 3332 12302
rect 3276 10610 3332 12236
rect 3836 12292 3892 12350
rect 3836 12226 3892 12236
rect 4328 12216 4384 12646
rect 4172 12180 4228 12190
rect 4328 12164 4330 12216
rect 4382 12164 4384 12216
rect 4328 12152 4384 12164
rect 4172 12086 4228 12124
rect 4124 11788 4388 11798
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4124 11722 4388 11732
rect 4508 11620 4564 13692
rect 4620 13636 4676 15820
rect 4732 15092 4788 15102
rect 4732 14530 4788 15036
rect 4732 14478 4734 14530
rect 4786 14478 4788 14530
rect 4732 14466 4788 14478
rect 4956 14532 5012 16158
rect 5628 15988 5684 15998
rect 5628 15370 5684 15932
rect 5628 15318 5630 15370
rect 5682 15318 5684 15370
rect 5740 15428 5796 17726
rect 6132 17666 6188 17948
rect 6132 17614 6134 17666
rect 6186 17614 6188 17666
rect 6132 17602 6188 17614
rect 6300 17668 6356 17678
rect 6020 17444 6076 17454
rect 6300 17444 6356 17612
rect 5852 17220 5908 17230
rect 5852 16882 5908 17164
rect 5852 16830 5854 16882
rect 5906 16830 5908 16882
rect 6020 16938 6076 17388
rect 6020 16886 6022 16938
rect 6074 16886 6076 16938
rect 6188 17388 6356 17444
rect 6412 17666 6468 17678
rect 6412 17614 6414 17666
rect 6466 17614 6468 17666
rect 6412 17444 6468 17614
rect 6188 16994 6244 17388
rect 6412 17378 6468 17388
rect 6412 17220 6468 17230
rect 6524 17220 6580 17948
rect 6468 17164 6580 17220
rect 6748 17666 6804 17678
rect 6748 17614 6750 17666
rect 6802 17614 6804 17666
rect 6188 16942 6190 16994
rect 6242 16942 6244 16994
rect 6188 16930 6244 16942
rect 6300 16996 6356 17006
rect 6020 16874 6076 16886
rect 6300 16882 6356 16940
rect 5852 16818 5908 16830
rect 6300 16830 6302 16882
rect 6354 16830 6356 16882
rect 6300 16818 6356 16830
rect 6412 16772 6468 17164
rect 6580 16996 6636 17006
rect 6748 16996 6804 17614
rect 6580 16994 6804 16996
rect 6580 16942 6582 16994
rect 6634 16942 6804 16994
rect 6580 16940 6804 16942
rect 6580 16930 6636 16940
rect 6860 16884 6916 18620
rect 7868 18450 7924 18462
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 6972 18228 7028 18238
rect 6972 18226 7364 18228
rect 6972 18174 6974 18226
rect 7026 18174 7364 18226
rect 6972 18172 7364 18174
rect 6972 18162 7028 18172
rect 7308 17444 7364 18172
rect 7532 18226 7588 18238
rect 7532 18174 7534 18226
rect 7586 18174 7588 18226
rect 7532 17892 7588 18174
rect 7532 17826 7588 17836
rect 7868 17892 7924 18398
rect 7868 17826 7924 17836
rect 8092 18228 8148 19180
rect 8316 19170 8372 19180
rect 7420 17668 7476 17678
rect 7924 17668 7980 17678
rect 7420 17666 7980 17668
rect 7420 17614 7422 17666
rect 7474 17614 7926 17666
rect 7978 17614 7980 17666
rect 7420 17612 7980 17614
rect 7420 17602 7476 17612
rect 7924 17602 7980 17612
rect 7532 17498 7588 17510
rect 7532 17446 7534 17498
rect 7586 17446 7588 17498
rect 7308 17388 7476 17444
rect 7036 17276 7300 17286
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7036 17210 7300 17220
rect 7420 17108 7476 17388
rect 6860 16790 6916 16828
rect 7196 17052 7476 17108
rect 7532 17108 7588 17446
rect 8092 17332 8148 18172
rect 8428 18116 8484 19852
rect 8540 19236 8596 20005
rect 8764 20020 8820 20030
rect 8988 20020 9044 20524
rect 8764 20018 9044 20020
rect 8764 19966 8766 20018
rect 8818 19966 9044 20018
rect 8764 19964 9044 19966
rect 9212 20020 9268 20030
rect 8764 19954 8820 19964
rect 8652 19236 8708 19246
rect 8540 19234 8708 19236
rect 8540 19182 8654 19234
rect 8706 19182 8708 19234
rect 8540 19180 8708 19182
rect 8652 19170 8708 19180
rect 8988 19124 9044 19134
rect 8988 19030 9044 19068
rect 9212 19124 9268 19964
rect 9212 19058 9268 19068
rect 9324 19012 9380 22092
rect 9903 21588 9959 21598
rect 9548 21586 9959 21588
rect 9548 21534 9905 21586
rect 9957 21534 9959 21586
rect 9548 21532 9959 21534
rect 9548 20914 9604 21532
rect 9903 21522 9959 21532
rect 10108 21476 10164 22316
rect 11340 21812 11396 22540
rect 11452 22370 11508 22382
rect 11452 22318 11454 22370
rect 11506 22318 11508 22370
rect 11452 21924 11508 22318
rect 11564 22372 11620 22382
rect 11564 22278 11620 22316
rect 11730 22370 11786 22540
rect 12124 22484 12180 22494
rect 11730 22318 11732 22370
rect 11784 22318 11786 22370
rect 11730 22306 11786 22318
rect 11900 22482 12180 22484
rect 11900 22430 12126 22482
rect 12178 22430 12180 22482
rect 11900 22428 12180 22430
rect 11900 22036 11956 22428
rect 12124 22418 12180 22428
rect 12796 22372 12852 25200
rect 15772 22764 16036 22774
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 15772 22698 16036 22708
rect 21308 22596 21364 25200
rect 22876 24052 22932 24062
rect 21596 22764 21860 22774
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21596 22698 21860 22708
rect 21308 22530 21364 22540
rect 22540 22596 22596 22606
rect 22540 22502 22596 22540
rect 21196 22482 21252 22494
rect 21196 22430 21198 22482
rect 21250 22430 21252 22482
rect 12796 22306 12852 22316
rect 13580 22372 13636 22382
rect 13580 22278 13636 22316
rect 13972 22372 14028 22382
rect 13972 22278 14028 22316
rect 19740 22370 19796 22382
rect 20748 22372 20804 22382
rect 19740 22318 19742 22370
rect 19794 22318 19796 22370
rect 19572 22260 19628 22270
rect 19572 22166 19628 22204
rect 19740 22260 19796 22318
rect 19740 22194 19796 22204
rect 20524 22370 20804 22372
rect 20524 22318 20750 22370
rect 20802 22318 20804 22370
rect 20524 22316 20804 22318
rect 13244 22148 13300 22158
rect 11676 21980 11956 22036
rect 12460 22146 13300 22148
rect 12460 22094 13246 22146
rect 13298 22094 13300 22146
rect 12460 22092 13300 22094
rect 11452 21868 11620 21924
rect 11340 21756 11508 21812
rect 10780 21588 10836 21598
rect 10780 21586 11060 21588
rect 10780 21534 10782 21586
rect 10834 21534 11060 21586
rect 10780 21532 11060 21534
rect 10780 21522 10836 21532
rect 9996 21420 10164 21476
rect 9660 21364 9716 21374
rect 9996 21364 10052 21420
rect 9660 21362 10052 21364
rect 9660 21310 9662 21362
rect 9714 21310 10052 21362
rect 9660 21308 10052 21310
rect 9660 21298 9716 21308
rect 9948 21196 10212 21206
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 9948 21130 10212 21140
rect 10332 21140 10388 21150
rect 9548 20862 9550 20914
rect 9602 20862 9604 20914
rect 9548 20850 9604 20862
rect 10332 20916 10388 21084
rect 9660 20804 9716 20814
rect 9884 20804 9940 20814
rect 9660 20711 9662 20748
rect 9714 20711 9716 20748
rect 9660 20188 9716 20711
rect 9548 20132 9716 20188
rect 9772 20802 9940 20804
rect 9772 20750 9886 20802
rect 9938 20750 9940 20802
rect 9772 20748 9940 20750
rect 9548 19684 9604 20132
rect 9660 20020 9716 20030
rect 9772 20020 9828 20748
rect 9884 20738 9940 20748
rect 10332 20188 10388 20860
rect 10444 20970 10500 20982
rect 10444 20918 10446 20970
rect 10498 20918 10500 20970
rect 10444 20580 10500 20918
rect 10892 20916 10948 20926
rect 11004 20916 11060 21532
rect 11340 21476 11396 21486
rect 11340 21382 11396 21420
rect 10948 20860 11060 20916
rect 11340 21140 11396 21150
rect 10556 20804 10612 20814
rect 10556 20710 10612 20748
rect 10892 20802 10948 20860
rect 10892 20750 10894 20802
rect 10946 20750 10948 20802
rect 10892 20738 10948 20750
rect 11340 20802 11396 21084
rect 11452 20970 11508 21756
rect 11452 20918 11454 20970
rect 11506 20918 11508 20970
rect 11452 20906 11508 20918
rect 11340 20750 11342 20802
rect 11394 20750 11396 20802
rect 11340 20738 11396 20750
rect 10444 20514 10500 20524
rect 11564 20244 11620 21868
rect 11676 21586 11732 21980
rect 11676 21534 11678 21586
rect 11730 21534 11732 21586
rect 11676 21522 11732 21534
rect 12012 21476 12068 21486
rect 12012 21474 12292 21476
rect 12012 21422 12014 21474
rect 12066 21422 12292 21474
rect 12012 21420 12292 21422
rect 12012 21410 12068 21420
rect 12124 20970 12180 20982
rect 12124 20918 12126 20970
rect 12178 20918 12180 20970
rect 11676 20804 11732 20814
rect 11676 20710 11732 20748
rect 12124 20804 12180 20918
rect 12124 20738 12180 20748
rect 12236 20916 12292 21420
rect 12236 20802 12292 20860
rect 12236 20750 12238 20802
rect 12290 20750 12292 20802
rect 12236 20738 12292 20750
rect 12236 20242 12292 20254
rect 12236 20190 12238 20242
rect 12290 20190 12292 20242
rect 12236 20188 12292 20190
rect 9716 19964 9828 20020
rect 9884 20132 9940 20142
rect 10332 20132 10500 20188
rect 11564 20178 11620 20188
rect 9884 20018 9940 20076
rect 9884 19966 9886 20018
rect 9938 19966 9940 20018
rect 9660 19926 9716 19964
rect 9884 19954 9940 19966
rect 10444 20018 10500 20132
rect 11900 20132 12292 20188
rect 10444 19966 10446 20018
rect 10498 19966 10500 20018
rect 10444 19954 10500 19966
rect 10668 20020 10724 20030
rect 11228 20020 11284 20030
rect 10668 19926 10724 19964
rect 10780 20018 11284 20020
rect 10780 19966 11230 20018
rect 11282 19966 11284 20018
rect 10780 19964 11284 19966
rect 10164 19796 10220 19806
rect 10780 19796 10836 19964
rect 11228 19954 11284 19964
rect 11452 20018 11508 20030
rect 11452 19966 11454 20018
rect 11506 19966 11508 20018
rect 10164 19794 10836 19796
rect 10164 19742 10166 19794
rect 10218 19742 10836 19794
rect 10164 19740 10836 19742
rect 10948 19796 11004 19806
rect 11452 19796 11508 19966
rect 11732 19908 11788 19918
rect 11732 19814 11788 19852
rect 10948 19794 11508 19796
rect 10948 19742 10950 19794
rect 11002 19742 11508 19794
rect 10948 19740 11508 19742
rect 10164 19730 10220 19740
rect 10948 19730 11004 19740
rect 9548 19628 9716 19684
rect 9492 19402 9548 19414
rect 9492 19350 9494 19402
rect 9546 19350 9548 19402
rect 9492 19236 9548 19350
rect 9492 19170 9548 19180
rect 9660 19348 9716 19628
rect 9948 19628 10212 19638
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 9948 19562 10212 19572
rect 11900 19460 11956 20132
rect 11116 19404 11956 19460
rect 12348 20020 12404 20030
rect 9660 19234 9716 19292
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 9660 19170 9716 19182
rect 9884 19346 9940 19358
rect 9884 19294 9886 19346
rect 9938 19294 9940 19346
rect 9884 19012 9940 19294
rect 10220 19236 10276 19246
rect 9324 18956 9940 19012
rect 9996 19190 10052 19202
rect 9996 19138 9998 19190
rect 10050 19138 10052 19190
rect 10220 19142 10276 19180
rect 10668 19234 10724 19246
rect 10668 19182 10670 19234
rect 10722 19182 10724 19234
rect 9996 18564 10052 19138
rect 9996 18498 10052 18508
rect 8428 18060 8932 18116
rect 8652 17892 8708 17902
rect 8092 17266 8148 17276
rect 8204 17666 8260 17678
rect 8204 17614 8206 17666
rect 8258 17614 8260 17666
rect 8204 17108 8260 17614
rect 8316 17668 8372 17678
rect 8316 17220 8372 17612
rect 8484 17668 8540 17678
rect 8484 17574 8540 17612
rect 8652 17666 8708 17836
rect 8652 17614 8654 17666
rect 8706 17614 8708 17666
rect 8652 17602 8708 17614
rect 8876 17666 8932 18060
rect 9948 18060 10212 18070
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 9948 17994 10212 18004
rect 10556 17780 10612 17790
rect 8876 17614 8878 17666
rect 8930 17614 8932 17666
rect 8540 17444 8596 17454
rect 8316 17154 8372 17164
rect 8502 17388 8540 17444
rect 8596 17388 8820 17444
rect 8502 17378 8596 17388
rect 7532 17052 8148 17108
rect 6412 16716 6804 16772
rect 6748 16660 6804 16716
rect 6748 16604 6916 16660
rect 6524 16212 6580 16222
rect 6524 16210 6804 16212
rect 6524 16158 6526 16210
rect 6578 16158 6804 16210
rect 6524 16156 6804 16158
rect 6524 16146 6580 16156
rect 5740 15362 5796 15372
rect 6300 16098 6356 16110
rect 6300 16046 6302 16098
rect 6354 16046 6356 16098
rect 6300 15876 6356 16046
rect 6636 16042 6692 16054
rect 6636 15990 6638 16042
rect 6690 15990 6692 16042
rect 6636 15988 6692 15990
rect 6636 15922 6692 15932
rect 6300 15370 6356 15820
rect 6748 15540 6804 16156
rect 6860 16098 6916 16604
rect 6860 16046 6862 16098
rect 6914 16046 6916 16098
rect 6860 16034 6916 16046
rect 7196 16098 7252 17052
rect 7868 16884 7980 16894
rect 7924 16882 7980 16884
rect 7924 16830 7926 16882
rect 7978 16830 7980 16882
rect 7924 16828 7980 16830
rect 7868 16818 7980 16828
rect 7196 16046 7198 16098
rect 7250 16046 7252 16098
rect 7196 16034 7252 16046
rect 7644 16660 7700 16670
rect 7644 16098 7700 16604
rect 7644 16046 7646 16098
rect 7698 16046 7700 16098
rect 7644 15988 7700 16046
rect 7644 15922 7700 15932
rect 7036 15708 7300 15718
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7036 15642 7300 15652
rect 6748 15484 7476 15540
rect 5628 15306 5684 15318
rect 6300 15318 6302 15370
rect 6354 15318 6356 15370
rect 6300 15306 6356 15318
rect 7254 15314 7310 15326
rect 7254 15262 7256 15314
rect 7308 15262 7310 15314
rect 7254 15204 7310 15262
rect 7420 15316 7476 15484
rect 7420 15222 7476 15260
rect 7532 15428 7588 15438
rect 7532 15316 7588 15372
rect 7756 15316 7812 15326
rect 7532 15314 7812 15316
rect 7532 15262 7534 15314
rect 7586 15262 7758 15314
rect 7810 15262 7812 15314
rect 7532 15260 7812 15262
rect 7532 15250 7588 15260
rect 7756 15250 7812 15260
rect 7254 15138 7310 15148
rect 6412 15092 6468 15102
rect 5796 14532 5852 14542
rect 4956 14476 5124 14532
rect 4900 14308 4956 14318
rect 4900 14214 4956 14252
rect 4844 13860 4900 13870
rect 4844 13746 4900 13804
rect 4844 13694 4846 13746
rect 4898 13694 4900 13746
rect 4844 13682 4900 13694
rect 4620 13570 4676 13580
rect 4900 13524 4956 13534
rect 4900 13074 4956 13468
rect 4900 13022 4902 13074
rect 4954 13022 4956 13074
rect 4900 13010 4956 13022
rect 5068 12964 5124 14476
rect 5796 14438 5852 14476
rect 6076 13412 6132 13422
rect 5068 12898 5124 12908
rect 5628 13130 5684 13142
rect 5628 13078 5630 13130
rect 5682 13078 5684 13130
rect 5180 12404 5236 12414
rect 4284 11564 4564 11620
rect 4732 12292 4788 12302
rect 3948 11508 4004 11518
rect 3948 11361 4004 11452
rect 3948 11309 3950 11361
rect 4002 11309 4004 11361
rect 3948 11297 4004 11309
rect 4284 11357 4340 11564
rect 4284 11305 4286 11357
rect 4338 11305 4340 11357
rect 4284 10836 4340 11305
rect 4060 10780 4340 10836
rect 4620 11338 4676 11350
rect 4620 11286 4622 11338
rect 4674 11286 4676 11338
rect 4620 11284 4676 11286
rect 4060 10668 4116 10780
rect 3276 10558 3278 10610
rect 3330 10558 3332 10610
rect 3556 10639 4116 10668
rect 3556 10587 3558 10639
rect 3610 10612 4116 10639
rect 3610 10587 3612 10612
rect 3556 10575 3612 10587
rect 4060 10610 4116 10612
rect 3276 10546 3332 10558
rect 4060 10558 4062 10610
rect 4114 10558 4116 10610
rect 4060 10546 4116 10558
rect 4284 10612 4340 10622
rect 4620 10612 4676 11228
rect 4284 10610 4676 10612
rect 4284 10558 4286 10610
rect 4338 10558 4676 10610
rect 4732 10666 4788 12236
rect 5068 12292 5124 12302
rect 4956 12180 5012 12190
rect 4956 11844 5012 12124
rect 5068 12178 5124 12236
rect 5068 12126 5070 12178
rect 5122 12126 5124 12178
rect 5068 12114 5124 12126
rect 5180 12010 5236 12348
rect 5404 12180 5460 12190
rect 5628 12180 5684 13078
rect 5740 12964 5796 12974
rect 5740 12870 5796 12908
rect 5964 12964 6020 12974
rect 5964 12740 6020 12908
rect 5964 12674 6020 12684
rect 5404 12086 5460 12124
rect 5516 12178 5684 12180
rect 5516 12126 5630 12178
rect 5682 12126 5684 12178
rect 5516 12124 5684 12126
rect 5180 11958 5182 12010
rect 5234 11958 5236 12010
rect 5180 11946 5236 11958
rect 4930 11788 5012 11844
rect 4930 11361 4986 11788
rect 4930 11309 4932 11361
rect 4984 11309 4986 11361
rect 4930 11297 4986 11309
rect 5068 11396 5124 11406
rect 4732 10614 4734 10666
rect 4786 10614 4788 10666
rect 5068 11282 5124 11340
rect 5068 11230 5070 11282
rect 5122 11230 5124 11282
rect 5068 10666 5124 11230
rect 5516 11060 5572 12124
rect 5628 12114 5684 12124
rect 5908 11956 5964 11966
rect 6076 11956 6132 13356
rect 5908 11954 6132 11956
rect 5908 11902 5910 11954
rect 5962 11902 6132 11954
rect 5908 11900 6132 11902
rect 5908 11890 5964 11900
rect 6076 11844 6132 11900
rect 6076 11620 6132 11788
rect 5964 11564 6132 11620
rect 6188 12292 6244 12302
rect 5796 11508 5852 11518
rect 5796 11450 5852 11452
rect 5628 11396 5684 11406
rect 5796 11398 5798 11450
rect 5850 11398 5852 11450
rect 5796 11386 5852 11398
rect 5964 11394 6020 11564
rect 5628 11302 5684 11340
rect 5964 11342 5966 11394
rect 6018 11342 6020 11394
rect 5964 11330 6020 11342
rect 6076 11396 6132 11406
rect 6188 11396 6244 12236
rect 6412 12180 6468 15036
rect 6860 15092 6916 15102
rect 6860 14998 6916 15036
rect 7420 15092 7476 15102
rect 7868 15092 7924 16818
rect 7980 16100 8036 16110
rect 7980 16006 8036 16044
rect 7980 15316 8036 15326
rect 7980 15222 8036 15260
rect 6524 14532 6580 14542
rect 6524 13748 6580 14476
rect 7036 14140 7300 14150
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7036 14074 7300 14084
rect 6972 13860 7028 13870
rect 6524 13524 6580 13692
rect 6524 13458 6580 13468
rect 6860 13746 6916 13758
rect 6860 13694 6862 13746
rect 6914 13694 6916 13746
rect 6748 13300 6804 13310
rect 6748 12964 6804 13244
rect 6860 13188 6916 13694
rect 6860 13122 6916 13132
rect 6972 13524 7028 13804
rect 7252 13802 7364 13860
rect 7252 13750 7254 13802
rect 7306 13750 7364 13802
rect 7252 13738 7364 13750
rect 7196 13634 7252 13646
rect 7196 13582 7198 13634
rect 7250 13582 7252 13634
rect 7196 13524 7252 13582
rect 6972 13468 7252 13524
rect 6860 12964 6916 12974
rect 6748 12962 6916 12964
rect 6748 12910 6862 12962
rect 6914 12910 6916 12962
rect 6748 12908 6916 12910
rect 6860 12898 6916 12908
rect 6524 12740 6580 12750
rect 6972 12740 7028 13468
rect 7084 13076 7140 13086
rect 7084 12962 7140 13020
rect 7308 12974 7364 13738
rect 7420 13746 7476 15036
rect 7756 15036 7924 15092
rect 7420 13694 7422 13746
rect 7474 13694 7476 13746
rect 7420 13682 7476 13694
rect 7532 13860 7588 13870
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 12898 7140 12910
rect 7252 12964 7364 12974
rect 7308 12908 7364 12964
rect 7420 13188 7476 13198
rect 7420 12962 7476 13132
rect 7420 12910 7422 12962
rect 7474 12910 7476 12962
rect 7252 12870 7308 12908
rect 7420 12898 7476 12910
rect 7532 12962 7588 13804
rect 7756 13748 7812 15036
rect 7756 13682 7812 13692
rect 7868 14532 7924 14542
rect 7868 13746 7924 14476
rect 8092 14308 8148 17052
rect 8204 17042 8260 17052
rect 8316 16996 8372 17006
rect 8204 16884 8260 16894
rect 8204 16790 8260 16828
rect 8316 16882 8372 16940
rect 8316 16830 8318 16882
rect 8370 16830 8372 16882
rect 8502 16920 8558 17378
rect 8502 16868 8504 16920
rect 8556 16868 8558 16920
rect 8502 16856 8558 16868
rect 8652 17220 8708 17230
rect 8316 16818 8372 16830
rect 8428 16660 8484 16670
rect 8428 15540 8484 16604
rect 8652 16322 8708 17164
rect 8764 16884 8820 17388
rect 8876 16996 8932 17614
rect 9212 17668 9268 17678
rect 9212 17444 9268 17612
rect 9212 17442 9380 17444
rect 9212 17390 9214 17442
rect 9266 17390 9380 17442
rect 9212 17388 9380 17390
rect 9212 17378 9268 17388
rect 8876 16930 8932 16940
rect 8988 17108 9044 17118
rect 8764 16818 8820 16828
rect 8652 16270 8654 16322
rect 8706 16270 8708 16322
rect 8652 16258 8708 16270
rect 8876 16658 8932 16670
rect 8876 16606 8878 16658
rect 8930 16606 8932 16658
rect 8708 15540 8764 15550
rect 8428 15538 8764 15540
rect 8428 15486 8710 15538
rect 8762 15486 8764 15538
rect 8428 15484 8764 15486
rect 8260 15090 8316 15102
rect 8260 15038 8262 15090
rect 8314 15038 8316 15090
rect 8260 14532 8316 15038
rect 8260 14466 8316 14476
rect 8428 14308 8484 15484
rect 8708 15474 8764 15484
rect 8876 15540 8932 16606
rect 8988 16098 9044 17052
rect 8988 16046 8990 16098
rect 9042 16046 9044 16098
rect 8988 16034 9044 16046
rect 9324 16098 9380 17388
rect 9884 16996 9940 17006
rect 9884 16938 9940 16940
rect 9548 16884 9604 16894
rect 9884 16886 9886 16938
rect 9938 16886 9940 16938
rect 9884 16874 9940 16886
rect 10220 16996 10276 17006
rect 10220 16882 10276 16940
rect 9548 16790 9604 16828
rect 10220 16830 10222 16882
rect 10274 16830 10276 16882
rect 10220 16818 10276 16830
rect 10556 16882 10612 17724
rect 10668 17444 10724 19182
rect 10836 19236 10892 19246
rect 10836 19142 10892 19180
rect 11116 19234 11172 19404
rect 11116 19182 11118 19234
rect 11170 19182 11172 19234
rect 11116 19170 11172 19182
rect 11004 19124 11060 19134
rect 11004 18450 11060 19068
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 18386 11060 18398
rect 11116 18564 11172 18574
rect 11116 18282 11172 18508
rect 11228 18452 11284 19404
rect 12068 19348 12124 19358
rect 12068 19290 12124 19292
rect 11396 19236 11452 19246
rect 11396 19142 11452 19180
rect 11900 19236 11956 19246
rect 12068 19238 12070 19290
rect 12122 19238 12124 19290
rect 12068 19226 12124 19238
rect 12348 19234 12404 19964
rect 11900 19142 11956 19180
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12236 19122 12292 19134
rect 12236 19070 12238 19122
rect 12290 19070 12292 19122
rect 11340 18452 11396 18462
rect 12012 18452 12068 18462
rect 11228 18450 11620 18452
rect 11228 18398 11342 18450
rect 11394 18398 11620 18450
rect 11228 18396 11620 18398
rect 11340 18386 11396 18396
rect 11116 18230 11118 18282
rect 11170 18230 11172 18282
rect 11116 18218 11172 18230
rect 11116 17892 11172 17902
rect 11116 17666 11172 17836
rect 11116 17614 11118 17666
rect 11170 17614 11172 17666
rect 11116 17602 11172 17614
rect 11564 17890 11620 18396
rect 12012 18358 12068 18396
rect 11564 17838 11566 17890
rect 11618 17838 11620 17890
rect 11564 17668 11620 17838
rect 11844 18226 11900 18238
rect 11844 18174 11846 18226
rect 11898 18174 11900 18226
rect 11844 17892 11900 18174
rect 11844 17826 11900 17836
rect 12124 18228 12180 18238
rect 11900 17668 11956 17678
rect 11564 17602 11620 17612
rect 11788 17666 11956 17668
rect 11788 17614 11902 17666
rect 11954 17614 11956 17666
rect 11788 17612 11956 17614
rect 10780 17444 10836 17454
rect 10668 17442 10836 17444
rect 10668 17390 10782 17442
rect 10834 17390 10836 17442
rect 10668 17388 10836 17390
rect 10556 16830 10558 16882
rect 10610 16830 10612 16882
rect 10556 16818 10612 16830
rect 9324 16046 9326 16098
rect 9378 16046 9380 16098
rect 9324 16034 9380 16046
rect 9772 16770 9828 16782
rect 9772 16718 9774 16770
rect 9826 16718 9828 16770
rect 9660 15876 9716 15886
rect 9660 15782 9716 15820
rect 8876 15474 8932 15484
rect 8876 15314 8932 15326
rect 8876 15262 8878 15314
rect 8930 15262 8932 15314
rect 8876 15204 8932 15262
rect 9772 15316 9828 16718
rect 9948 16492 10212 16502
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 9948 16426 10212 16436
rect 10556 15876 10612 15886
rect 10220 15540 10276 15550
rect 9660 15204 9716 15214
rect 8876 15202 9716 15204
rect 8876 15150 9662 15202
rect 9714 15150 9716 15202
rect 8876 15148 9716 15150
rect 8764 14502 8820 14514
rect 8764 14450 8766 14502
rect 8818 14450 8820 14502
rect 8764 14420 8820 14450
rect 8764 14354 8820 14364
rect 8092 14252 8182 14308
rect 7868 13694 7870 13746
rect 7922 13694 7924 13746
rect 7532 12910 7534 12962
rect 7586 12910 7588 12962
rect 7532 12852 7588 12910
rect 7532 12786 7588 12796
rect 7644 13524 7700 13534
rect 7644 13076 7700 13468
rect 7868 13076 7924 13694
rect 7980 13860 8036 13870
rect 7980 13746 8036 13804
rect 7980 13694 7982 13746
rect 8034 13694 8036 13746
rect 7980 13682 8036 13694
rect 8126 13784 8182 14252
rect 8316 14252 8484 14308
rect 8316 13860 8372 14252
rect 8316 13794 8372 13804
rect 8126 13732 8128 13784
rect 8180 13732 8182 13784
rect 8126 13300 8182 13732
rect 8540 13524 8596 13534
rect 8540 13430 8596 13468
rect 8126 13234 8182 13244
rect 7868 13020 8148 13076
rect 6524 12738 6838 12740
rect 6524 12686 6526 12738
rect 6578 12686 6838 12738
rect 6524 12684 6838 12686
rect 6972 12684 7476 12740
rect 6524 12674 6580 12684
rect 6636 12292 6692 12302
rect 6524 12180 6580 12190
rect 6412 12178 6580 12180
rect 6412 12126 6526 12178
rect 6578 12126 6580 12178
rect 6412 12124 6580 12126
rect 6412 11508 6468 12124
rect 6524 12114 6580 12124
rect 6636 12178 6692 12236
rect 6636 12126 6638 12178
rect 6690 12126 6692 12178
rect 6636 12114 6692 12126
rect 6782 12216 6838 12684
rect 7036 12572 7300 12582
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7036 12506 7300 12516
rect 7420 12292 7476 12684
rect 7644 12628 7700 13020
rect 7812 12852 7868 12862
rect 7812 12850 8036 12852
rect 7812 12798 7814 12850
rect 7866 12798 8036 12850
rect 7812 12796 8036 12798
rect 7812 12786 7868 12796
rect 7644 12572 7868 12628
rect 7644 12292 7700 12302
rect 7420 12290 7700 12292
rect 7420 12238 7646 12290
rect 7698 12238 7700 12290
rect 7420 12236 7700 12238
rect 7644 12226 7700 12236
rect 7812 12234 7868 12572
rect 6782 12180 6784 12216
rect 6836 12180 6838 12216
rect 6782 12086 6838 12124
rect 7196 12180 7252 12190
rect 7812 12182 7814 12234
rect 7866 12182 7868 12234
rect 7812 12170 7868 12182
rect 7196 12066 7252 12124
rect 7196 12014 7198 12066
rect 7250 12014 7252 12066
rect 7196 12002 7252 12014
rect 7420 12068 7476 12078
rect 6412 11442 6468 11452
rect 6860 11844 6916 11854
rect 6076 11394 6244 11396
rect 6076 11342 6078 11394
rect 6130 11342 6244 11394
rect 6076 11340 6244 11342
rect 6076 11284 6132 11340
rect 6356 11284 6412 11294
rect 6076 11218 6132 11228
rect 6300 11282 6412 11284
rect 6300 11230 6358 11282
rect 6410 11230 6412 11282
rect 6300 11218 6412 11230
rect 5516 11004 5952 11060
rect 4732 10602 4788 10614
rect 4844 10638 4900 10650
rect 4284 10556 4676 10558
rect 4844 10586 4846 10638
rect 4898 10586 4900 10638
rect 5068 10614 5070 10666
rect 5122 10614 5124 10666
rect 5068 10602 5124 10614
rect 5292 10638 5348 10650
rect 5292 10612 5294 10638
rect 5346 10612 5348 10638
rect 4284 10546 4340 10556
rect 3612 10498 3668 10510
rect 4844 10500 4900 10586
rect 5896 10648 5952 11004
rect 5896 10596 5898 10648
rect 5950 10596 5952 10648
rect 5896 10584 5952 10596
rect 5292 10546 5348 10556
rect 3612 10446 3614 10498
rect 3666 10446 3668 10498
rect 3612 10388 3668 10446
rect 4396 10444 4900 10500
rect 4396 10442 4452 10444
rect 4396 10390 4398 10442
rect 4450 10390 4452 10442
rect 4396 10378 4452 10390
rect 5572 10388 5628 10398
rect 5516 10386 5628 10388
rect 3612 10322 3668 10332
rect 5516 10334 5574 10386
rect 5626 10334 5628 10386
rect 5516 10322 5628 10334
rect 4124 10220 4388 10230
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4124 10154 4388 10164
rect 4956 9042 5012 9054
rect 4956 8990 4958 9042
rect 5010 8990 5012 9042
rect 4124 8652 4388 8662
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4124 8586 4388 8596
rect 4956 8428 5012 8990
rect 4956 8372 5236 8428
rect 5180 7474 5236 8316
rect 5516 8258 5572 10322
rect 6300 9268 6356 11218
rect 6860 10668 6916 11788
rect 7420 11394 7476 12012
rect 7420 11342 7422 11394
rect 7474 11342 7476 11394
rect 7420 11060 7476 11342
rect 7036 11004 7300 11014
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7420 10994 7476 11004
rect 7532 11562 7588 11574
rect 7532 11510 7534 11562
rect 7586 11510 7588 11562
rect 7036 10938 7300 10948
rect 7308 10836 7364 10846
rect 7532 10836 7588 11510
rect 6412 10612 6468 10622
rect 6412 10442 6468 10556
rect 6412 10390 6414 10442
rect 6466 10390 6468 10442
rect 6412 10378 6468 10390
rect 6692 10610 6748 10622
rect 6860 10612 7252 10668
rect 6692 10558 6694 10610
rect 6746 10558 6748 10610
rect 6692 10052 6748 10558
rect 7196 10610 7252 10612
rect 7196 10558 7198 10610
rect 7250 10558 7252 10610
rect 7196 10546 7252 10558
rect 6692 9958 6748 9996
rect 6972 10500 7028 10510
rect 6972 9826 7028 10444
rect 7308 10388 7364 10780
rect 6972 9774 6974 9826
rect 7026 9774 7028 9826
rect 6972 9762 7028 9774
rect 7196 10332 7364 10388
rect 7420 10780 7588 10836
rect 7756 11394 7812 11406
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 7756 10836 7812 11342
rect 7980 11284 8036 12796
rect 8092 12068 8148 13020
rect 8652 12964 8708 12974
rect 8876 12964 8932 15148
rect 9660 15138 9716 15148
rect 9772 14980 9828 15260
rect 10052 15314 10108 15326
rect 10052 15262 10054 15314
rect 10106 15262 10108 15314
rect 10052 15204 10108 15262
rect 10052 15138 10108 15148
rect 10220 15314 10276 15484
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 10220 15092 10276 15262
rect 10332 15316 10388 15326
rect 10332 15222 10388 15260
rect 10556 15314 10612 15820
rect 10556 15262 10558 15314
rect 10610 15262 10612 15314
rect 10556 15250 10612 15262
rect 10780 15316 10836 17388
rect 11788 16882 11844 17612
rect 11900 17602 11956 17612
rect 12124 16884 12180 18172
rect 12236 17834 12292 19070
rect 12348 18564 12404 19182
rect 12348 18498 12404 18508
rect 12460 18452 12516 22092
rect 13244 22082 13300 22092
rect 20076 22146 20132 22158
rect 20076 22094 20078 22146
rect 20130 22094 20132 22146
rect 12860 21980 13124 21990
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 12860 21914 13124 21924
rect 18684 21980 18948 21990
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18684 21914 18948 21924
rect 20076 21924 20132 22094
rect 20076 21858 20132 21868
rect 17836 21700 17892 21710
rect 14700 21586 14756 21598
rect 14924 21588 14980 21598
rect 15260 21588 15316 21598
rect 14700 21534 14702 21586
rect 14754 21534 14756 21586
rect 13916 21476 13972 21486
rect 13916 21382 13972 21420
rect 14700 20804 14756 21534
rect 14812 21586 14980 21588
rect 14812 21534 14926 21586
rect 14978 21534 14980 21586
rect 14812 21532 14980 21534
rect 14812 21140 14868 21532
rect 14924 21522 14980 21532
rect 15036 21586 15316 21588
rect 15036 21534 15262 21586
rect 15314 21534 15316 21586
rect 15036 21532 15316 21534
rect 15036 21252 15092 21532
rect 15260 21522 15316 21532
rect 15596 21586 15652 21598
rect 17276 21588 17332 21598
rect 15596 21534 15598 21586
rect 15650 21534 15652 21586
rect 14812 21074 14868 21084
rect 14924 21196 15092 21252
rect 15260 21418 15316 21430
rect 15260 21366 15262 21418
rect 15314 21366 15316 21418
rect 14924 20970 14980 21196
rect 12912 20764 12968 20776
rect 12912 20712 12914 20764
rect 12966 20712 12968 20764
rect 12912 20580 12968 20712
rect 12684 20524 12968 20580
rect 14136 20764 14192 20776
rect 14136 20712 14138 20764
rect 14190 20712 14192 20764
rect 14700 20738 14756 20748
rect 14812 20916 14868 20926
rect 14924 20918 14926 20970
rect 14978 20918 14980 20970
rect 14924 20906 14980 20918
rect 14812 20802 14868 20860
rect 14812 20750 14814 20802
rect 14866 20750 14868 20802
rect 14812 20738 14868 20750
rect 15148 20804 15204 20814
rect 12684 20242 12740 20524
rect 14136 20468 14192 20712
rect 15148 20710 15204 20748
rect 15260 20580 15316 21366
rect 15260 20524 15350 20580
rect 12860 20412 13124 20422
rect 14136 20412 14196 20468
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 12860 20346 13124 20356
rect 12684 20190 12686 20242
rect 12738 20190 12740 20242
rect 12684 20178 12740 20190
rect 13804 20132 13860 20142
rect 13580 19348 13636 19358
rect 13580 19254 13636 19292
rect 13692 19236 13748 19246
rect 12628 19124 12684 19134
rect 12628 19122 13412 19124
rect 12628 19070 12630 19122
rect 12682 19070 13412 19122
rect 12628 19068 13412 19070
rect 12628 19058 12684 19068
rect 12860 18844 13124 18854
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 12860 18778 13124 18788
rect 12460 18386 12516 18396
rect 12908 18452 12964 18462
rect 12908 18358 12964 18396
rect 13356 18450 13412 19068
rect 13356 18398 13358 18450
rect 13410 18398 13412 18450
rect 13356 18386 13412 18398
rect 13692 18450 13748 19180
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13692 18386 13748 18398
rect 12572 18228 12628 18238
rect 12572 18134 12628 18172
rect 12236 17782 12238 17834
rect 12290 17782 12292 17834
rect 13692 17892 13748 17902
rect 13804 17892 13860 20076
rect 14140 20132 14196 20412
rect 14140 20066 14196 20076
rect 15148 20132 15204 20142
rect 15036 20020 15092 20030
rect 14364 20018 15092 20020
rect 14364 19966 15038 20018
rect 15090 19966 15092 20018
rect 14364 19964 15092 19966
rect 14364 18228 14420 19964
rect 15036 19954 15092 19964
rect 15148 20018 15204 20076
rect 15148 19966 15150 20018
rect 15202 19966 15204 20018
rect 15294 20056 15350 20524
rect 15294 20004 15296 20056
rect 15348 20004 15350 20056
rect 15294 19992 15350 20004
rect 15148 19954 15204 19966
rect 15596 19908 15652 21534
rect 17052 21532 17276 21588
rect 15932 21364 15988 21374
rect 15932 21362 16212 21364
rect 15932 21310 15934 21362
rect 15986 21310 16212 21362
rect 15932 21308 16212 21310
rect 15932 21298 15988 21308
rect 15772 21196 16036 21206
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 15772 21130 16036 21140
rect 15932 20916 15988 20926
rect 16156 20916 16212 21308
rect 15932 20914 16212 20916
rect 15932 20862 15934 20914
rect 15986 20862 16212 20914
rect 15932 20860 16212 20862
rect 15932 20850 15988 20860
rect 17052 20804 17108 21532
rect 17276 21494 17332 21532
rect 17836 20916 17892 21644
rect 17836 20822 17892 20860
rect 18060 21474 18116 21486
rect 18060 21422 18062 21474
rect 18114 21422 18116 21474
rect 15708 19908 15764 19918
rect 15596 19906 15764 19908
rect 15596 19854 15710 19906
rect 15762 19854 15764 19906
rect 15596 19852 15764 19854
rect 15708 19842 15764 19852
rect 15772 19628 16036 19638
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 15772 19562 16036 19572
rect 17052 19348 17108 20748
rect 18060 20242 18116 21422
rect 19964 21476 20020 21486
rect 19964 21474 20132 21476
rect 19964 21422 19966 21474
rect 20018 21422 20132 21474
rect 19964 21420 20132 21422
rect 19964 21410 20020 21420
rect 19292 20916 19348 20926
rect 19516 20916 19908 20972
rect 19292 20914 19572 20916
rect 19292 20862 19294 20914
rect 19346 20862 19572 20914
rect 19292 20860 19572 20862
rect 19292 20850 19348 20860
rect 18956 20804 19012 20814
rect 19628 20802 19684 20814
rect 18956 20710 19012 20748
rect 19180 20758 19236 20770
rect 19180 20706 19182 20758
rect 19234 20706 19236 20758
rect 18684 20412 18948 20422
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18684 20346 18948 20356
rect 19180 20356 19236 20706
rect 19180 20290 19236 20300
rect 19628 20750 19630 20802
rect 19682 20750 19684 20802
rect 18060 20190 18062 20242
rect 18114 20190 18116 20242
rect 18060 20178 18116 20190
rect 18396 20244 18452 20254
rect 18396 20018 18452 20188
rect 19404 20020 19460 20030
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19954 18452 19966
rect 19292 19964 19404 20020
rect 19628 20020 19684 20750
rect 19852 20804 19908 20916
rect 20076 20804 20132 21420
rect 19852 20748 19964 20804
rect 19908 20746 19964 20748
rect 19908 20694 19910 20746
rect 19962 20694 19964 20746
rect 20076 20738 20132 20748
rect 20300 21028 20356 21038
rect 20300 20802 20356 20972
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 20300 20738 20356 20750
rect 20412 20804 20468 20814
rect 19908 20682 19964 20694
rect 19740 20634 19796 20646
rect 19740 20582 19742 20634
rect 19794 20582 19796 20634
rect 19740 20244 19796 20582
rect 20412 20580 20468 20748
rect 19740 20178 19796 20188
rect 20356 20524 20468 20580
rect 20356 20074 20412 20524
rect 19740 20020 19796 20030
rect 20188 20020 20244 20030
rect 19628 20018 20020 20020
rect 19628 19966 19742 20018
rect 19794 19966 20020 20018
rect 19628 19964 20020 19966
rect 19292 19918 19348 19964
rect 19404 19926 19460 19964
rect 19740 19954 19796 19964
rect 18788 19908 18844 19918
rect 19236 19908 19348 19918
rect 18788 19906 19348 19908
rect 18788 19854 18790 19906
rect 18842 19854 19238 19906
rect 19290 19854 19348 19906
rect 18788 19852 19348 19854
rect 18788 19842 18844 19852
rect 19236 19842 19348 19852
rect 16828 19292 17332 19348
rect 15484 19236 15540 19246
rect 15484 19142 15540 19180
rect 16268 19236 16324 19246
rect 16828 19236 16884 19292
rect 16268 19234 16884 19236
rect 16268 19182 16270 19234
rect 16322 19182 16830 19234
rect 16882 19182 16884 19234
rect 16268 19180 16884 19182
rect 16268 19170 16324 19180
rect 16828 19170 16884 19180
rect 15148 18452 15204 18462
rect 15148 18450 15428 18452
rect 15148 18398 15150 18450
rect 15202 18398 15428 18450
rect 15148 18396 15428 18398
rect 15148 18386 15204 18396
rect 14364 18172 14644 18228
rect 13692 17890 13860 17892
rect 13692 17838 13694 17890
rect 13746 17838 13860 17890
rect 13692 17836 13860 17838
rect 13692 17826 13748 17836
rect 12236 17770 12292 17782
rect 14588 17780 14644 18172
rect 14588 17686 14644 17724
rect 15148 17780 15204 17790
rect 12236 17668 12292 17678
rect 12236 17574 12292 17612
rect 12460 17666 12516 17678
rect 13356 17668 13412 17678
rect 12460 17614 12462 17666
rect 12514 17614 12516 17666
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16212 11844 16830
rect 11788 16146 11844 16156
rect 12012 16828 12124 16884
rect 10780 15250 10836 15260
rect 11228 16098 11284 16110
rect 11228 16046 11230 16098
rect 11282 16046 11284 16098
rect 11228 15316 11284 16046
rect 11452 16100 11508 16110
rect 11452 16006 11508 16044
rect 12012 16098 12068 16828
rect 12124 16818 12180 16828
rect 12348 16882 12404 16894
rect 12348 16830 12350 16882
rect 12402 16830 12404 16882
rect 12348 16436 12404 16830
rect 12012 16046 12014 16098
rect 12066 16046 12068 16098
rect 12012 16034 12068 16046
rect 12124 16380 12404 16436
rect 11732 15988 11788 15998
rect 11732 15894 11788 15932
rect 11228 15250 11284 15260
rect 12012 15316 12068 15326
rect 12124 15316 12180 16380
rect 12460 16324 12516 17614
rect 13244 17666 13412 17668
rect 13244 17614 13358 17666
rect 13410 17614 13412 17666
rect 13244 17612 13412 17614
rect 12860 17276 13124 17286
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 12860 17210 13124 17220
rect 12572 17052 12628 17062
rect 12572 17050 13076 17052
rect 12572 16998 12574 17050
rect 12626 16998 13076 17050
rect 12572 16996 13076 16998
rect 12572 16986 12628 16996
rect 12908 16884 12964 16894
rect 13020 16884 13076 16996
rect 13132 16884 13188 16894
rect 13244 16884 13300 17612
rect 13356 17602 13412 17612
rect 14476 16996 14980 17052
rect 13020 16882 13300 16884
rect 13020 16830 13134 16882
rect 13186 16830 13300 16882
rect 13020 16828 13300 16830
rect 13412 16884 13468 16894
rect 12908 16790 12964 16828
rect 13132 16818 13188 16828
rect 13412 16790 13468 16828
rect 14252 16884 14308 16894
rect 12348 16268 12516 16324
rect 12236 16100 12292 16110
rect 12236 16006 12292 16044
rect 12348 15540 12404 16268
rect 12516 16100 12572 16110
rect 12516 16006 12572 16044
rect 14252 15876 14308 16828
rect 14476 16334 14532 16996
rect 14588 16917 14644 16929
rect 14588 16865 14590 16917
rect 14642 16865 14644 16917
rect 14588 16548 14644 16865
rect 14700 16910 14756 16922
rect 14700 16884 14702 16910
rect 14754 16884 14756 16910
rect 14924 16910 14980 16996
rect 14924 16858 14926 16910
rect 14978 16858 14980 16910
rect 15148 16938 15204 17724
rect 15372 17006 15428 18396
rect 15484 18228 15540 18238
rect 15484 18226 16548 18228
rect 15484 18174 15486 18226
rect 15538 18174 16548 18226
rect 15484 18172 16548 18174
rect 15484 18162 15540 18172
rect 15772 18060 16036 18070
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 15772 17994 16036 18004
rect 16492 17778 16548 18172
rect 16492 17726 16494 17778
rect 16546 17726 16548 17778
rect 16492 17714 16548 17726
rect 17276 17668 17332 19292
rect 17612 19236 17668 19246
rect 17612 19234 17892 19236
rect 17612 19182 17614 19234
rect 17666 19182 17892 19234
rect 17612 19180 17892 19182
rect 17612 19170 17668 19180
rect 17836 18674 17892 19180
rect 18684 18844 18948 18854
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18684 18778 18948 18788
rect 17836 18622 17838 18674
rect 17890 18622 17892 18674
rect 17836 18610 17892 18622
rect 18172 18452 18228 18462
rect 18172 18358 18228 18396
rect 17388 17668 17444 17678
rect 17276 17666 17444 17668
rect 17276 17614 17278 17666
rect 17330 17614 17390 17666
rect 17442 17614 17444 17666
rect 17276 17612 17444 17614
rect 17276 17602 17332 17612
rect 15372 16994 15484 17006
rect 15372 16942 15430 16994
rect 15482 16942 15484 16994
rect 15372 16940 15484 16942
rect 15148 16886 15150 16938
rect 15202 16886 15204 16938
rect 15428 16930 15484 16940
rect 15148 16874 15204 16886
rect 14924 16846 14980 16858
rect 14700 16818 14756 16828
rect 14588 16492 14868 16548
rect 14476 16324 14588 16334
rect 14476 16322 14756 16324
rect 14476 16270 14534 16322
rect 14586 16270 14756 16322
rect 14476 16268 14756 16270
rect 14532 16258 14588 16268
rect 14364 16100 14420 16110
rect 14420 16044 14644 16100
rect 14364 16006 14420 16044
rect 14252 15820 14532 15876
rect 12860 15708 13124 15718
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 12860 15642 13124 15652
rect 12348 15446 12404 15484
rect 13580 15540 13636 15550
rect 12012 15314 12180 15316
rect 12012 15262 12014 15314
rect 12066 15262 12180 15314
rect 12012 15260 12180 15262
rect 10892 15204 10948 15214
rect 10892 15110 10948 15148
rect 12012 15204 12068 15260
rect 10220 15036 10388 15092
rect 9548 14924 9828 14980
rect 9948 14924 10212 14934
rect 9436 14642 9492 14654
rect 9436 14590 9438 14642
rect 9490 14590 9492 14642
rect 9100 14530 9156 14542
rect 9100 14478 9102 14530
rect 9154 14478 9156 14530
rect 9100 14308 9156 14478
rect 9100 14242 9156 14252
rect 9212 13748 9268 13758
rect 9044 13076 9100 13086
rect 9212 13076 9268 13692
rect 9044 13074 9268 13076
rect 9044 13022 9046 13074
rect 9098 13022 9268 13074
rect 9044 13020 9268 13022
rect 9044 13010 9100 13020
rect 8652 12962 8932 12964
rect 8652 12910 8654 12962
rect 8706 12910 8932 12962
rect 8652 12908 8932 12910
rect 9212 12962 9268 13020
rect 9212 12910 9214 12962
rect 9266 12910 9268 12962
rect 8652 12898 8708 12908
rect 9212 12898 9268 12910
rect 8316 12740 8372 12750
rect 8204 12738 8372 12740
rect 8204 12686 8318 12738
rect 8370 12686 8372 12738
rect 8204 12684 8372 12686
rect 8204 12292 8260 12684
rect 8316 12674 8372 12684
rect 8204 12226 8260 12236
rect 8316 12180 8372 12190
rect 8316 12086 8372 12124
rect 8558 12180 8614 12190
rect 8558 12086 8614 12124
rect 9436 12178 9492 14590
rect 9548 14491 9604 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 9948 14858 10212 14868
rect 10332 14756 10388 15036
rect 9548 14439 9550 14491
rect 9602 14439 9604 14491
rect 9772 14700 10388 14756
rect 9772 14530 9828 14700
rect 9772 14478 9774 14530
rect 9826 14478 9828 14530
rect 9772 14466 9828 14478
rect 10108 14530 10164 14542
rect 10108 14478 10110 14530
rect 10162 14478 10164 14530
rect 9548 14427 9604 14439
rect 10108 13524 10164 14478
rect 11116 14420 11172 14430
rect 10948 13636 11004 13646
rect 10948 13542 11004 13580
rect 10108 13458 10164 13468
rect 9948 13356 10212 13366
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 9948 13290 10212 13300
rect 9996 12962 10052 12974
rect 9996 12910 9998 12962
rect 10050 12910 10052 12962
rect 9996 12404 10052 12910
rect 9996 12338 10052 12348
rect 10668 12404 10724 12414
rect 10500 12292 10556 12302
rect 10500 12234 10556 12236
rect 9436 12126 9438 12178
rect 9490 12126 9492 12178
rect 8092 12002 8148 12012
rect 9436 11620 9492 12126
rect 9660 12180 9716 12190
rect 9660 12086 9716 12124
rect 10332 12178 10388 12190
rect 10332 12126 10334 12178
rect 10386 12126 10388 12178
rect 10500 12182 10502 12234
rect 10554 12182 10556 12234
rect 10500 12170 10556 12182
rect 10332 12068 10388 12126
rect 10332 12002 10388 12012
rect 9940 11956 9996 11966
rect 9772 11954 9996 11956
rect 9772 11902 9942 11954
rect 9994 11902 9996 11954
rect 9772 11900 9996 11902
rect 8876 11564 9604 11620
rect 7980 11218 8036 11228
rect 8428 11284 8484 11294
rect 7196 9826 7252 10332
rect 7196 9774 7198 9826
rect 7250 9774 7252 9826
rect 7196 9762 7252 9774
rect 7308 10052 7364 10062
rect 7308 9826 7364 9996
rect 7420 9940 7476 10780
rect 7756 10770 7812 10780
rect 8428 10666 8484 11228
rect 7532 10610 7588 10622
rect 8204 10612 8260 10622
rect 7532 10558 7534 10610
rect 7586 10558 7588 10610
rect 7532 10052 7588 10558
rect 7644 10610 8260 10612
rect 7644 10558 8206 10610
rect 8258 10558 8260 10610
rect 8428 10614 8430 10666
rect 8482 10614 8484 10666
rect 8428 10602 8484 10614
rect 8876 10610 8932 11564
rect 7644 10556 8260 10558
rect 7644 10442 7700 10556
rect 8204 10546 8260 10556
rect 8876 10558 8878 10610
rect 8930 10558 8932 10610
rect 8876 10546 8932 10558
rect 7644 10390 7646 10442
rect 7698 10390 7700 10442
rect 7644 10378 7700 10390
rect 8652 10498 8708 10510
rect 8652 10446 8654 10498
rect 8706 10446 8708 10498
rect 7532 9986 7588 9996
rect 7644 10276 7700 10286
rect 7420 9874 7476 9884
rect 7308 9774 7310 9826
rect 7362 9774 7364 9826
rect 7308 9762 7364 9774
rect 7532 9828 7588 9838
rect 7644 9828 7700 10220
rect 7532 9826 7700 9828
rect 7532 9774 7534 9826
rect 7586 9774 7700 9826
rect 7532 9772 7700 9774
rect 8652 9828 8708 10446
rect 7532 9762 7588 9772
rect 8652 9762 8708 9772
rect 7812 9716 7868 9726
rect 7812 9714 7924 9716
rect 7812 9662 7814 9714
rect 7866 9662 7924 9714
rect 7812 9650 7924 9662
rect 7036 9436 7300 9446
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7036 9370 7300 9380
rect 5964 9212 6356 9268
rect 5740 8930 5796 8942
rect 5740 8878 5742 8930
rect 5794 8878 5796 8930
rect 5740 8484 5796 8878
rect 5852 8484 5908 8494
rect 5740 8482 5908 8484
rect 5740 8430 5854 8482
rect 5906 8430 5908 8482
rect 5740 8428 5908 8430
rect 5852 8418 5908 8428
rect 5964 8428 6020 9212
rect 7644 8932 7700 8942
rect 7644 8838 7700 8876
rect 7756 8820 7812 8830
rect 7756 8428 7812 8764
rect 5964 8372 6244 8428
rect 5516 8206 5518 8258
rect 5570 8206 5572 8258
rect 5516 8194 5572 8206
rect 6188 8258 6244 8372
rect 6188 8206 6190 8258
rect 6242 8206 6244 8258
rect 6188 8194 6244 8206
rect 6860 8372 6916 8382
rect 6860 8258 6916 8316
rect 6860 8206 6862 8258
rect 6914 8206 6916 8258
rect 6860 8194 6916 8206
rect 7532 8372 7588 8382
rect 6524 8036 6580 8046
rect 5180 7422 5182 7474
rect 5234 7422 5236 7474
rect 5180 7410 5236 7422
rect 5964 8034 6580 8036
rect 5964 7982 6526 8034
rect 6578 7982 6580 8034
rect 5964 7980 6580 7982
rect 5964 7474 6020 7980
rect 6524 7970 6580 7980
rect 7036 7868 7300 7878
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7036 7802 7300 7812
rect 5964 7422 5966 7474
rect 6018 7422 6020 7474
rect 5964 7410 6020 7422
rect 4124 7084 4388 7094
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4124 7018 4388 7028
rect 7532 6690 7588 8316
rect 7644 8372 7812 8428
rect 7644 8370 7700 8372
rect 7644 8318 7646 8370
rect 7698 8318 7700 8370
rect 7644 8306 7700 8318
rect 7868 7924 7924 9650
rect 8092 9042 8148 9054
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 8092 8596 8148 8990
rect 9548 9042 9604 11564
rect 9660 11396 9716 11406
rect 9772 11396 9828 11900
rect 9940 11890 9996 11900
rect 9948 11788 10212 11798
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 9948 11722 10212 11732
rect 9996 11396 10052 11406
rect 9772 11394 10052 11396
rect 9772 11342 9998 11394
rect 10050 11342 10052 11394
rect 9772 11340 10052 11342
rect 9660 11302 9716 11340
rect 9996 11330 10052 11340
rect 10108 11394 10164 11406
rect 10108 11342 10110 11394
rect 10162 11342 10164 11394
rect 9660 10612 9716 10622
rect 10108 10612 10164 11342
rect 9660 10610 10164 10612
rect 9660 10558 9662 10610
rect 9714 10558 10164 10610
rect 9660 10556 10164 10558
rect 9660 9940 9716 10556
rect 10444 10500 10500 10510
rect 10332 10498 10500 10500
rect 10332 10446 10446 10498
rect 10498 10446 10500 10498
rect 10332 10444 10500 10446
rect 9948 10220 10212 10230
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 9948 10154 10212 10164
rect 10332 10052 10388 10444
rect 10444 10434 10500 10444
rect 9996 9996 10388 10052
rect 9884 9940 9940 9950
rect 9660 9938 9828 9940
rect 9660 9886 9662 9938
rect 9714 9886 9828 9938
rect 9660 9884 9828 9886
rect 9660 9874 9716 9884
rect 9548 8990 9550 9042
rect 9602 8990 9604 9042
rect 9548 8978 9604 8990
rect 8092 8530 8148 8540
rect 9772 8372 9828 9884
rect 9884 9042 9940 9884
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9884 8978 9940 8990
rect 9996 8874 10052 9996
rect 10220 9828 10276 9838
rect 10220 9042 10276 9772
rect 10668 9798 10724 12348
rect 11116 12404 11172 14364
rect 11396 13748 11452 13758
rect 11564 13748 11620 13758
rect 11452 13746 11620 13748
rect 11452 13694 11566 13746
rect 11618 13694 11620 13746
rect 11452 13692 11620 13694
rect 11396 13654 11452 13692
rect 11564 13682 11620 13692
rect 11116 12338 11172 12348
rect 11788 13636 11844 13646
rect 11788 12205 11844 13580
rect 11900 12850 11956 12862
rect 11900 12798 11902 12850
rect 11954 12798 11956 12850
rect 11900 12292 11956 12798
rect 11900 12226 11956 12236
rect 11004 12180 11060 12190
rect 11788 12153 11790 12205
rect 11842 12153 11844 12205
rect 11788 12141 11844 12153
rect 11004 12086 11060 12124
rect 12012 12068 12068 15148
rect 13580 14644 13636 15484
rect 14476 15370 14532 15820
rect 14308 15330 14364 15342
rect 14308 15316 14310 15330
rect 14140 15278 14310 15316
rect 14362 15278 14364 15330
rect 14476 15318 14478 15370
rect 14530 15318 14532 15370
rect 14476 15306 14532 15318
rect 14140 15260 14364 15278
rect 13580 14586 13692 14644
rect 13020 14532 13076 14542
rect 13020 14438 13076 14476
rect 13580 14534 13638 14586
rect 13690 14534 13692 14586
rect 13580 14522 13692 14534
rect 14140 14530 14196 15260
rect 13468 14420 13524 14430
rect 13468 14326 13524 14364
rect 12684 14308 12740 14318
rect 12348 14306 12740 14308
rect 12348 14254 12686 14306
rect 12738 14254 12740 14306
rect 12348 14252 12740 14254
rect 12348 13746 12404 14252
rect 12684 14242 12740 14252
rect 12860 14140 13124 14150
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 12860 14074 13124 14084
rect 12348 13694 12350 13746
rect 12402 13694 12404 13746
rect 12348 13682 12404 13694
rect 13580 13524 13636 14522
rect 14140 14478 14142 14530
rect 14194 14478 14196 14530
rect 13468 13468 13636 13524
rect 13804 14420 13860 14430
rect 13356 13188 13412 13198
rect 12860 12572 13124 12582
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 12860 12506 13124 12516
rect 13356 12404 13412 13132
rect 13356 12310 13412 12348
rect 11246 11954 11302 11966
rect 11246 11902 11248 11954
rect 11300 11902 11302 11954
rect 11246 11732 11302 11902
rect 11246 11666 11302 11676
rect 10892 11396 10948 11406
rect 10892 11302 10948 11340
rect 10668 9746 10670 9798
rect 10722 9746 10724 9798
rect 11900 9828 11956 9838
rect 12012 9828 12068 12012
rect 12684 11732 12740 11742
rect 12348 10498 12404 10510
rect 12348 10446 12350 10498
rect 12402 10446 12404 10498
rect 12348 9940 12404 10446
rect 12348 9874 12404 9884
rect 11900 9826 12068 9828
rect 11900 9774 11902 9826
rect 11954 9774 12068 9826
rect 11900 9772 12068 9774
rect 11900 9762 11956 9772
rect 10668 9734 10724 9746
rect 12236 9604 12292 9614
rect 12684 9604 12740 11676
rect 12796 11282 12852 11294
rect 12796 11230 12798 11282
rect 12850 11230 12852 11282
rect 12796 11172 12852 11230
rect 12796 11106 12852 11116
rect 12860 11004 13124 11014
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 12860 10938 13124 10948
rect 13468 10722 13524 13468
rect 13468 10670 13470 10722
rect 13522 10670 13524 10722
rect 13468 9826 13524 10670
rect 13636 11172 13692 11182
rect 13636 10666 13692 11116
rect 13636 10614 13638 10666
rect 13690 10614 13692 10666
rect 13636 10602 13692 10614
rect 13468 9774 13470 9826
rect 13522 9774 13524 9826
rect 13636 9940 13692 9950
rect 13636 9882 13692 9884
rect 13636 9830 13638 9882
rect 13690 9830 13692 9882
rect 13636 9818 13692 9830
rect 13468 9762 13524 9774
rect 12236 9602 12404 9604
rect 12236 9550 12238 9602
rect 12290 9550 12404 9602
rect 12236 9548 12404 9550
rect 12684 9548 12796 9604
rect 12236 9538 12292 9548
rect 10220 8990 10222 9042
rect 10274 8990 10276 9042
rect 10220 8978 10276 8990
rect 11676 9044 11732 9054
rect 11994 9044 12050 9054
rect 11676 9042 12050 9044
rect 11676 8990 11678 9042
rect 11730 8990 11996 9042
rect 12048 8990 12050 9042
rect 11676 8988 12050 8990
rect 11676 8978 11732 8988
rect 11994 8978 12050 8988
rect 12236 9042 12292 9054
rect 12236 8990 12238 9042
rect 12290 8990 12292 9042
rect 9996 8822 9998 8874
rect 10050 8822 10052 8874
rect 9996 8810 10052 8822
rect 10556 8820 10612 8830
rect 11340 8820 11396 8830
rect 10556 8726 10612 8764
rect 10668 8818 11396 8820
rect 10668 8766 11342 8818
rect 11394 8766 11396 8818
rect 10668 8764 11396 8766
rect 9948 8652 10212 8662
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 9948 8586 10212 8596
rect 9772 8260 9828 8316
rect 10668 8370 10724 8764
rect 11340 8754 11396 8764
rect 10668 8318 10670 8370
rect 10722 8318 10724 8370
rect 10668 8306 10724 8318
rect 9884 8260 9940 8270
rect 9772 8258 9940 8260
rect 9772 8206 9886 8258
rect 9938 8206 9940 8258
rect 9772 8204 9940 8206
rect 9548 8146 9604 8158
rect 9548 8094 9550 8146
rect 9602 8094 9604 8146
rect 7868 7868 8036 7924
rect 7980 7476 8036 7868
rect 9548 7588 9604 8094
rect 9548 7522 9604 7532
rect 8204 7476 8260 7486
rect 7980 7474 8260 7476
rect 7980 7422 8206 7474
rect 8258 7422 8260 7474
rect 7980 7420 8260 7422
rect 8204 7410 8260 7420
rect 7868 7364 7924 7374
rect 7868 7270 7924 7308
rect 8540 7252 8596 7262
rect 8316 7250 8596 7252
rect 8316 7198 8542 7250
rect 8594 7198 8596 7250
rect 8316 7196 8596 7198
rect 8316 6802 8372 7196
rect 8540 7186 8596 7196
rect 8316 6750 8318 6802
rect 8370 6750 8372 6802
rect 8316 6738 8372 6750
rect 7532 6638 7534 6690
rect 7586 6638 7588 6690
rect 7532 6626 7588 6638
rect 7036 6300 7300 6310
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7036 6234 7300 6244
rect 4124 5516 4388 5526
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4124 5450 4388 5460
rect 9772 5122 9828 8204
rect 9884 8194 9940 8204
rect 12236 8148 12292 8990
rect 12348 8372 12404 9548
rect 12740 9098 12796 9548
rect 12860 9436 13124 9446
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 12860 9370 13124 9380
rect 12740 9046 12742 9098
rect 12794 9046 12796 9098
rect 12908 9156 12964 9166
rect 12908 9062 12964 9100
rect 13244 9156 13300 9166
rect 12740 9034 12796 9046
rect 12348 8306 12404 8316
rect 12572 8148 12628 8158
rect 12236 8146 12628 8148
rect 12236 8094 12574 8146
rect 12626 8094 12628 8146
rect 12236 8092 12628 8094
rect 11116 8036 11172 8046
rect 11116 7586 11172 7980
rect 11116 7534 11118 7586
rect 11170 7534 11172 7586
rect 11116 7522 11172 7534
rect 11676 8036 11732 8046
rect 11284 7418 11340 7430
rect 11284 7366 11286 7418
rect 11338 7366 11340 7418
rect 11284 7364 11340 7366
rect 11284 7298 11340 7308
rect 9948 7084 10212 7094
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 9948 7018 10212 7028
rect 10220 6692 10276 6702
rect 10220 6598 10276 6636
rect 11676 6690 11732 7980
rect 11788 7476 11844 7486
rect 12236 7476 12292 8092
rect 12572 8082 12628 8092
rect 12860 7868 13124 7878
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 12860 7802 13124 7812
rect 11788 7474 12292 7476
rect 11788 7422 11790 7474
rect 11842 7422 12292 7474
rect 11788 7420 12292 7422
rect 11788 7410 11844 7420
rect 12030 7252 12086 7262
rect 12030 7250 12516 7252
rect 12030 7198 12032 7250
rect 12084 7198 12516 7250
rect 12030 7196 12516 7198
rect 12030 7186 12086 7196
rect 11676 6638 11678 6690
rect 11730 6638 11732 6690
rect 11676 6626 11732 6638
rect 11844 6692 11900 6702
rect 11844 6598 11900 6636
rect 12348 6690 12404 6702
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 11228 5908 11284 5918
rect 11228 5814 11284 5852
rect 11770 5908 11826 5918
rect 11770 5814 11826 5852
rect 12012 5906 12068 5918
rect 12012 5854 12014 5906
rect 12066 5854 12068 5906
rect 10892 5684 10948 5694
rect 10556 5682 10948 5684
rect 10556 5630 10894 5682
rect 10946 5630 10948 5682
rect 10556 5628 10948 5630
rect 9948 5516 10212 5526
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 9948 5450 10212 5460
rect 10556 5234 10612 5628
rect 10892 5618 10948 5628
rect 10556 5182 10558 5234
rect 10610 5182 10612 5234
rect 10556 5170 10612 5182
rect 12012 5236 12068 5854
rect 12348 5236 12404 6638
rect 12460 6356 12516 7196
rect 12590 6580 12646 6590
rect 12590 6486 12646 6524
rect 12460 6300 12572 6356
rect 12516 5962 12572 6300
rect 12860 6300 13124 6310
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 12860 6234 13124 6244
rect 12516 5910 12518 5962
rect 12570 5910 12572 5962
rect 12684 6020 12740 6030
rect 12684 5926 12740 5964
rect 13244 6020 13300 9100
rect 13804 9156 13860 14364
rect 14140 13860 14196 14478
rect 14382 14532 14438 14542
rect 14382 14438 14438 14476
rect 14252 13860 14308 13870
rect 14140 13858 14308 13860
rect 14140 13806 14254 13858
rect 14306 13806 14308 13858
rect 14140 13804 14308 13806
rect 14252 13794 14308 13804
rect 14588 13748 14644 16044
rect 14700 15370 14756 16268
rect 14700 15318 14702 15370
rect 14754 15318 14756 15370
rect 14700 15306 14756 15318
rect 14364 13746 14644 13748
rect 14364 13694 14590 13746
rect 14642 13694 14644 13746
rect 14364 13692 14644 13694
rect 14084 12906 14140 12918
rect 13916 12850 13972 12862
rect 13916 12798 13918 12850
rect 13970 12798 13972 12850
rect 13916 11956 13972 12798
rect 14084 12854 14086 12906
rect 14138 12854 14140 12906
rect 14084 12404 14140 12854
rect 14084 12348 14308 12404
rect 13916 11890 13972 11900
rect 14252 10724 14308 12348
rect 14364 12178 14420 13692
rect 14588 13682 14644 13692
rect 14812 13524 14868 16492
rect 15772 16492 16036 16502
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 15772 16426 16036 16436
rect 17388 16324 17444 17612
rect 18172 17666 18228 17678
rect 18172 17614 18174 17666
rect 18226 17614 18228 17666
rect 18172 17106 18228 17614
rect 19292 17444 19348 19842
rect 19516 19124 19572 19134
rect 19516 19030 19572 19068
rect 19964 18450 20020 19964
rect 20356 20022 20358 20074
rect 20410 20022 20412 20074
rect 20524 20132 20580 22316
rect 20748 22306 20804 22316
rect 21084 22326 21140 22338
rect 21084 22274 21086 22326
rect 21138 22274 21140 22326
rect 20860 21588 20916 21598
rect 20860 21494 20916 21532
rect 21084 21028 21140 22274
rect 21084 20962 21140 20972
rect 20524 20038 20580 20076
rect 20636 20356 20692 20366
rect 20356 20010 20412 20022
rect 20636 20018 20692 20300
rect 20188 19926 20244 19964
rect 20636 19966 20638 20018
rect 20690 19966 20692 20018
rect 20636 19796 20692 19966
rect 21196 20020 21252 22430
rect 21532 22342 21588 22354
rect 21532 22290 21534 22342
rect 21586 22290 21588 22342
rect 21532 21700 21588 22290
rect 21532 21634 21588 21644
rect 21644 21476 21700 21486
rect 21532 21474 21700 21476
rect 21532 21422 21646 21474
rect 21698 21422 21700 21474
rect 21532 21420 21700 21422
rect 21532 21364 21588 21420
rect 21644 21410 21700 21420
rect 21476 21308 21588 21364
rect 21364 21028 21420 21038
rect 21476 21028 21532 21308
rect 21980 21252 22036 21262
rect 21596 21196 21860 21206
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21596 21130 21860 21140
rect 21476 20972 21588 21028
rect 21364 20934 21420 20972
rect 21532 20186 21588 20972
rect 21644 20802 21700 20814
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20356 21700 20750
rect 21868 20804 21924 20814
rect 21980 20804 22036 21196
rect 22204 20804 22260 20814
rect 21980 20802 22260 20804
rect 21980 20750 22206 20802
rect 22258 20750 22260 20802
rect 21980 20748 22260 20750
rect 21868 20710 21924 20748
rect 22204 20738 22260 20748
rect 21644 20290 21700 20300
rect 22876 20356 22932 23996
rect 24508 21980 24772 21990
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24508 21914 24772 21924
rect 23548 21474 23604 21486
rect 23548 21422 23550 21474
rect 23602 21422 23604 21474
rect 23080 20804 23136 20814
rect 23080 20710 23136 20748
rect 23324 20690 23380 20702
rect 23324 20638 23326 20690
rect 23378 20638 23380 20690
rect 23324 20356 23380 20638
rect 22876 20290 22932 20300
rect 22988 20300 23380 20356
rect 21532 20134 21534 20186
rect 21586 20134 21588 20186
rect 22316 20244 22372 20254
rect 22316 20242 22820 20244
rect 22316 20190 22318 20242
rect 22370 20190 22820 20242
rect 22316 20188 22820 20190
rect 22316 20178 22372 20188
rect 21532 20122 21588 20134
rect 21588 20047 21644 20059
rect 21308 20020 21364 20030
rect 21588 20020 21590 20047
rect 21196 20018 21364 20020
rect 21196 19966 21310 20018
rect 21362 19966 21364 20018
rect 21196 19964 21364 19966
rect 21308 19954 21364 19964
rect 21532 19995 21590 20020
rect 21642 19995 21644 20047
rect 21532 19964 21644 19995
rect 22764 20020 22820 20188
rect 22876 20020 22932 20030
rect 22764 20018 22932 20020
rect 20356 19740 20692 19796
rect 20916 19796 20972 19806
rect 21532 19796 21588 19964
rect 20916 19794 21588 19796
rect 20916 19742 20918 19794
rect 20970 19742 21588 19794
rect 20916 19740 21588 19742
rect 22652 19962 22708 19974
rect 22764 19966 22878 20018
rect 22930 19966 22932 20018
rect 22764 19964 22932 19966
rect 22652 19910 22654 19962
rect 22706 19910 22708 19962
rect 22876 19954 22932 19964
rect 22988 20020 23044 20300
rect 23548 20132 23604 21422
rect 24276 21476 24332 21486
rect 24276 21474 24388 21476
rect 24276 21422 24278 21474
rect 24330 21422 24388 21474
rect 24276 21410 24388 21422
rect 24332 20802 24388 21410
rect 24332 20750 24334 20802
rect 24386 20750 24388 20802
rect 24332 20692 24388 20750
rect 24332 20636 24948 20692
rect 23996 20580 24052 20590
rect 23996 20578 24388 20580
rect 23996 20526 23998 20578
rect 24050 20526 24388 20578
rect 23996 20524 24388 20526
rect 23996 20514 24052 20524
rect 23604 20076 23808 20132
rect 23548 20066 23604 20076
rect 23752 20074 23808 20076
rect 23752 20022 23754 20074
rect 23806 20022 23808 20074
rect 23752 20010 23808 20022
rect 22988 19954 23044 19964
rect 22652 19908 22708 19910
rect 20356 19460 20412 19740
rect 20916 19730 20972 19740
rect 21596 19628 21860 19638
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21596 19562 21860 19572
rect 20300 19458 20412 19460
rect 20300 19406 20358 19458
rect 20410 19406 20412 19458
rect 20300 19394 20412 19406
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19180 17388 19348 17444
rect 19404 17556 19460 17566
rect 18684 17276 18948 17286
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18684 17210 18948 17220
rect 18172 17054 18174 17106
rect 18226 17054 18228 17106
rect 18172 17042 18228 17054
rect 18508 17108 18564 17118
rect 18508 16882 18564 17052
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18508 16818 18564 16830
rect 17276 16322 17444 16324
rect 17276 16270 17390 16322
rect 17442 16270 17444 16322
rect 17276 16268 17444 16270
rect 16716 16070 16772 16082
rect 16716 16018 16718 16070
rect 16770 16018 16772 16070
rect 14962 15330 15018 15342
rect 14962 15278 14964 15330
rect 15016 15316 15018 15330
rect 15204 15316 15260 15326
rect 15484 15316 15540 15326
rect 15016 15278 15092 15316
rect 14962 15260 15092 15278
rect 14924 14420 14980 14430
rect 14924 13970 14980 14364
rect 14924 13918 14926 13970
rect 14978 13918 14980 13970
rect 14924 13906 14980 13918
rect 15036 14420 15092 15260
rect 15204 15314 15540 15316
rect 15204 15262 15206 15314
rect 15258 15262 15486 15314
rect 15538 15262 15540 15314
rect 15204 15260 15540 15262
rect 15204 15250 15260 15260
rect 15484 15250 15540 15260
rect 15820 15092 15876 15130
rect 15820 15026 15876 15036
rect 15772 14924 16036 14934
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 15772 14858 16036 14868
rect 16716 14868 16772 16018
rect 17276 15316 17332 16268
rect 17388 16258 17444 16268
rect 19180 15988 19236 17388
rect 19404 16882 19460 17500
rect 19404 16830 19406 16882
rect 19458 16830 19460 16882
rect 19404 16818 19460 16830
rect 19628 16897 19684 16909
rect 19628 16845 19630 16897
rect 19682 16845 19684 16897
rect 19628 16660 19684 16845
rect 19740 16884 19796 16894
rect 19964 16884 20020 18398
rect 20188 18618 20244 18630
rect 20188 18566 20190 18618
rect 20242 18566 20244 18618
rect 20188 18452 20244 18566
rect 20188 18386 20244 18396
rect 20300 18340 20356 19394
rect 22652 19358 22708 19852
rect 23996 19794 24052 19806
rect 23996 19742 23998 19794
rect 24050 19742 24052 19794
rect 21308 19346 21364 19358
rect 21308 19294 21310 19346
rect 21362 19294 21364 19346
rect 20636 19236 20692 19246
rect 20636 19142 20692 19180
rect 20860 19234 20916 19246
rect 20860 19182 20862 19234
rect 20914 19182 20916 19234
rect 20860 19124 20916 19182
rect 20860 19058 20916 19068
rect 21308 18900 21364 19294
rect 22596 19346 22708 19358
rect 22596 19294 22598 19346
rect 22650 19294 22708 19346
rect 22596 19292 22708 19294
rect 22876 19684 22932 19694
rect 22596 19282 22652 19292
rect 20412 18844 21364 18900
rect 21420 19236 21476 19268
rect 21420 19138 21422 19180
rect 21474 19138 21476 19180
rect 21756 19236 21812 19246
rect 21756 19142 21812 19180
rect 20412 18506 20468 18844
rect 20412 18454 20414 18506
rect 20466 18454 20468 18506
rect 20412 18442 20468 18454
rect 20636 18450 20692 18462
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20636 18340 20692 18398
rect 20300 18284 20692 18340
rect 20076 17556 20132 17566
rect 20076 17462 20132 17500
rect 20188 17108 20244 17118
rect 21420 17052 21476 19138
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22036 18340 22092 18350
rect 22036 18246 22092 18284
rect 22764 18340 22820 18398
rect 22876 18452 22932 19628
rect 23996 19684 24052 19742
rect 23996 19618 24052 19628
rect 23436 19572 23492 19582
rect 23231 19236 23287 19246
rect 23231 19142 23287 19180
rect 22988 19124 23044 19134
rect 22988 19122 23156 19124
rect 22988 19070 22990 19122
rect 23042 19070 23156 19122
rect 22988 19068 23156 19070
rect 22988 19058 23044 19068
rect 22988 18452 23044 18462
rect 22876 18450 23044 18452
rect 22876 18398 22990 18450
rect 23042 18398 23044 18450
rect 22876 18396 23044 18398
rect 22988 18386 23044 18396
rect 23100 18452 23156 19068
rect 23436 18506 23492 19516
rect 24108 19236 24164 19246
rect 24332 19236 24388 20524
rect 24508 20412 24772 20422
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24508 20346 24772 20356
rect 24892 20020 24948 20636
rect 24892 19954 24948 19964
rect 24108 19234 24388 19236
rect 24108 19182 24110 19234
rect 24162 19182 24388 19234
rect 24108 19180 24388 19182
rect 24108 19170 24164 19180
rect 24508 18844 24772 18854
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24508 18778 24772 18788
rect 23436 18454 23438 18506
rect 23490 18454 23492 18506
rect 23436 18442 23492 18454
rect 23660 18452 23716 18462
rect 23996 18452 24052 18462
rect 23660 18450 23940 18452
rect 23100 18386 23156 18396
rect 23660 18398 23662 18450
rect 23714 18398 23940 18450
rect 23660 18396 23940 18398
rect 23660 18386 23716 18396
rect 22428 18226 22484 18238
rect 22428 18174 22430 18226
rect 22482 18174 22484 18226
rect 22428 18116 22484 18174
rect 21596 18060 21860 18070
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 22428 18050 22484 18060
rect 21596 17994 21860 18004
rect 22764 18004 22820 18284
rect 22764 17938 22820 17948
rect 23324 18338 23380 18350
rect 23324 18286 23326 18338
rect 23378 18286 23380 18338
rect 22092 17668 22148 17678
rect 22092 17574 22148 17612
rect 22968 17610 23024 17622
rect 22204 17556 22260 17566
rect 21532 17052 21588 17062
rect 20188 17050 20244 17052
rect 20188 16998 20190 17050
rect 20242 16998 20244 17050
rect 20188 16986 20244 16998
rect 20748 17050 21588 17052
rect 20748 16998 21534 17050
rect 21586 16998 21588 17050
rect 20748 16996 21588 16998
rect 20412 16909 20468 16922
rect 20076 16884 20132 16894
rect 19740 16770 19796 16828
rect 19740 16718 19742 16770
rect 19794 16718 19796 16770
rect 19740 16706 19796 16718
rect 19852 16882 20132 16884
rect 19852 16830 20078 16882
rect 20130 16830 20132 16882
rect 19852 16828 20132 16830
rect 19628 16594 19684 16604
rect 19292 16100 19348 16110
rect 19292 16006 19348 16044
rect 19628 16100 19684 16110
rect 19852 16100 19908 16828
rect 20076 16818 20132 16828
rect 20412 16884 20414 16909
rect 20466 16884 20468 16909
rect 20412 16818 20468 16828
rect 20748 16882 20804 16996
rect 21532 16986 21588 16996
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20748 16818 20804 16830
rect 21756 16882 21812 16894
rect 21756 16830 21758 16882
rect 21810 16830 21812 16882
rect 19628 16098 19908 16100
rect 19628 16046 19630 16098
rect 19682 16046 19908 16098
rect 19628 16044 19908 16046
rect 20076 16660 20132 16670
rect 21756 16660 21812 16830
rect 22204 16884 22260 17500
rect 22968 17558 22970 17610
rect 23022 17558 23024 17610
rect 22968 17556 23024 17558
rect 22968 17490 23024 17500
rect 23212 17554 23268 17566
rect 23212 17502 23214 17554
rect 23266 17502 23268 17554
rect 23100 17050 23156 17062
rect 23100 16998 23102 17050
rect 23154 16998 23156 17050
rect 23100 16996 23156 16998
rect 23100 16930 23156 16940
rect 22316 16884 22372 16894
rect 22204 16882 22372 16884
rect 22204 16830 22318 16882
rect 22370 16830 22372 16882
rect 22204 16828 22372 16830
rect 22316 16818 22372 16828
rect 22988 16882 23044 16894
rect 22988 16830 22990 16882
rect 23042 16830 23044 16882
rect 22988 16660 23044 16830
rect 21756 16604 22036 16660
rect 20076 16100 20132 16604
rect 21596 16492 21860 16502
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21596 16426 21860 16436
rect 20636 16100 20692 16110
rect 20076 16098 20244 16100
rect 20076 16046 20078 16098
rect 20130 16046 20244 16098
rect 20076 16044 20244 16046
rect 19628 16034 19684 16044
rect 20076 16034 20132 16044
rect 18684 15708 18948 15718
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18684 15642 18948 15652
rect 17276 15314 17892 15316
rect 17276 15262 17278 15314
rect 17330 15262 17892 15314
rect 17276 15260 17892 15262
rect 17276 15250 17332 15260
rect 17052 15092 17108 15102
rect 16716 14812 16884 14868
rect 15148 14420 15204 14430
rect 15036 14418 15204 14420
rect 15036 14366 15150 14418
rect 15202 14366 15204 14418
rect 15036 14364 15204 14366
rect 14588 13468 14868 13524
rect 14588 13076 14644 13468
rect 14588 12962 14644 13020
rect 14588 12910 14590 12962
rect 14642 12910 14644 12962
rect 14588 12898 14644 12910
rect 14830 12852 14886 12862
rect 14830 12758 14886 12796
rect 14364 12126 14366 12178
rect 14418 12126 14420 12178
rect 14364 12114 14420 12126
rect 15036 12180 15092 14364
rect 15148 14354 15204 14364
rect 16828 14308 16884 14812
rect 17052 14642 17108 15036
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14578 17108 14590
rect 17836 14532 17892 15260
rect 18060 15202 18116 15214
rect 18060 15150 18062 15202
rect 18114 15150 18116 15202
rect 18060 14756 18116 15150
rect 18508 14980 18564 14990
rect 18172 14756 18228 14766
rect 18060 14754 18228 14756
rect 18060 14702 18174 14754
rect 18226 14702 18228 14754
rect 18060 14700 18228 14702
rect 18172 14690 18228 14700
rect 17836 14530 18116 14532
rect 17836 14478 17838 14530
rect 17890 14478 18116 14530
rect 17836 14476 18116 14478
rect 17836 14466 17892 14476
rect 16716 14252 16884 14308
rect 15772 13356 16036 13366
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 15772 13290 16036 13300
rect 16716 13300 16772 14252
rect 18060 13748 18116 14476
rect 18508 14530 18564 14924
rect 18508 14478 18510 14530
rect 18562 14478 18564 14530
rect 18508 14466 18564 14478
rect 18684 14140 18948 14150
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18684 14074 18948 14084
rect 18172 13748 18228 13758
rect 18060 13746 18228 13748
rect 18060 13694 18174 13746
rect 18226 13694 18228 13746
rect 18060 13692 18228 13694
rect 18172 13682 18228 13692
rect 18956 13634 19012 13646
rect 18956 13582 18958 13634
rect 19010 13582 19012 13634
rect 16716 13234 16772 13244
rect 17724 13300 17780 13310
rect 15372 13076 15428 13086
rect 15372 12982 15428 13020
rect 17276 12962 17332 12974
rect 17276 12910 17278 12962
rect 17330 12910 17332 12962
rect 15036 12114 15092 12124
rect 15596 12852 15652 12862
rect 15596 12178 15652 12796
rect 15932 12404 15988 12414
rect 15932 12310 15988 12348
rect 17276 12404 17332 12910
rect 17276 12338 17332 12348
rect 15596 12126 15598 12178
rect 15650 12126 15652 12178
rect 15596 12114 15652 12126
rect 14700 11956 14756 11966
rect 14700 11508 14756 11900
rect 15772 11788 16036 11798
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 15772 11722 16036 11732
rect 14700 11452 14980 11508
rect 14756 11338 14812 11350
rect 14756 11286 14758 11338
rect 14810 11286 14812 11338
rect 14382 10724 14438 10734
rect 14756 10724 14812 11286
rect 14252 10722 14438 10724
rect 14252 10670 14384 10722
rect 14436 10670 14438 10722
rect 14252 10668 14438 10670
rect 14382 10658 14438 10668
rect 14588 10668 14812 10724
rect 14924 11226 14980 11452
rect 14924 11174 14926 11226
rect 14978 11174 14980 11226
rect 14140 10612 14196 10622
rect 14140 10518 14196 10556
rect 14588 10164 14644 10668
rect 14924 10612 14980 11174
rect 14382 10108 14644 10164
rect 14812 10556 14980 10612
rect 15260 11394 15316 11406
rect 15260 11342 15262 11394
rect 15314 11342 15316 11394
rect 15260 11284 15316 11342
rect 15260 10612 15316 11228
rect 15502 11284 15558 11294
rect 16044 11284 16100 11294
rect 15502 11282 15988 11284
rect 15502 11230 15504 11282
rect 15556 11230 15988 11282
rect 15502 11228 15988 11230
rect 15502 11218 15558 11228
rect 14382 10050 14438 10108
rect 14382 9998 14384 10050
rect 14436 9998 14438 10050
rect 14382 9986 14438 9998
rect 14140 9828 14196 9838
rect 14140 9734 14196 9772
rect 14812 9714 14868 10556
rect 15260 10546 15316 10556
rect 15932 10610 15988 11228
rect 16044 11190 16100 11228
rect 16268 10836 16324 10846
rect 16268 10742 16324 10780
rect 15932 10558 15934 10610
rect 15986 10558 15988 10610
rect 17724 10637 17780 13244
rect 18956 13188 19012 13582
rect 19068 13188 19124 13198
rect 18956 13186 19124 13188
rect 18956 13134 19070 13186
rect 19122 13134 19124 13186
rect 18956 13132 19124 13134
rect 19068 13122 19124 13132
rect 18060 12964 18116 12974
rect 19180 12964 19236 15932
rect 20076 15930 20132 15942
rect 20076 15878 20078 15930
rect 20130 15878 20132 15930
rect 19964 15316 20020 15326
rect 19964 15222 20020 15260
rect 20076 15204 20132 15878
rect 20188 15428 20244 16044
rect 20188 15362 20244 15372
rect 20412 16042 20468 16054
rect 20412 15990 20414 16042
rect 20466 15990 20468 16042
rect 20636 16006 20692 16044
rect 21084 16100 21140 16110
rect 20076 15138 20132 15148
rect 20412 15202 20468 15990
rect 20412 15150 20414 15202
rect 20466 15150 20468 15202
rect 20412 15138 20468 15150
rect 20524 15329 20580 15341
rect 20524 15277 20526 15329
rect 20578 15277 20580 15329
rect 20356 14756 20412 14766
rect 20356 14662 20412 14700
rect 20524 14756 20580 15277
rect 20860 15316 20916 15326
rect 20860 15222 20916 15260
rect 20524 14690 20580 14700
rect 21084 14644 21140 16044
rect 21756 16100 21812 16110
rect 21252 15428 21308 15438
rect 21252 15334 21308 15372
rect 21532 15314 21588 15326
rect 21532 15262 21534 15314
rect 21586 15262 21588 15314
rect 21532 15148 21588 15262
rect 21756 15316 21812 16044
rect 21980 15876 22036 16604
rect 22652 16604 23044 16660
rect 21980 15810 22036 15820
rect 22428 16100 22484 16110
rect 21756 15222 21812 15260
rect 21420 15092 21588 15148
rect 21420 14756 21476 15092
rect 22428 14980 22484 16044
rect 22540 15986 22596 15998
rect 22540 15934 22542 15986
rect 22594 15934 22596 15986
rect 22540 15316 22596 15934
rect 22540 15250 22596 15260
rect 22652 15204 22708 16604
rect 23212 16548 23268 17502
rect 23324 16938 23380 18286
rect 23884 17668 23940 18396
rect 23996 18358 24052 18396
rect 23884 17612 24164 17668
rect 23996 17444 24052 17454
rect 23324 16886 23326 16938
rect 23378 16886 23380 16938
rect 23884 17442 24052 17444
rect 23884 17390 23998 17442
rect 24050 17390 24052 17442
rect 23884 17388 24052 17390
rect 23324 16874 23380 16886
rect 23660 16884 23716 16894
rect 23660 16790 23716 16828
rect 22988 16492 23268 16548
rect 22783 16100 22839 16138
rect 22783 16034 22839 16044
rect 22652 15138 22708 15148
rect 22764 15876 22820 15886
rect 21596 14924 21860 14934
rect 22428 14924 22708 14980
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21596 14858 21860 14868
rect 21084 14588 21364 14644
rect 20636 14530 20692 14542
rect 20636 14478 20638 14530
rect 20690 14478 20692 14530
rect 20636 13636 20692 14478
rect 20860 14530 20916 14542
rect 20860 14478 20862 14530
rect 20914 14478 20916 14530
rect 20860 13748 20916 14478
rect 20860 13654 20916 13692
rect 20636 13570 20692 13580
rect 18060 12962 18452 12964
rect 18060 12910 18062 12962
rect 18114 12910 18452 12962
rect 18060 12908 18452 12910
rect 18060 12898 18116 12908
rect 18396 12178 18452 12908
rect 19068 12908 19236 12964
rect 19404 13412 19460 13422
rect 19404 12962 19460 13356
rect 19404 12910 19406 12962
rect 19458 12910 19460 12962
rect 18684 12572 18948 12582
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18684 12506 18948 12516
rect 18396 12126 18398 12178
rect 18450 12126 18452 12178
rect 17948 11394 18004 11406
rect 17948 11342 17950 11394
rect 18002 11342 18004 11394
rect 17948 10836 18004 11342
rect 18396 11396 18452 12126
rect 19068 11844 19124 12908
rect 19404 12898 19460 12910
rect 21084 12852 21140 12862
rect 21084 12290 21140 12796
rect 21084 12238 21086 12290
rect 21138 12238 21140 12290
rect 21084 12226 21140 12238
rect 21196 12180 21252 14588
rect 21308 14530 21364 14588
rect 21308 14478 21310 14530
rect 21362 14478 21364 14530
rect 21308 14466 21364 14478
rect 21420 14532 21476 14700
rect 21980 14532 22036 14542
rect 21420 14476 21644 14532
rect 21588 14474 21644 14476
rect 21588 14422 21590 14474
rect 21642 14422 21644 14474
rect 21588 14410 21644 14422
rect 21756 14530 22036 14532
rect 21756 14478 21982 14530
rect 22034 14478 22036 14530
rect 21756 14476 22036 14478
rect 21420 14362 21476 14374
rect 21420 14310 21422 14362
rect 21474 14310 21476 14362
rect 21308 13748 21364 13758
rect 21308 13654 21364 13692
rect 21420 13524 21476 14310
rect 21644 13761 21700 13773
rect 21644 13709 21646 13761
rect 21698 13709 21700 13761
rect 21644 13636 21700 13709
rect 21644 13570 21700 13580
rect 21756 13634 21812 14476
rect 21980 14466 22036 14476
rect 22652 13802 22708 14924
rect 22428 13748 22484 13758
rect 21756 13582 21758 13634
rect 21810 13582 21812 13634
rect 21756 13570 21812 13582
rect 22204 13746 22484 13748
rect 22204 13694 22430 13746
rect 22482 13694 22484 13746
rect 22652 13750 22654 13802
rect 22706 13750 22708 13802
rect 22652 13738 22708 13750
rect 22204 13692 22484 13694
rect 22204 13636 22260 13692
rect 22428 13682 22484 13692
rect 21420 13458 21476 13468
rect 21596 13356 21860 13366
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21596 13290 21860 13300
rect 22204 12516 22260 13580
rect 22764 13634 22820 15820
rect 22988 15428 23044 16492
rect 23660 16100 23716 16110
rect 23884 16100 23940 17388
rect 23996 17378 24052 17388
rect 23660 16098 23940 16100
rect 23660 16046 23662 16098
rect 23714 16046 23940 16098
rect 23660 16044 23940 16046
rect 23660 16034 23716 16044
rect 22988 15372 23212 15428
rect 23156 15370 23212 15372
rect 22764 13582 22766 13634
rect 22818 13582 22820 13634
rect 22764 13570 22820 13582
rect 22876 15314 22932 15326
rect 22876 15262 22878 15314
rect 22930 15262 22932 15314
rect 23156 15318 23158 15370
rect 23210 15318 23212 15370
rect 23156 15306 23212 15318
rect 23548 15316 23604 15326
rect 22876 13412 22932 15262
rect 22988 15204 23044 15242
rect 23548 15222 23604 15260
rect 23884 15314 23940 15326
rect 23884 15262 23886 15314
rect 23938 15262 23940 15314
rect 22988 15138 23044 15148
rect 23212 15204 23268 15214
rect 23100 14756 23156 14766
rect 23212 14756 23268 15148
rect 23884 15148 23940 15262
rect 24108 15204 24164 17612
rect 24332 17666 24388 17678
rect 24332 17614 24334 17666
rect 24386 17614 24388 17666
rect 24332 15998 24388 17614
rect 24508 17276 24772 17286
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24508 17210 24772 17220
rect 24276 15988 24388 15998
rect 24332 15932 24388 15988
rect 25004 16884 25060 16894
rect 24276 15894 24332 15932
rect 24508 15708 24772 15718
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24508 15642 24772 15652
rect 23884 15092 24052 15148
rect 24108 15138 24164 15148
rect 23996 14980 24052 15092
rect 23996 14924 24948 14980
rect 23100 14754 23268 14756
rect 23100 14702 23102 14754
rect 23154 14702 23268 14754
rect 23100 14700 23268 14702
rect 23100 14690 23156 14700
rect 24220 14530 24276 14542
rect 23343 14474 23399 14486
rect 23343 14422 23345 14474
rect 23397 14422 23399 14474
rect 23343 14084 23399 14422
rect 23100 14028 23399 14084
rect 24220 14478 24222 14530
rect 24274 14478 24276 14530
rect 23100 13748 23156 14028
rect 23604 13972 23660 13982
rect 23604 13878 23660 13916
rect 23772 13972 23828 13982
rect 23100 13654 23156 13692
rect 23772 13746 23828 13916
rect 24108 13972 24164 13982
rect 24220 13972 24276 14478
rect 24508 14140 24772 14150
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24508 14074 24772 14084
rect 24108 13970 24276 13972
rect 24108 13918 24110 13970
rect 24162 13918 24276 13970
rect 24108 13916 24276 13918
rect 24108 13906 24164 13916
rect 23772 13694 23774 13746
rect 23826 13694 23828 13746
rect 23772 13682 23828 13694
rect 22316 13356 22932 13412
rect 22316 13186 22372 13356
rect 22316 13134 22318 13186
rect 22370 13134 22372 13186
rect 22316 13122 22372 13134
rect 23436 12964 23492 12974
rect 21980 12460 22260 12516
rect 22559 12906 22615 12918
rect 22559 12854 22561 12906
rect 22613 12854 22615 12906
rect 23436 12870 23492 12908
rect 23996 12964 24052 12974
rect 23996 12870 24052 12908
rect 24332 12962 24388 12974
rect 24332 12910 24334 12962
rect 24386 12910 24388 12962
rect 22559 12852 22615 12854
rect 22559 12516 22615 12796
rect 22559 12460 23044 12516
rect 21980 12234 22036 12460
rect 22204 12404 22260 12460
rect 21532 12180 21588 12190
rect 21196 12178 21588 12180
rect 21196 12126 21534 12178
rect 21586 12126 21588 12178
rect 21980 12182 21982 12234
rect 22034 12182 22036 12234
rect 21980 12170 22036 12182
rect 22092 12346 22148 12358
rect 22204 12348 22932 12404
rect 22092 12294 22094 12346
rect 22146 12294 22148 12346
rect 21196 12124 21588 12126
rect 19180 12068 19236 12078
rect 19180 12066 19460 12068
rect 19180 12014 19182 12066
rect 19234 12014 19460 12066
rect 19180 12012 19460 12014
rect 19180 12002 19236 12012
rect 19068 11788 19348 11844
rect 18732 11396 18788 11406
rect 18396 11394 18788 11396
rect 18396 11342 18734 11394
rect 18786 11342 18788 11394
rect 18396 11340 18788 11342
rect 17948 10770 18004 10780
rect 18508 10836 18564 11340
rect 18732 11330 18788 11340
rect 18684 11004 18948 11014
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18684 10938 18948 10948
rect 18732 10836 18788 10846
rect 18508 10834 19236 10836
rect 18508 10782 18734 10834
rect 18786 10782 19236 10834
rect 18508 10780 19236 10782
rect 17724 10585 17726 10637
rect 17778 10585 17780 10637
rect 17724 10573 17780 10585
rect 15932 10546 15988 10558
rect 15772 10220 16036 10230
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 15772 10154 16036 10164
rect 15484 9828 15540 9838
rect 14812 9662 14814 9714
rect 14866 9662 14868 9714
rect 14812 9604 14868 9662
rect 13804 9090 13860 9100
rect 14140 9548 14868 9604
rect 14980 9770 15036 9782
rect 14980 9718 14982 9770
rect 15034 9718 15036 9770
rect 15484 9734 15540 9772
rect 16492 9828 16548 9838
rect 16492 9734 16548 9772
rect 18396 9826 18452 9838
rect 18396 9774 18398 9826
rect 18450 9774 18452 9826
rect 13580 9042 13636 9054
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8428 13636 8990
rect 13748 8986 13804 8998
rect 13748 8934 13750 8986
rect 13802 8934 13804 8986
rect 13748 8932 13804 8934
rect 13748 8866 13804 8876
rect 13468 8372 13636 8428
rect 13468 7586 13524 8316
rect 14140 8260 14196 9548
rect 14980 9268 15036 9718
rect 15726 9716 15782 9726
rect 14494 9212 15036 9268
rect 15708 9714 15782 9716
rect 15708 9662 15728 9714
rect 15780 9662 15782 9714
rect 15708 9650 15782 9662
rect 14494 9154 14550 9212
rect 14494 9102 14496 9154
rect 14548 9102 14550 9154
rect 14494 9090 14550 9102
rect 14252 9042 14308 9054
rect 14252 8990 14254 9042
rect 14306 8990 14308 9042
rect 14252 8428 14308 8990
rect 15708 9044 15764 9650
rect 16604 9268 16660 9278
rect 16604 9174 16660 9212
rect 18396 9268 18452 9774
rect 18396 9202 18452 9212
rect 16268 9044 16324 9054
rect 15708 9042 16324 9044
rect 15708 8990 16270 9042
rect 16322 8990 16324 9042
rect 15708 8988 16324 8990
rect 16268 8978 16324 8988
rect 15772 8652 16036 8662
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 15772 8586 16036 8596
rect 18508 8428 18564 10780
rect 18732 10770 18788 10780
rect 19180 9826 19236 10780
rect 19180 9774 19182 9826
rect 19234 9774 19236 9826
rect 19180 9604 19236 9774
rect 19292 9828 19348 11788
rect 19404 11620 19460 12012
rect 19852 11844 19908 11854
rect 19516 11620 19572 11630
rect 19404 11618 19572 11620
rect 19404 11566 19518 11618
rect 19570 11566 19572 11618
rect 19404 11564 19572 11566
rect 19516 11554 19572 11564
rect 19852 11394 19908 11788
rect 19852 11342 19854 11394
rect 19906 11342 19908 11394
rect 19852 11330 19908 11342
rect 21308 11394 21364 12124
rect 21532 12114 21588 12124
rect 22092 12068 22148 12294
rect 22876 12346 22932 12348
rect 22876 12294 22878 12346
rect 22930 12294 22932 12346
rect 22876 12282 22932 12294
rect 22092 12002 22148 12012
rect 22204 12178 22260 12190
rect 22204 12126 22206 12178
rect 22258 12126 22260 12178
rect 21596 11788 21860 11798
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21596 11722 21860 11732
rect 21308 11342 21310 11394
rect 21362 11342 21364 11394
rect 21308 11330 21364 11342
rect 21756 11508 21812 11518
rect 22204 11508 22260 12126
rect 22876 12178 22932 12190
rect 22876 12126 22878 12178
rect 22930 12126 22932 12178
rect 22876 11620 22932 12126
rect 22876 11554 22932 11564
rect 22988 12180 23044 12460
rect 24052 12346 24108 12358
rect 23212 12292 23268 12302
rect 23212 12234 23268 12236
rect 23212 12182 23214 12234
rect 23266 12182 23268 12234
rect 24052 12294 24054 12346
rect 24106 12294 24108 12346
rect 24052 12292 24108 12294
rect 24052 12226 24108 12236
rect 23212 12170 23268 12182
rect 23436 12178 23492 12190
rect 22540 11508 22596 11518
rect 22204 11506 22596 11508
rect 22204 11454 22542 11506
rect 22594 11454 22596 11506
rect 22204 11452 22596 11454
rect 21756 11355 21812 11452
rect 22540 11442 22596 11452
rect 22652 11508 22708 11518
rect 21756 11303 21758 11355
rect 21810 11303 21812 11355
rect 21980 11396 22036 11406
rect 21980 11394 22484 11396
rect 21980 11342 21982 11394
rect 22034 11342 22484 11394
rect 21980 11340 22484 11342
rect 21980 11330 22036 11340
rect 21756 11291 21812 11303
rect 21532 11226 21588 11238
rect 21532 11174 21534 11226
rect 21586 11174 21588 11226
rect 21532 10948 21588 11174
rect 21532 10892 21812 10948
rect 21756 10610 21812 10892
rect 22428 10724 22484 11340
rect 22652 11379 22708 11452
rect 22652 11327 22654 11379
rect 22706 11327 22708 11379
rect 22876 11396 22932 11406
rect 22988 11396 23044 12124
rect 23436 12126 23438 12178
rect 23490 12126 23492 12178
rect 23324 11508 23380 11518
rect 23324 11414 23380 11452
rect 22876 11394 23044 11396
rect 22876 11342 22878 11394
rect 22930 11342 23044 11394
rect 22876 11340 23044 11342
rect 23436 11350 23492 12126
rect 23884 12180 23940 12190
rect 23884 12086 23940 12124
rect 24332 11966 24388 12910
rect 24508 12572 24772 12582
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24508 12506 24772 12516
rect 24276 11956 24388 11966
rect 24332 11900 24388 11956
rect 23660 11620 23716 11630
rect 23660 11396 23716 11564
rect 24276 11506 24332 11900
rect 24276 11454 24278 11506
rect 24330 11454 24332 11506
rect 24276 11442 24332 11454
rect 22876 11330 22932 11340
rect 22652 11315 22708 11327
rect 23436 11298 23438 11350
rect 23490 11298 23492 11350
rect 23436 11284 23492 11298
rect 22988 11228 23492 11284
rect 23548 11394 23716 11396
rect 23548 11342 23662 11394
rect 23714 11342 23716 11394
rect 23548 11340 23716 11342
rect 22596 10724 22652 10734
rect 22428 10722 22652 10724
rect 22428 10670 22598 10722
rect 22650 10670 22652 10722
rect 22428 10668 22652 10670
rect 22596 10658 22652 10668
rect 21756 10558 21758 10610
rect 21810 10558 21812 10610
rect 21756 10546 21812 10558
rect 22876 10610 22932 10622
rect 22876 10558 22878 10610
rect 22930 10558 22932 10610
rect 22260 10498 22316 10510
rect 22260 10446 22262 10498
rect 22314 10446 22316 10498
rect 21420 10386 21476 10398
rect 21420 10334 21422 10386
rect 21474 10334 21476 10386
rect 21420 9940 21476 10334
rect 21596 10220 21860 10230
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21596 10154 21860 10164
rect 22260 10164 22316 10446
rect 22876 10388 22932 10558
rect 22988 10388 23044 11228
rect 23548 11172 23604 11340
rect 23660 11330 23716 11340
rect 23380 11116 23604 11172
rect 23380 10836 23436 11116
rect 24508 11004 24772 11014
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24508 10938 24772 10948
rect 23100 10834 23436 10836
rect 23100 10782 23382 10834
rect 23434 10782 23436 10834
rect 23100 10780 23436 10782
rect 23100 10610 23156 10780
rect 23380 10770 23436 10780
rect 23100 10558 23102 10610
rect 23154 10558 23156 10610
rect 23100 10546 23156 10558
rect 23548 10610 23604 10622
rect 23548 10558 23550 10610
rect 23602 10558 23604 10610
rect 22876 10332 23156 10388
rect 22260 10098 22316 10108
rect 21420 9874 21476 9884
rect 21980 9940 22036 9950
rect 21980 9846 22036 9884
rect 19852 9828 19908 9838
rect 19292 9826 19908 9828
rect 19292 9774 19854 9826
rect 19906 9774 19908 9826
rect 19292 9772 19908 9774
rect 19180 9538 19236 9548
rect 18684 9436 18948 9446
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18684 9370 18948 9380
rect 19124 9268 19180 9278
rect 19404 9268 19460 9772
rect 19852 9762 19908 9772
rect 21196 9826 21252 9838
rect 21196 9774 21198 9826
rect 21250 9774 21252 9826
rect 19124 9266 19460 9268
rect 19124 9214 19126 9266
rect 19178 9214 19460 9266
rect 19124 9212 19460 9214
rect 19516 9602 19572 9614
rect 19516 9550 19518 9602
rect 19570 9550 19572 9602
rect 19124 9202 19180 9212
rect 14252 8372 14420 8428
rect 14364 8306 14420 8316
rect 14924 8372 14980 8382
rect 14252 8260 14308 8270
rect 14140 8258 14308 8260
rect 14140 8206 14254 8258
rect 14306 8206 14308 8258
rect 14924 8258 14980 8316
rect 15708 8372 15764 8382
rect 15708 8278 15764 8316
rect 18396 8372 18564 8428
rect 19516 8428 19572 9550
rect 21196 9604 21252 9774
rect 23100 9604 23156 10332
rect 21196 9538 21252 9548
rect 22540 9548 23156 9604
rect 23343 9604 23399 9614
rect 21596 8652 21860 8662
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21596 8586 21860 8596
rect 19516 8372 19796 8428
rect 14140 8204 14308 8206
rect 14252 8194 14308 8204
rect 14420 8202 14476 8214
rect 14420 8150 14422 8202
rect 14474 8150 14476 8202
rect 14924 8206 14926 8258
rect 14978 8206 14980 8258
rect 14924 8194 14980 8206
rect 17612 8258 17668 8270
rect 17612 8206 17614 8258
rect 17666 8206 17668 8258
rect 14420 7598 14476 8150
rect 15166 8146 15222 8158
rect 15166 8094 15168 8146
rect 15220 8094 15222 8146
rect 15166 7812 15222 8094
rect 15166 7756 15876 7812
rect 13468 7534 13470 7586
rect 13522 7534 13524 7586
rect 13468 7522 13524 7534
rect 13636 7588 13692 7598
rect 13636 7530 13692 7532
rect 13636 7478 13638 7530
rect 13690 7478 13692 7530
rect 14382 7586 14476 7598
rect 14382 7534 14384 7586
rect 14436 7534 14476 7586
rect 14382 7532 14476 7534
rect 14382 7522 14438 7532
rect 13636 7466 13692 7478
rect 14140 7476 14196 7486
rect 13916 7474 14196 7476
rect 13916 7422 14142 7474
rect 14194 7422 14196 7474
rect 13916 7420 14196 7422
rect 13916 6802 13972 7420
rect 14140 7410 14196 7420
rect 15820 7474 15876 7756
rect 16156 7700 16212 7710
rect 16156 7606 16212 7644
rect 17612 7700 17668 8206
rect 18396 8258 18452 8372
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 18396 7700 18452 8206
rect 19740 8260 19796 8372
rect 22092 8426 22148 8438
rect 22092 8374 22094 8426
rect 22146 8374 22148 8426
rect 19964 8260 20020 8283
rect 19740 8258 19908 8260
rect 19740 8206 19742 8258
rect 19794 8206 19908 8258
rect 19740 8204 19908 8206
rect 19740 8194 19796 8204
rect 19740 8090 19796 8102
rect 19740 8038 19742 8090
rect 19794 8038 19796 8090
rect 18684 7868 18948 7878
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18684 7802 18948 7812
rect 18396 7644 19012 7700
rect 17612 7634 17668 7644
rect 15820 7422 15822 7474
rect 15874 7422 15876 7474
rect 15820 7410 15876 7422
rect 18396 7489 18452 7501
rect 18396 7437 18398 7489
rect 18450 7437 18452 7489
rect 18284 7364 18340 7374
rect 17500 7362 18340 7364
rect 17500 7310 18286 7362
rect 18338 7310 18340 7362
rect 17500 7308 18340 7310
rect 15772 7084 16036 7094
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 15772 7018 16036 7028
rect 13916 6750 13918 6802
rect 13970 6750 13972 6802
rect 13356 6580 13412 6590
rect 13412 6524 13468 6580
rect 13356 6514 13468 6524
rect 13244 5926 13300 5964
rect 13412 5962 13468 6514
rect 12516 5898 12572 5910
rect 13412 5910 13414 5962
rect 13466 5910 13468 5962
rect 13412 5898 13468 5910
rect 13916 5906 13972 6750
rect 14700 6804 14756 6814
rect 14700 6132 14756 6748
rect 15820 6804 15876 6814
rect 15820 6710 15876 6748
rect 17500 6802 17556 7308
rect 18284 7298 18340 7308
rect 18396 7028 18452 7437
rect 18732 7476 18788 7486
rect 18732 7382 18788 7420
rect 18956 7474 19012 7644
rect 18956 7422 18958 7474
rect 19010 7422 19012 7474
rect 18396 6972 18676 7028
rect 17500 6750 17502 6802
rect 17554 6750 17556 6802
rect 17500 6738 17556 6750
rect 16604 6692 16660 6702
rect 16716 6692 16772 6702
rect 16604 6690 16772 6692
rect 16604 6638 16606 6690
rect 16658 6638 16718 6690
rect 16770 6638 16772 6690
rect 16604 6636 16772 6638
rect 16604 6626 16660 6636
rect 16716 6468 16772 6636
rect 16716 6402 16772 6412
rect 18284 6468 18340 6478
rect 18620 6468 18676 6972
rect 14812 6132 14868 6142
rect 14700 6130 14868 6132
rect 14700 6078 14814 6130
rect 14866 6078 14868 6130
rect 14700 6076 14868 6078
rect 14812 6066 14868 6076
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13916 5842 13972 5854
rect 14158 5908 14214 5918
rect 14476 5908 14532 5918
rect 14158 5906 14532 5908
rect 14158 5854 14160 5906
rect 14212 5854 14478 5906
rect 14530 5854 14532 5906
rect 14158 5852 14532 5854
rect 14158 5842 14214 5852
rect 14476 5842 14532 5852
rect 15772 5516 16036 5526
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 15772 5450 16036 5460
rect 12460 5236 12516 5246
rect 12012 5234 12516 5236
rect 12012 5182 12462 5234
rect 12514 5182 12516 5234
rect 12012 5180 12516 5182
rect 12460 5170 12516 5180
rect 9772 5070 9774 5122
rect 9826 5070 9828 5122
rect 9772 5058 9828 5070
rect 18284 5124 18340 6412
rect 18508 6412 18676 6468
rect 18956 6468 19012 7422
rect 19740 7474 19796 8038
rect 19740 7422 19742 7474
rect 19794 7422 19796 7474
rect 19740 7410 19796 7422
rect 19852 7476 19908 8204
rect 19964 8191 19966 8204
rect 20018 8191 20020 8204
rect 22092 8260 22148 8374
rect 22092 8194 22148 8204
rect 22204 8260 22260 8270
rect 22204 8258 22372 8260
rect 22204 8206 22206 8258
rect 22258 8206 22372 8258
rect 22204 8204 22372 8206
rect 22204 8194 22260 8204
rect 19964 8179 20020 8191
rect 21644 7700 21700 7710
rect 21644 7588 21700 7644
rect 19852 6692 19908 7420
rect 21420 7586 21700 7588
rect 21420 7534 21646 7586
rect 21698 7534 21700 7586
rect 21420 7532 21700 7534
rect 21420 6916 21476 7532
rect 21644 7522 21700 7532
rect 21980 7588 22036 7598
rect 21596 7084 21860 7094
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21596 7018 21860 7028
rect 21420 6860 21700 6916
rect 19964 6692 20020 6702
rect 20524 6692 20580 6702
rect 19852 6690 20132 6692
rect 19852 6638 19966 6690
rect 20018 6638 20132 6690
rect 20412 6690 20580 6692
rect 19852 6636 20132 6638
rect 19964 6626 20020 6636
rect 19404 6580 19460 6590
rect 19404 6578 19684 6580
rect 19404 6526 19406 6578
rect 19458 6526 19684 6578
rect 19404 6524 19684 6526
rect 19404 6514 19460 6524
rect 18508 6018 18564 6412
rect 18956 6402 19012 6412
rect 18684 6300 18948 6310
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18684 6234 18948 6244
rect 18508 5966 18510 6018
rect 18562 5966 18564 6018
rect 18508 5954 18564 5966
rect 18751 6132 18807 6142
rect 18751 5962 18807 6076
rect 18751 5910 18753 5962
rect 18805 5910 18807 5962
rect 18751 5898 18807 5910
rect 19628 6020 19684 6524
rect 19964 6522 20020 6534
rect 19964 6470 19966 6522
rect 20018 6470 20020 6522
rect 19964 6020 20020 6470
rect 19628 5906 19684 5964
rect 19628 5854 19630 5906
rect 19682 5854 19684 5906
rect 19628 5842 19684 5854
rect 19852 5964 20020 6020
rect 19740 5124 19796 5134
rect 19852 5124 19908 5964
rect 20076 5950 20132 6636
rect 20300 6634 20356 6646
rect 20300 6582 20302 6634
rect 20354 6582 20356 6634
rect 20300 6132 20356 6582
rect 20300 6066 20356 6076
rect 20412 6638 20526 6690
rect 20578 6638 20580 6690
rect 20412 6636 20580 6638
rect 20076 5898 20078 5950
rect 20130 5898 20132 5950
rect 20300 5908 20356 5918
rect 20076 5886 20132 5898
rect 20188 5906 20356 5908
rect 20188 5854 20302 5906
rect 20354 5854 20356 5906
rect 20188 5852 20356 5854
rect 19740 5122 19908 5124
rect 7036 4732 7300 4742
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7036 4666 7300 4676
rect 12860 4732 13124 4742
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 12860 4666 13124 4676
rect 18284 4338 18340 5068
rect 19068 5053 19572 5109
rect 19740 5070 19742 5122
rect 19794 5070 19908 5122
rect 19740 5068 19908 5070
rect 19964 5794 20020 5806
rect 19964 5742 19966 5794
rect 20018 5742 20020 5794
rect 19740 5058 19796 5068
rect 18684 4732 18948 4742
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18684 4666 18948 4676
rect 18284 4286 18286 4338
rect 18338 4286 18340 4338
rect 18284 4274 18340 4286
rect 19068 4338 19124 5053
rect 19404 4898 19460 4910
rect 19404 4846 19406 4898
rect 19458 4846 19460 4898
rect 19404 4564 19460 4846
rect 19516 4900 19572 5053
rect 19964 4900 20020 5742
rect 20188 5796 20244 5852
rect 20300 5842 20356 5852
rect 20076 5124 20132 5134
rect 20188 5124 20244 5740
rect 20076 5122 20244 5124
rect 20076 5070 20078 5122
rect 20130 5070 20244 5122
rect 20076 5068 20244 5070
rect 20300 5684 20356 5694
rect 20300 5107 20356 5628
rect 20412 5234 20468 6636
rect 20524 6626 20580 6636
rect 21644 6690 21700 6860
rect 21644 6638 21646 6690
rect 21698 6638 21700 6690
rect 21644 6626 21700 6638
rect 21812 6634 21868 6646
rect 21812 6582 21814 6634
rect 21866 6582 21868 6634
rect 21812 6524 21868 6582
rect 21756 6468 21868 6524
rect 21980 6578 22036 7532
rect 22204 7474 22260 7486
rect 22204 7422 22206 7474
rect 22258 7422 22260 7474
rect 21980 6526 21982 6578
rect 22034 6526 22036 6578
rect 21980 6468 22036 6526
rect 20804 6132 20860 6142
rect 20804 6018 20860 6076
rect 20804 5966 20806 6018
rect 20858 5966 20860 6018
rect 20804 5954 20860 5966
rect 20412 5182 20414 5234
rect 20466 5182 20468 5234
rect 20412 5170 20468 5182
rect 20972 5908 21028 5918
rect 20972 5236 21028 5852
rect 21084 5906 21140 5918
rect 21084 5854 21086 5906
rect 21138 5854 21140 5906
rect 21084 5684 21140 5854
rect 21196 5906 21252 5918
rect 21196 5854 21198 5906
rect 21250 5854 21252 5906
rect 21196 5796 21252 5854
rect 21420 5908 21476 5918
rect 21420 5814 21476 5852
rect 21196 5730 21252 5740
rect 21756 5796 21812 6468
rect 21756 5702 21812 5740
rect 21084 5618 21140 5628
rect 21980 5684 22036 6412
rect 22092 6690 22148 6702
rect 22092 6638 22094 6690
rect 22146 6638 22148 6690
rect 22092 6020 22148 6638
rect 22092 5954 22148 5964
rect 22204 5908 22260 7422
rect 22316 6926 22372 8204
rect 22540 8258 22596 9548
rect 23343 9098 23399 9548
rect 23548 9604 23604 10558
rect 23772 10610 23828 10622
rect 23772 10558 23774 10610
rect 23826 10558 23828 10610
rect 23772 10164 23828 10558
rect 24108 10388 24164 10398
rect 24108 10386 24276 10388
rect 24108 10334 24110 10386
rect 24162 10334 24276 10386
rect 24108 10332 24276 10334
rect 24108 10322 24164 10332
rect 23772 10098 23828 10108
rect 23548 9538 23604 9548
rect 23884 9714 23940 9726
rect 23884 9662 23886 9714
rect 23938 9662 23940 9714
rect 23884 9604 23940 9662
rect 23884 9538 23940 9548
rect 23343 9046 23345 9098
rect 23397 9046 23399 9098
rect 23343 9034 23399 9046
rect 24220 9042 24276 10332
rect 24508 9436 24772 9446
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24508 9370 24772 9380
rect 24220 8990 24222 9042
rect 24274 8990 24276 9042
rect 24220 8978 24276 8990
rect 22708 8930 22764 8942
rect 22708 8878 22710 8930
rect 22762 8878 22764 8930
rect 22708 8428 22764 8878
rect 23100 8820 23156 8830
rect 23100 8818 23268 8820
rect 23100 8766 23102 8818
rect 23154 8766 23268 8818
rect 23100 8764 23268 8766
rect 23100 8754 23156 8764
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22428 7588 22484 7598
rect 22428 7530 22484 7532
rect 22428 7478 22430 7530
rect 22482 7478 22484 7530
rect 22428 7466 22484 7478
rect 22428 7364 22484 7374
rect 22540 7364 22596 8206
rect 22428 7362 22596 7364
rect 22428 7310 22430 7362
rect 22482 7310 22596 7362
rect 22428 7308 22596 7310
rect 22652 8372 22764 8428
rect 23100 8372 23156 8382
rect 22428 7298 22484 7308
rect 22316 6914 22428 6926
rect 22316 6862 22374 6914
rect 22426 6862 22428 6914
rect 22316 6860 22428 6862
rect 22372 6850 22428 6860
rect 22652 6244 22708 8372
rect 23100 8278 23156 8316
rect 23100 7700 23156 7710
rect 22652 6178 22708 6188
rect 22764 7474 22820 7486
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22559 6020 22615 6030
rect 22764 6020 22820 7422
rect 23100 7474 23156 7644
rect 23100 7422 23102 7474
rect 23154 7422 23156 7474
rect 23100 7410 23156 7422
rect 23212 6916 23268 8764
rect 24892 8372 24948 14924
rect 24892 8306 24948 8316
rect 24220 8258 24276 8270
rect 23343 8202 23399 8214
rect 23343 8150 23345 8202
rect 23397 8150 23399 8202
rect 23343 7700 23399 8150
rect 24220 8206 24222 8258
rect 24274 8206 24276 8258
rect 23343 7634 23399 7644
rect 23772 7700 23828 7710
rect 23772 7476 23828 7644
rect 24108 7700 24164 7710
rect 24220 7700 24276 8206
rect 24508 7868 24772 7878
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24508 7802 24772 7812
rect 24108 7698 24276 7700
rect 24108 7646 24110 7698
rect 24162 7646 24276 7698
rect 24108 7644 24276 7646
rect 24108 7634 24164 7644
rect 23212 6850 23268 6860
rect 23604 7474 23828 7476
rect 23604 7422 23774 7474
rect 23826 7422 23828 7474
rect 23604 7420 23828 7422
rect 23604 6802 23660 7420
rect 23772 7410 23828 7420
rect 23604 6750 23606 6802
rect 23658 6750 23660 6802
rect 23604 6738 23660 6750
rect 23884 6916 23940 6926
rect 23212 6692 23268 6702
rect 23212 6690 23492 6692
rect 23212 6638 23214 6690
rect 23266 6638 23492 6690
rect 23212 6636 23492 6638
rect 23212 6626 23268 6636
rect 22876 6468 22932 6478
rect 22876 6374 22932 6412
rect 23436 6132 23492 6636
rect 23436 6076 23828 6132
rect 22615 5964 22820 6020
rect 22559 5962 22615 5964
rect 22559 5910 22561 5962
rect 22613 5910 22615 5962
rect 22559 5898 22615 5910
rect 23436 5908 23492 5946
rect 22204 5842 22260 5852
rect 23436 5842 23492 5852
rect 21980 5618 22036 5628
rect 22316 5684 22372 5694
rect 22316 5682 22820 5684
rect 22316 5630 22318 5682
rect 22370 5630 22820 5682
rect 22316 5628 22820 5630
rect 22316 5618 22372 5628
rect 21596 5516 21860 5526
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21596 5450 21860 5460
rect 20076 5058 20132 5068
rect 20300 5055 20302 5107
rect 20354 5055 20356 5107
rect 20300 5043 20356 5055
rect 19516 4844 20020 4900
rect 19404 4498 19460 4508
rect 20972 4450 21028 5180
rect 22428 5348 22484 5358
rect 22764 5348 22820 5628
rect 22764 5292 23044 5348
rect 20972 4398 20974 4450
rect 21026 4398 21028 4450
rect 20972 4386 21028 4398
rect 21308 5124 21364 5134
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 21308 4338 21364 5068
rect 21420 5124 21476 5134
rect 21532 5124 21588 5134
rect 21420 5122 21532 5124
rect 21420 5070 21422 5122
rect 21474 5070 21532 5122
rect 21420 5068 21532 5070
rect 21420 5058 21476 5068
rect 21532 5058 21588 5068
rect 22296 5066 22352 5078
rect 22296 5014 22298 5066
rect 22350 5014 22352 5066
rect 22296 4676 22352 5014
rect 22204 4620 22352 4676
rect 21308 4286 21310 4338
rect 21362 4286 21364 4338
rect 21308 4274 21364 4286
rect 22092 4340 22148 4350
rect 22092 4246 22148 4284
rect 22204 4116 22260 4620
rect 22428 4564 22484 5292
rect 22540 5124 22596 5134
rect 22540 5030 22596 5068
rect 22988 5122 23044 5292
rect 23324 5236 23380 5246
rect 23324 5142 23380 5180
rect 22988 5070 22990 5122
rect 23042 5070 23044 5122
rect 23660 5124 23716 5134
rect 22988 5058 23044 5070
rect 23436 5066 23492 5078
rect 22372 4508 22484 4564
rect 23436 5014 23438 5066
rect 23490 5014 23492 5066
rect 23660 5030 23716 5068
rect 22372 4452 22428 4508
rect 21980 4060 22260 4116
rect 22316 4396 22428 4452
rect 4124 3948 4388 3958
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4124 3882 4388 3892
rect 9948 3948 10212 3958
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 9948 3882 10212 3892
rect 15772 3948 16036 3958
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 15772 3882 16036 3892
rect 21596 3948 21860 3958
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21596 3882 21860 3892
rect 21868 3780 21924 3790
rect 21980 3780 22036 4060
rect 22316 3892 22372 4396
rect 21868 3778 22036 3780
rect 21868 3726 21870 3778
rect 21922 3726 22036 3778
rect 21868 3724 22036 3726
rect 22092 3836 22372 3892
rect 23192 4004 23248 4014
rect 21868 3714 21924 3724
rect 21532 3554 21588 3566
rect 21532 3502 21534 3554
rect 21586 3502 21588 3554
rect 21364 3444 21420 3454
rect 21532 3444 21588 3502
rect 22092 3556 22148 3836
rect 22316 3556 22372 3566
rect 22092 3554 22372 3556
rect 22092 3502 22318 3554
rect 22370 3502 22372 3554
rect 22092 3500 22372 3502
rect 22316 3490 22372 3500
rect 23192 3554 23248 3948
rect 23436 3778 23492 5014
rect 23772 4788 23828 6076
rect 23884 5124 23940 6860
rect 24332 6692 24388 6702
rect 24220 6690 24388 6692
rect 24220 6638 24334 6690
rect 24386 6638 24388 6690
rect 24220 6636 24388 6638
rect 23996 6466 24052 6478
rect 23996 6414 23998 6466
rect 24050 6414 24052 6466
rect 23996 5908 24052 6414
rect 23996 5842 24052 5852
rect 24220 5908 24276 6636
rect 24332 6626 24388 6636
rect 24508 6300 24772 6310
rect 23996 5682 24052 5694
rect 23996 5630 23998 5682
rect 24050 5630 24052 5682
rect 23996 5348 24052 5630
rect 23996 5282 24052 5292
rect 23996 5124 24052 5134
rect 23884 5122 24052 5124
rect 23884 5070 23998 5122
rect 24050 5070 24052 5122
rect 23884 5068 24052 5070
rect 23996 5058 24052 5068
rect 23772 4732 24052 4788
rect 23996 4450 24052 4732
rect 23996 4398 23998 4450
rect 24050 4398 24052 4450
rect 23996 4004 24052 4398
rect 23996 3938 24052 3948
rect 23436 3726 23438 3778
rect 23490 3726 23492 3778
rect 23436 3714 23492 3726
rect 24052 3668 24108 3678
rect 24220 3668 24276 5852
rect 24332 6244 24388 6254
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24508 6234 24772 6244
rect 24332 5906 24388 6188
rect 24332 5854 24334 5906
rect 24386 5854 24388 5906
rect 24332 3892 24388 5854
rect 25004 5236 25060 16828
rect 25004 5170 25060 5180
rect 24508 4732 24772 4742
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24508 4666 24772 4676
rect 24332 3826 24388 3836
rect 24052 3666 24276 3668
rect 24052 3614 24054 3666
rect 24106 3614 24276 3666
rect 24052 3612 24276 3614
rect 24052 3602 24108 3612
rect 23192 3502 23194 3554
rect 23246 3502 23248 3554
rect 23192 3490 23248 3502
rect 21364 3442 21588 3444
rect 21364 3390 21366 3442
rect 21418 3390 21588 3442
rect 21364 3388 21588 3390
rect 21364 3378 21420 3388
rect 7036 3164 7300 3174
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7036 3098 7300 3108
rect 12860 3164 13124 3174
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 12860 3098 13124 3108
rect 18684 3164 18948 3174
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18684 3098 18948 3108
rect 21532 1876 21588 3388
rect 24508 3164 24772 3174
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24508 3098 24772 3108
rect 21532 1810 21588 1820
<< via2 >>
rect 4124 22762 4180 22764
rect 4124 22710 4126 22762
rect 4126 22710 4178 22762
rect 4178 22710 4180 22762
rect 4124 22708 4180 22710
rect 4228 22762 4284 22764
rect 4228 22710 4230 22762
rect 4230 22710 4282 22762
rect 4282 22710 4284 22762
rect 4228 22708 4284 22710
rect 4332 22762 4388 22764
rect 4332 22710 4334 22762
rect 4334 22710 4386 22762
rect 4386 22710 4388 22762
rect 4332 22708 4388 22710
rect 4124 21194 4180 21196
rect 4124 21142 4126 21194
rect 4126 21142 4178 21194
rect 4178 21142 4180 21194
rect 4124 21140 4180 21142
rect 4228 21194 4284 21196
rect 4228 21142 4230 21194
rect 4230 21142 4282 21194
rect 4282 21142 4284 21194
rect 4228 21140 4284 21142
rect 4332 21194 4388 21196
rect 4332 21142 4334 21194
rect 4334 21142 4386 21194
rect 4386 21142 4388 21194
rect 4332 21140 4388 21142
rect 4124 19626 4180 19628
rect 4124 19574 4126 19626
rect 4126 19574 4178 19626
rect 4178 19574 4180 19626
rect 4124 19572 4180 19574
rect 4228 19626 4284 19628
rect 4228 19574 4230 19626
rect 4230 19574 4282 19626
rect 4282 19574 4284 19626
rect 4228 19572 4284 19574
rect 4332 19626 4388 19628
rect 4332 19574 4334 19626
rect 4334 19574 4386 19626
rect 4386 19574 4388 19626
rect 4332 19572 4388 19574
rect 2828 18620 2884 18676
rect 4284 18450 4340 18452
rect 4284 18398 4286 18450
rect 4286 18398 4338 18450
rect 4338 18398 4340 18450
rect 4284 18396 4340 18398
rect 4124 18058 4180 18060
rect 4124 18006 4126 18058
rect 4126 18006 4178 18058
rect 4178 18006 4180 18058
rect 4124 18004 4180 18006
rect 4228 18058 4284 18060
rect 4228 18006 4230 18058
rect 4230 18006 4282 18058
rect 4282 18006 4284 18058
rect 4228 18004 4284 18006
rect 4332 18058 4388 18060
rect 4332 18006 4334 18058
rect 4334 18006 4386 18058
rect 4386 18006 4388 18058
rect 4332 18004 4388 18006
rect 3276 16940 3332 16996
rect 3724 17052 3780 17108
rect 2380 16828 2436 16884
rect 3388 16828 3444 16884
rect 2828 16098 2884 16100
rect 2828 16046 2830 16098
rect 2830 16046 2882 16098
rect 2882 16046 2884 16098
rect 2828 16044 2884 16046
rect 3052 16156 3108 16212
rect 3164 15708 3220 15764
rect 4172 17666 4228 17668
rect 4172 17614 4174 17666
rect 4174 17614 4226 17666
rect 4226 17614 4228 17666
rect 4172 17612 4228 17614
rect 4060 16940 4116 16996
rect 4284 17276 4340 17332
rect 4396 16940 4452 16996
rect 3612 16716 3668 16772
rect 3612 16156 3668 16212
rect 3500 16098 3556 16100
rect 3500 16046 3502 16098
rect 3502 16046 3554 16098
rect 3554 16046 3556 16098
rect 3500 16044 3556 16046
rect 3500 14252 3556 14308
rect 2828 13746 2884 13748
rect 2828 13694 2830 13746
rect 2830 13694 2882 13746
rect 2882 13694 2884 13746
rect 2828 13692 2884 13694
rect 1596 13468 1652 13524
rect 7196 22092 7252 22148
rect 7036 21978 7092 21980
rect 7036 21926 7038 21978
rect 7038 21926 7090 21978
rect 7090 21926 7092 21978
rect 7036 21924 7092 21926
rect 7140 21978 7196 21980
rect 7140 21926 7142 21978
rect 7142 21926 7194 21978
rect 7194 21926 7196 21978
rect 7140 21924 7196 21926
rect 7244 21978 7300 21980
rect 7244 21926 7246 21978
rect 7246 21926 7298 21978
rect 7298 21926 7300 21978
rect 7244 21924 7300 21926
rect 9948 22762 10004 22764
rect 9948 22710 9950 22762
rect 9950 22710 10002 22762
rect 10002 22710 10004 22762
rect 9948 22708 10004 22710
rect 10052 22762 10108 22764
rect 10052 22710 10054 22762
rect 10054 22710 10106 22762
rect 10106 22710 10108 22762
rect 10052 22708 10108 22710
rect 10156 22762 10212 22764
rect 10156 22710 10158 22762
rect 10158 22710 10210 22762
rect 10210 22710 10212 22762
rect 10156 22708 10212 22710
rect 7420 21532 7476 21588
rect 5516 21474 5572 21476
rect 5516 21422 5518 21474
rect 5518 21422 5570 21474
rect 5570 21422 5572 21474
rect 5516 21420 5572 21422
rect 7980 21474 8036 21476
rect 7980 21422 7982 21474
rect 7982 21422 8034 21474
rect 8034 21422 8036 21474
rect 7980 21420 8036 21422
rect 10108 22316 10164 22372
rect 8428 22092 8484 22148
rect 8204 21586 8260 21588
rect 8204 21534 8206 21586
rect 8206 21534 8258 21586
rect 8258 21534 8260 21586
rect 8204 21532 8260 21534
rect 7980 20860 8036 20916
rect 4676 20242 4732 20244
rect 4676 20190 4678 20242
rect 4678 20190 4730 20242
rect 4730 20190 4732 20242
rect 4676 20188 4732 20190
rect 5516 20188 5572 20244
rect 7036 20410 7092 20412
rect 7036 20358 7038 20410
rect 7038 20358 7090 20410
rect 7090 20358 7092 20410
rect 7036 20356 7092 20358
rect 7140 20410 7196 20412
rect 7140 20358 7142 20410
rect 7142 20358 7194 20410
rect 7194 20358 7196 20410
rect 7140 20356 7196 20358
rect 7244 20410 7300 20412
rect 7244 20358 7246 20410
rect 7246 20358 7298 20410
rect 7298 20358 7300 20410
rect 7244 20356 7300 20358
rect 6300 20188 6356 20244
rect 4732 18844 4788 18900
rect 4676 17666 4732 17668
rect 4676 17614 4678 17666
rect 4678 17614 4730 17666
rect 4730 17614 4732 17666
rect 4676 17612 4732 17614
rect 4620 17052 4676 17108
rect 6188 19852 6244 19908
rect 5068 18844 5124 18900
rect 5068 18284 5124 18340
rect 9324 22092 9380 22148
rect 8092 20748 8148 20804
rect 9212 20802 9268 20804
rect 9212 20750 9214 20802
rect 9214 20750 9266 20802
rect 9266 20750 9268 20802
rect 9212 20748 9268 20750
rect 8764 20188 8820 20244
rect 8988 20524 9044 20580
rect 7036 18842 7092 18844
rect 7036 18790 7038 18842
rect 7038 18790 7090 18842
rect 7090 18790 7092 18842
rect 7036 18788 7092 18790
rect 7140 18842 7196 18844
rect 7140 18790 7142 18842
rect 7142 18790 7194 18842
rect 7194 18790 7196 18842
rect 7140 18788 7196 18790
rect 7244 18842 7300 18844
rect 7244 18790 7246 18842
rect 7246 18790 7298 18842
rect 7298 18790 7300 18842
rect 7244 18788 7300 18790
rect 5292 18450 5348 18452
rect 5292 18398 5294 18450
rect 5294 18398 5346 18450
rect 5346 18398 5348 18450
rect 5292 18396 5348 18398
rect 6728 18284 6784 18340
rect 4956 17500 5012 17556
rect 5068 17052 5124 17108
rect 4956 16828 5012 16884
rect 4124 16490 4180 16492
rect 4124 16438 4126 16490
rect 4126 16438 4178 16490
rect 4178 16438 4180 16490
rect 4124 16436 4180 16438
rect 4228 16490 4284 16492
rect 4228 16438 4230 16490
rect 4230 16438 4282 16490
rect 4282 16438 4284 16490
rect 4228 16436 4284 16438
rect 4332 16490 4388 16492
rect 4332 16438 4334 16490
rect 4334 16438 4386 16490
rect 4386 16438 4388 16490
rect 4332 16436 4388 16438
rect 3836 15708 3892 15764
rect 4396 16156 4452 16212
rect 4562 16044 4618 16100
rect 4284 15820 4340 15876
rect 3948 15372 4004 15428
rect 4508 15372 4564 15428
rect 3724 13020 3780 13076
rect 2380 12962 2436 12964
rect 2380 12910 2382 12962
rect 2382 12910 2434 12962
rect 2434 12910 2436 12962
rect 2380 12908 2436 12910
rect 3836 12908 3892 12964
rect 4124 14922 4180 14924
rect 4124 14870 4126 14922
rect 4126 14870 4178 14922
rect 4178 14870 4180 14922
rect 4124 14868 4180 14870
rect 4228 14922 4284 14924
rect 4228 14870 4230 14922
rect 4230 14870 4282 14922
rect 4282 14870 4284 14922
rect 4228 14868 4284 14870
rect 4332 14922 4388 14924
rect 4332 14870 4334 14922
rect 4334 14870 4386 14922
rect 4386 14870 4388 14922
rect 4332 14868 4388 14870
rect 4508 13746 4564 13748
rect 4508 13694 4510 13746
rect 4510 13694 4562 13746
rect 4562 13694 4564 13746
rect 4508 13692 4564 13694
rect 4124 13354 4180 13356
rect 4124 13302 4126 13354
rect 4126 13302 4178 13354
rect 4178 13302 4180 13354
rect 4124 13300 4180 13302
rect 4228 13354 4284 13356
rect 4228 13302 4230 13354
rect 4230 13302 4282 13354
rect 4282 13302 4284 13354
rect 4228 13300 4284 13302
rect 4332 13354 4388 13356
rect 4332 13302 4334 13354
rect 4334 13302 4386 13354
rect 4386 13302 4388 13354
rect 4332 13300 4388 13302
rect 4284 13074 4340 13076
rect 4284 13022 4286 13074
rect 4286 13022 4338 13074
rect 4338 13022 4340 13074
rect 4284 13020 4340 13022
rect 4284 12684 4340 12740
rect 3276 12236 3332 12292
rect 3836 12236 3892 12292
rect 4172 12178 4228 12180
rect 4172 12126 4174 12178
rect 4174 12126 4226 12178
rect 4226 12126 4228 12178
rect 4172 12124 4228 12126
rect 4124 11786 4180 11788
rect 4124 11734 4126 11786
rect 4126 11734 4178 11786
rect 4178 11734 4180 11786
rect 4124 11732 4180 11734
rect 4228 11786 4284 11788
rect 4228 11734 4230 11786
rect 4230 11734 4282 11786
rect 4282 11734 4284 11786
rect 4228 11732 4284 11734
rect 4332 11786 4388 11788
rect 4332 11734 4334 11786
rect 4334 11734 4386 11786
rect 4386 11734 4388 11786
rect 4332 11732 4388 11734
rect 4732 15036 4788 15092
rect 5628 15932 5684 15988
rect 6524 17948 6580 18004
rect 6300 17666 6356 17668
rect 6300 17614 6302 17666
rect 6302 17614 6354 17666
rect 6354 17614 6356 17666
rect 6300 17612 6356 17614
rect 6020 17388 6076 17444
rect 5852 17164 5908 17220
rect 6412 17388 6468 17444
rect 6412 17164 6468 17220
rect 6300 16940 6356 16996
rect 7532 17836 7588 17892
rect 7868 17836 7924 17892
rect 8092 18172 8148 18228
rect 7036 17274 7092 17276
rect 7036 17222 7038 17274
rect 7038 17222 7090 17274
rect 7090 17222 7092 17274
rect 7036 17220 7092 17222
rect 7140 17274 7196 17276
rect 7140 17222 7142 17274
rect 7142 17222 7194 17274
rect 7194 17222 7196 17274
rect 7140 17220 7196 17222
rect 7244 17274 7300 17276
rect 7244 17222 7246 17274
rect 7246 17222 7298 17274
rect 7298 17222 7300 17274
rect 7244 17220 7300 17222
rect 6860 16882 6916 16884
rect 6860 16830 6862 16882
rect 6862 16830 6914 16882
rect 6914 16830 6916 16882
rect 6860 16828 6916 16830
rect 9212 19964 9268 20020
rect 8988 19122 9044 19124
rect 8988 19070 8990 19122
rect 8990 19070 9042 19122
rect 9042 19070 9044 19122
rect 8988 19068 9044 19070
rect 9212 19068 9268 19124
rect 11564 22370 11620 22372
rect 11564 22318 11566 22370
rect 11566 22318 11618 22370
rect 11618 22318 11620 22370
rect 11564 22316 11620 22318
rect 15772 22762 15828 22764
rect 15772 22710 15774 22762
rect 15774 22710 15826 22762
rect 15826 22710 15828 22762
rect 15772 22708 15828 22710
rect 15876 22762 15932 22764
rect 15876 22710 15878 22762
rect 15878 22710 15930 22762
rect 15930 22710 15932 22762
rect 15876 22708 15932 22710
rect 15980 22762 16036 22764
rect 15980 22710 15982 22762
rect 15982 22710 16034 22762
rect 16034 22710 16036 22762
rect 15980 22708 16036 22710
rect 22876 23996 22932 24052
rect 21596 22762 21652 22764
rect 21596 22710 21598 22762
rect 21598 22710 21650 22762
rect 21650 22710 21652 22762
rect 21596 22708 21652 22710
rect 21700 22762 21756 22764
rect 21700 22710 21702 22762
rect 21702 22710 21754 22762
rect 21754 22710 21756 22762
rect 21700 22708 21756 22710
rect 21804 22762 21860 22764
rect 21804 22710 21806 22762
rect 21806 22710 21858 22762
rect 21858 22710 21860 22762
rect 21804 22708 21860 22710
rect 21308 22540 21364 22596
rect 22540 22594 22596 22596
rect 22540 22542 22542 22594
rect 22542 22542 22594 22594
rect 22594 22542 22596 22594
rect 22540 22540 22596 22542
rect 12796 22316 12852 22372
rect 13580 22370 13636 22372
rect 13580 22318 13582 22370
rect 13582 22318 13634 22370
rect 13634 22318 13636 22370
rect 13580 22316 13636 22318
rect 13972 22370 14028 22372
rect 13972 22318 13974 22370
rect 13974 22318 14026 22370
rect 14026 22318 14028 22370
rect 13972 22316 14028 22318
rect 19572 22258 19628 22260
rect 19572 22206 19574 22258
rect 19574 22206 19626 22258
rect 19626 22206 19628 22258
rect 19572 22204 19628 22206
rect 19740 22204 19796 22260
rect 9948 21194 10004 21196
rect 9948 21142 9950 21194
rect 9950 21142 10002 21194
rect 10002 21142 10004 21194
rect 9948 21140 10004 21142
rect 10052 21194 10108 21196
rect 10052 21142 10054 21194
rect 10054 21142 10106 21194
rect 10106 21142 10108 21194
rect 10052 21140 10108 21142
rect 10156 21194 10212 21196
rect 10156 21142 10158 21194
rect 10158 21142 10210 21194
rect 10210 21142 10212 21194
rect 10156 21140 10212 21142
rect 10332 21084 10388 21140
rect 10332 20860 10388 20916
rect 9660 20763 9716 20804
rect 9660 20748 9662 20763
rect 9662 20748 9714 20763
rect 9714 20748 9716 20763
rect 11340 21474 11396 21476
rect 11340 21422 11342 21474
rect 11342 21422 11394 21474
rect 11394 21422 11396 21474
rect 11340 21420 11396 21422
rect 10892 20860 10948 20916
rect 11340 21084 11396 21140
rect 10556 20802 10612 20804
rect 10556 20750 10558 20802
rect 10558 20750 10610 20802
rect 10610 20750 10612 20802
rect 10556 20748 10612 20750
rect 10444 20524 10500 20580
rect 11676 20802 11732 20804
rect 11676 20750 11678 20802
rect 11678 20750 11730 20802
rect 11730 20750 11732 20802
rect 11676 20748 11732 20750
rect 12124 20748 12180 20804
rect 12236 20860 12292 20916
rect 11564 20188 11620 20244
rect 9660 20018 9716 20020
rect 9660 19966 9662 20018
rect 9662 19966 9714 20018
rect 9714 19966 9716 20018
rect 9660 19964 9716 19966
rect 9884 20076 9940 20132
rect 10668 20018 10724 20020
rect 10668 19966 10670 20018
rect 10670 19966 10722 20018
rect 10722 19966 10724 20018
rect 10668 19964 10724 19966
rect 11732 19906 11788 19908
rect 11732 19854 11734 19906
rect 11734 19854 11786 19906
rect 11786 19854 11788 19906
rect 11732 19852 11788 19854
rect 9492 19180 9548 19236
rect 9948 19626 10004 19628
rect 9948 19574 9950 19626
rect 9950 19574 10002 19626
rect 10002 19574 10004 19626
rect 9948 19572 10004 19574
rect 10052 19626 10108 19628
rect 10052 19574 10054 19626
rect 10054 19574 10106 19626
rect 10106 19574 10108 19626
rect 10052 19572 10108 19574
rect 10156 19626 10212 19628
rect 10156 19574 10158 19626
rect 10158 19574 10210 19626
rect 10210 19574 10212 19626
rect 10156 19572 10212 19574
rect 12348 19964 12404 20020
rect 9660 19292 9716 19348
rect 10220 19234 10276 19236
rect 10220 19182 10222 19234
rect 10222 19182 10274 19234
rect 10274 19182 10276 19234
rect 10220 19180 10276 19182
rect 9996 18508 10052 18564
rect 8652 17836 8708 17892
rect 8092 17276 8148 17332
rect 8316 17666 8372 17668
rect 8316 17614 8318 17666
rect 8318 17614 8370 17666
rect 8370 17614 8372 17666
rect 8316 17612 8372 17614
rect 8484 17666 8540 17668
rect 8484 17614 8486 17666
rect 8486 17614 8538 17666
rect 8538 17614 8540 17666
rect 8484 17612 8540 17614
rect 9948 18058 10004 18060
rect 9948 18006 9950 18058
rect 9950 18006 10002 18058
rect 10002 18006 10004 18058
rect 9948 18004 10004 18006
rect 10052 18058 10108 18060
rect 10052 18006 10054 18058
rect 10054 18006 10106 18058
rect 10106 18006 10108 18058
rect 10052 18004 10108 18006
rect 10156 18058 10212 18060
rect 10156 18006 10158 18058
rect 10158 18006 10210 18058
rect 10210 18006 10212 18058
rect 10156 18004 10212 18006
rect 10556 17724 10612 17780
rect 8316 17164 8372 17220
rect 8540 17388 8596 17444
rect 5740 15372 5796 15428
rect 6636 15932 6692 15988
rect 6300 15820 6356 15876
rect 7868 16828 7924 16884
rect 7644 16604 7700 16660
rect 7644 15932 7700 15988
rect 7036 15706 7092 15708
rect 7036 15654 7038 15706
rect 7038 15654 7090 15706
rect 7090 15654 7092 15706
rect 7036 15652 7092 15654
rect 7140 15706 7196 15708
rect 7140 15654 7142 15706
rect 7142 15654 7194 15706
rect 7194 15654 7196 15706
rect 7140 15652 7196 15654
rect 7244 15706 7300 15708
rect 7244 15654 7246 15706
rect 7246 15654 7298 15706
rect 7298 15654 7300 15706
rect 7244 15652 7300 15654
rect 7420 15314 7476 15316
rect 7420 15262 7422 15314
rect 7422 15262 7474 15314
rect 7474 15262 7476 15314
rect 7420 15260 7476 15262
rect 7532 15372 7588 15428
rect 7254 15148 7310 15204
rect 6412 15036 6468 15092
rect 4900 14306 4956 14308
rect 4900 14254 4902 14306
rect 4902 14254 4954 14306
rect 4954 14254 4956 14306
rect 4900 14252 4956 14254
rect 4844 13804 4900 13860
rect 4620 13580 4676 13636
rect 4900 13468 4956 13524
rect 5796 14530 5852 14532
rect 5796 14478 5798 14530
rect 5798 14478 5850 14530
rect 5850 14478 5852 14530
rect 5796 14476 5852 14478
rect 6076 13356 6132 13412
rect 5068 12908 5124 12964
rect 5180 12348 5236 12404
rect 4732 12236 4788 12292
rect 3948 11452 4004 11508
rect 4620 11228 4676 11284
rect 5068 12236 5124 12292
rect 4956 12124 5012 12180
rect 5740 12962 5796 12964
rect 5740 12910 5742 12962
rect 5742 12910 5794 12962
rect 5794 12910 5796 12962
rect 5740 12908 5796 12910
rect 5964 12962 6020 12964
rect 5964 12910 5966 12962
rect 5966 12910 6018 12962
rect 6018 12910 6020 12962
rect 5964 12908 6020 12910
rect 5964 12684 6020 12740
rect 5404 12178 5460 12180
rect 5404 12126 5406 12178
rect 5406 12126 5458 12178
rect 5458 12126 5460 12178
rect 5404 12124 5460 12126
rect 5068 11340 5124 11396
rect 6076 11788 6132 11844
rect 6188 12236 6244 12292
rect 5796 11452 5852 11508
rect 5628 11394 5684 11396
rect 5628 11342 5630 11394
rect 5630 11342 5682 11394
rect 5682 11342 5684 11394
rect 5628 11340 5684 11342
rect 6860 15090 6916 15092
rect 6860 15038 6862 15090
rect 6862 15038 6914 15090
rect 6914 15038 6916 15090
rect 6860 15036 6916 15038
rect 7980 16098 8036 16100
rect 7980 16046 7982 16098
rect 7982 16046 8034 16098
rect 8034 16046 8036 16098
rect 7980 16044 8036 16046
rect 7980 15314 8036 15316
rect 7980 15262 7982 15314
rect 7982 15262 8034 15314
rect 8034 15262 8036 15314
rect 7980 15260 8036 15262
rect 7420 15036 7476 15092
rect 6524 14530 6580 14532
rect 6524 14478 6526 14530
rect 6526 14478 6578 14530
rect 6578 14478 6580 14530
rect 6524 14476 6580 14478
rect 7036 14138 7092 14140
rect 7036 14086 7038 14138
rect 7038 14086 7090 14138
rect 7090 14086 7092 14138
rect 7036 14084 7092 14086
rect 7140 14138 7196 14140
rect 7140 14086 7142 14138
rect 7142 14086 7194 14138
rect 7194 14086 7196 14138
rect 7140 14084 7196 14086
rect 7244 14138 7300 14140
rect 7244 14086 7246 14138
rect 7246 14086 7298 14138
rect 7298 14086 7300 14138
rect 7244 14084 7300 14086
rect 6972 13804 7028 13860
rect 6524 13692 6580 13748
rect 6524 13468 6580 13524
rect 6748 13244 6804 13300
rect 6860 13132 6916 13188
rect 7084 13020 7140 13076
rect 7532 13804 7588 13860
rect 7252 12962 7308 12964
rect 7252 12910 7254 12962
rect 7254 12910 7306 12962
rect 7306 12910 7308 12962
rect 7252 12908 7308 12910
rect 7420 13132 7476 13188
rect 7756 13692 7812 13748
rect 7868 14476 7924 14532
rect 8204 17052 8260 17108
rect 8316 16940 8372 16996
rect 8204 16882 8260 16884
rect 8204 16830 8206 16882
rect 8206 16830 8258 16882
rect 8258 16830 8260 16882
rect 8204 16828 8260 16830
rect 8652 17164 8708 17220
rect 8428 16604 8484 16660
rect 9212 17612 9268 17668
rect 8876 16940 8932 16996
rect 8988 17052 9044 17108
rect 8764 16828 8820 16884
rect 8260 14476 8316 14532
rect 9884 16940 9940 16996
rect 9548 16882 9604 16884
rect 9548 16830 9550 16882
rect 9550 16830 9602 16882
rect 9602 16830 9604 16882
rect 10220 16940 10276 16996
rect 9548 16828 9604 16830
rect 10836 19234 10892 19236
rect 10836 19182 10838 19234
rect 10838 19182 10890 19234
rect 10890 19182 10892 19234
rect 10836 19180 10892 19182
rect 11004 19122 11060 19124
rect 11004 19070 11006 19122
rect 11006 19070 11058 19122
rect 11058 19070 11060 19122
rect 11004 19068 11060 19070
rect 11116 18508 11172 18564
rect 12068 19292 12124 19348
rect 11396 19234 11452 19236
rect 11396 19182 11398 19234
rect 11398 19182 11450 19234
rect 11450 19182 11452 19234
rect 11396 19180 11452 19182
rect 11900 19234 11956 19236
rect 11900 19182 11902 19234
rect 11902 19182 11954 19234
rect 11954 19182 11956 19234
rect 11900 19180 11956 19182
rect 11116 17836 11172 17892
rect 12012 18450 12068 18452
rect 12012 18398 12014 18450
rect 12014 18398 12066 18450
rect 12066 18398 12068 18450
rect 12012 18396 12068 18398
rect 11844 17836 11900 17892
rect 12124 18172 12180 18228
rect 11564 17612 11620 17668
rect 9660 15874 9716 15876
rect 9660 15822 9662 15874
rect 9662 15822 9714 15874
rect 9714 15822 9716 15874
rect 9660 15820 9716 15822
rect 8876 15484 8932 15540
rect 9948 16490 10004 16492
rect 9948 16438 9950 16490
rect 9950 16438 10002 16490
rect 10002 16438 10004 16490
rect 9948 16436 10004 16438
rect 10052 16490 10108 16492
rect 10052 16438 10054 16490
rect 10054 16438 10106 16490
rect 10106 16438 10108 16490
rect 10052 16436 10108 16438
rect 10156 16490 10212 16492
rect 10156 16438 10158 16490
rect 10158 16438 10210 16490
rect 10210 16438 10212 16490
rect 10156 16436 10212 16438
rect 10556 15820 10612 15876
rect 10220 15484 10276 15540
rect 9772 15260 9828 15316
rect 8764 14364 8820 14420
rect 7532 12796 7588 12852
rect 7644 13468 7700 13524
rect 7644 13020 7700 13076
rect 7980 13804 8036 13860
rect 8316 13804 8372 13860
rect 8540 13522 8596 13524
rect 8540 13470 8542 13522
rect 8542 13470 8594 13522
rect 8594 13470 8596 13522
rect 8540 13468 8596 13470
rect 8126 13244 8182 13300
rect 6636 12236 6692 12292
rect 7036 12570 7092 12572
rect 7036 12518 7038 12570
rect 7038 12518 7090 12570
rect 7090 12518 7092 12570
rect 7036 12516 7092 12518
rect 7140 12570 7196 12572
rect 7140 12518 7142 12570
rect 7142 12518 7194 12570
rect 7194 12518 7196 12570
rect 7140 12516 7196 12518
rect 7244 12570 7300 12572
rect 7244 12518 7246 12570
rect 7246 12518 7298 12570
rect 7298 12518 7300 12570
rect 7244 12516 7300 12518
rect 6782 12164 6784 12180
rect 6784 12164 6836 12180
rect 6836 12164 6838 12180
rect 6782 12124 6838 12164
rect 7196 12124 7252 12180
rect 7420 12012 7476 12068
rect 6412 11452 6468 11508
rect 6860 11788 6916 11844
rect 6076 11228 6132 11284
rect 5292 10586 5294 10612
rect 5294 10586 5346 10612
rect 5346 10586 5348 10612
rect 5292 10556 5348 10586
rect 3612 10332 3668 10388
rect 4124 10218 4180 10220
rect 4124 10166 4126 10218
rect 4126 10166 4178 10218
rect 4178 10166 4180 10218
rect 4124 10164 4180 10166
rect 4228 10218 4284 10220
rect 4228 10166 4230 10218
rect 4230 10166 4282 10218
rect 4282 10166 4284 10218
rect 4228 10164 4284 10166
rect 4332 10218 4388 10220
rect 4332 10166 4334 10218
rect 4334 10166 4386 10218
rect 4386 10166 4388 10218
rect 4332 10164 4388 10166
rect 4124 8650 4180 8652
rect 4124 8598 4126 8650
rect 4126 8598 4178 8650
rect 4178 8598 4180 8650
rect 4124 8596 4180 8598
rect 4228 8650 4284 8652
rect 4228 8598 4230 8650
rect 4230 8598 4282 8650
rect 4282 8598 4284 8650
rect 4228 8596 4284 8598
rect 4332 8650 4388 8652
rect 4332 8598 4334 8650
rect 4334 8598 4386 8650
rect 4386 8598 4388 8650
rect 4332 8596 4388 8598
rect 5180 8316 5236 8372
rect 7036 11002 7092 11004
rect 7036 10950 7038 11002
rect 7038 10950 7090 11002
rect 7090 10950 7092 11002
rect 7036 10948 7092 10950
rect 7140 11002 7196 11004
rect 7140 10950 7142 11002
rect 7142 10950 7194 11002
rect 7194 10950 7196 11002
rect 7140 10948 7196 10950
rect 7244 11002 7300 11004
rect 7244 10950 7246 11002
rect 7246 10950 7298 11002
rect 7298 10950 7300 11002
rect 7420 11004 7476 11060
rect 7244 10948 7300 10950
rect 7308 10780 7364 10836
rect 6412 10556 6468 10612
rect 6692 10050 6748 10052
rect 6692 9998 6694 10050
rect 6694 9998 6746 10050
rect 6746 9998 6748 10050
rect 6692 9996 6748 9998
rect 6972 10444 7028 10500
rect 10052 15148 10108 15204
rect 10332 15314 10388 15316
rect 10332 15262 10334 15314
rect 10334 15262 10386 15314
rect 10386 15262 10388 15314
rect 10332 15260 10388 15262
rect 12348 18508 12404 18564
rect 12860 21978 12916 21980
rect 12860 21926 12862 21978
rect 12862 21926 12914 21978
rect 12914 21926 12916 21978
rect 12860 21924 12916 21926
rect 12964 21978 13020 21980
rect 12964 21926 12966 21978
rect 12966 21926 13018 21978
rect 13018 21926 13020 21978
rect 12964 21924 13020 21926
rect 13068 21978 13124 21980
rect 13068 21926 13070 21978
rect 13070 21926 13122 21978
rect 13122 21926 13124 21978
rect 13068 21924 13124 21926
rect 18684 21978 18740 21980
rect 18684 21926 18686 21978
rect 18686 21926 18738 21978
rect 18738 21926 18740 21978
rect 18684 21924 18740 21926
rect 18788 21978 18844 21980
rect 18788 21926 18790 21978
rect 18790 21926 18842 21978
rect 18842 21926 18844 21978
rect 18788 21924 18844 21926
rect 18892 21978 18948 21980
rect 18892 21926 18894 21978
rect 18894 21926 18946 21978
rect 18946 21926 18948 21978
rect 18892 21924 18948 21926
rect 20076 21868 20132 21924
rect 17836 21644 17892 21700
rect 13916 21474 13972 21476
rect 13916 21422 13918 21474
rect 13918 21422 13970 21474
rect 13970 21422 13972 21474
rect 13916 21420 13972 21422
rect 14812 21084 14868 21140
rect 14700 20748 14756 20804
rect 14812 20860 14868 20916
rect 15148 20802 15204 20804
rect 15148 20750 15150 20802
rect 15150 20750 15202 20802
rect 15202 20750 15204 20802
rect 15148 20748 15204 20750
rect 12860 20410 12916 20412
rect 12860 20358 12862 20410
rect 12862 20358 12914 20410
rect 12914 20358 12916 20410
rect 12860 20356 12916 20358
rect 12964 20410 13020 20412
rect 12964 20358 12966 20410
rect 12966 20358 13018 20410
rect 13018 20358 13020 20410
rect 12964 20356 13020 20358
rect 13068 20410 13124 20412
rect 13068 20358 13070 20410
rect 13070 20358 13122 20410
rect 13122 20358 13124 20410
rect 13068 20356 13124 20358
rect 13804 20076 13860 20132
rect 13580 19346 13636 19348
rect 13580 19294 13582 19346
rect 13582 19294 13634 19346
rect 13634 19294 13636 19346
rect 13580 19292 13636 19294
rect 13692 19180 13748 19236
rect 12860 18842 12916 18844
rect 12860 18790 12862 18842
rect 12862 18790 12914 18842
rect 12914 18790 12916 18842
rect 12860 18788 12916 18790
rect 12964 18842 13020 18844
rect 12964 18790 12966 18842
rect 12966 18790 13018 18842
rect 13018 18790 13020 18842
rect 12964 18788 13020 18790
rect 13068 18842 13124 18844
rect 13068 18790 13070 18842
rect 13070 18790 13122 18842
rect 13122 18790 13124 18842
rect 13068 18788 13124 18790
rect 12460 18396 12516 18452
rect 12908 18450 12964 18452
rect 12908 18398 12910 18450
rect 12910 18398 12962 18450
rect 12962 18398 12964 18450
rect 12908 18396 12964 18398
rect 12572 18226 12628 18228
rect 12572 18174 12574 18226
rect 12574 18174 12626 18226
rect 12626 18174 12628 18226
rect 12572 18172 12628 18174
rect 14140 20076 14196 20132
rect 15148 20076 15204 20132
rect 17276 21586 17332 21588
rect 17276 21534 17278 21586
rect 17278 21534 17330 21586
rect 17330 21534 17332 21586
rect 17276 21532 17332 21534
rect 15772 21194 15828 21196
rect 15772 21142 15774 21194
rect 15774 21142 15826 21194
rect 15826 21142 15828 21194
rect 15772 21140 15828 21142
rect 15876 21194 15932 21196
rect 15876 21142 15878 21194
rect 15878 21142 15930 21194
rect 15930 21142 15932 21194
rect 15876 21140 15932 21142
rect 15980 21194 16036 21196
rect 15980 21142 15982 21194
rect 15982 21142 16034 21194
rect 16034 21142 16036 21194
rect 15980 21140 16036 21142
rect 17836 20914 17892 20916
rect 17836 20862 17838 20914
rect 17838 20862 17890 20914
rect 17890 20862 17892 20914
rect 17836 20860 17892 20862
rect 17052 20748 17108 20804
rect 15772 19626 15828 19628
rect 15772 19574 15774 19626
rect 15774 19574 15826 19626
rect 15826 19574 15828 19626
rect 15772 19572 15828 19574
rect 15876 19626 15932 19628
rect 15876 19574 15878 19626
rect 15878 19574 15930 19626
rect 15930 19574 15932 19626
rect 15876 19572 15932 19574
rect 15980 19626 16036 19628
rect 15980 19574 15982 19626
rect 15982 19574 16034 19626
rect 16034 19574 16036 19626
rect 15980 19572 16036 19574
rect 18956 20802 19012 20804
rect 18956 20750 18958 20802
rect 18958 20750 19010 20802
rect 19010 20750 19012 20802
rect 18956 20748 19012 20750
rect 18684 20410 18740 20412
rect 18684 20358 18686 20410
rect 18686 20358 18738 20410
rect 18738 20358 18740 20410
rect 18684 20356 18740 20358
rect 18788 20410 18844 20412
rect 18788 20358 18790 20410
rect 18790 20358 18842 20410
rect 18842 20358 18844 20410
rect 18788 20356 18844 20358
rect 18892 20410 18948 20412
rect 18892 20358 18894 20410
rect 18894 20358 18946 20410
rect 18946 20358 18948 20410
rect 18892 20356 18948 20358
rect 19180 20300 19236 20356
rect 18396 20188 18452 20244
rect 19404 20018 19460 20020
rect 19404 19966 19406 20018
rect 19406 19966 19458 20018
rect 19458 19966 19460 20018
rect 19404 19964 19460 19966
rect 20076 20748 20132 20804
rect 20300 20972 20356 21028
rect 20412 20748 20468 20804
rect 19740 20188 19796 20244
rect 15484 19234 15540 19236
rect 15484 19182 15486 19234
rect 15486 19182 15538 19234
rect 15538 19182 15540 19234
rect 15484 19180 15540 19182
rect 14588 17778 14644 17780
rect 14588 17726 14590 17778
rect 14590 17726 14642 17778
rect 14642 17726 14644 17778
rect 14588 17724 14644 17726
rect 15148 17724 15204 17780
rect 12236 17666 12292 17668
rect 12236 17614 12238 17666
rect 12238 17614 12290 17666
rect 12290 17614 12292 17666
rect 12236 17612 12292 17614
rect 11788 16156 11844 16212
rect 12124 16828 12180 16884
rect 10780 15260 10836 15316
rect 11452 16098 11508 16100
rect 11452 16046 11454 16098
rect 11454 16046 11506 16098
rect 11506 16046 11508 16098
rect 11452 16044 11508 16046
rect 11732 15986 11788 15988
rect 11732 15934 11734 15986
rect 11734 15934 11786 15986
rect 11786 15934 11788 15986
rect 11732 15932 11788 15934
rect 11228 15260 11284 15316
rect 12860 17274 12916 17276
rect 12860 17222 12862 17274
rect 12862 17222 12914 17274
rect 12914 17222 12916 17274
rect 12860 17220 12916 17222
rect 12964 17274 13020 17276
rect 12964 17222 12966 17274
rect 12966 17222 13018 17274
rect 13018 17222 13020 17274
rect 12964 17220 13020 17222
rect 13068 17274 13124 17276
rect 13068 17222 13070 17274
rect 13070 17222 13122 17274
rect 13122 17222 13124 17274
rect 13068 17220 13124 17222
rect 12908 16882 12964 16884
rect 12908 16830 12910 16882
rect 12910 16830 12962 16882
rect 12962 16830 12964 16882
rect 12908 16828 12964 16830
rect 13412 16882 13468 16884
rect 13412 16830 13414 16882
rect 13414 16830 13466 16882
rect 13466 16830 13468 16882
rect 13412 16828 13468 16830
rect 14252 16828 14308 16884
rect 12236 16098 12292 16100
rect 12236 16046 12238 16098
rect 12238 16046 12290 16098
rect 12290 16046 12292 16098
rect 12236 16044 12292 16046
rect 12516 16098 12572 16100
rect 12516 16046 12518 16098
rect 12518 16046 12570 16098
rect 12570 16046 12572 16098
rect 12516 16044 12572 16046
rect 14700 16858 14702 16884
rect 14702 16858 14754 16884
rect 14754 16858 14756 16884
rect 14700 16828 14756 16858
rect 15772 18058 15828 18060
rect 15772 18006 15774 18058
rect 15774 18006 15826 18058
rect 15826 18006 15828 18058
rect 15772 18004 15828 18006
rect 15876 18058 15932 18060
rect 15876 18006 15878 18058
rect 15878 18006 15930 18058
rect 15930 18006 15932 18058
rect 15876 18004 15932 18006
rect 15980 18058 16036 18060
rect 15980 18006 15982 18058
rect 15982 18006 16034 18058
rect 16034 18006 16036 18058
rect 15980 18004 16036 18006
rect 18684 18842 18740 18844
rect 18684 18790 18686 18842
rect 18686 18790 18738 18842
rect 18738 18790 18740 18842
rect 18684 18788 18740 18790
rect 18788 18842 18844 18844
rect 18788 18790 18790 18842
rect 18790 18790 18842 18842
rect 18842 18790 18844 18842
rect 18788 18788 18844 18790
rect 18892 18842 18948 18844
rect 18892 18790 18894 18842
rect 18894 18790 18946 18842
rect 18946 18790 18948 18842
rect 18892 18788 18948 18790
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 14364 16098 14420 16100
rect 14364 16046 14366 16098
rect 14366 16046 14418 16098
rect 14418 16046 14420 16098
rect 14364 16044 14420 16046
rect 12860 15706 12916 15708
rect 12860 15654 12862 15706
rect 12862 15654 12914 15706
rect 12914 15654 12916 15706
rect 12860 15652 12916 15654
rect 12964 15706 13020 15708
rect 12964 15654 12966 15706
rect 12966 15654 13018 15706
rect 13018 15654 13020 15706
rect 12964 15652 13020 15654
rect 13068 15706 13124 15708
rect 13068 15654 13070 15706
rect 13070 15654 13122 15706
rect 13122 15654 13124 15706
rect 13068 15652 13124 15654
rect 12348 15538 12404 15540
rect 12348 15486 12350 15538
rect 12350 15486 12402 15538
rect 12402 15486 12404 15538
rect 12348 15484 12404 15486
rect 13580 15484 13636 15540
rect 10892 15202 10948 15204
rect 10892 15150 10894 15202
rect 10894 15150 10946 15202
rect 10946 15150 10948 15202
rect 10892 15148 10948 15150
rect 12012 15148 12068 15204
rect 9100 14252 9156 14308
rect 9212 13692 9268 13748
rect 8204 12236 8260 12292
rect 8316 12178 8372 12180
rect 8316 12126 8318 12178
rect 8318 12126 8370 12178
rect 8370 12126 8372 12178
rect 8316 12124 8372 12126
rect 8558 12178 8614 12180
rect 8558 12126 8560 12178
rect 8560 12126 8612 12178
rect 8612 12126 8614 12178
rect 8558 12124 8614 12126
rect 9948 14922 10004 14924
rect 9948 14870 9950 14922
rect 9950 14870 10002 14922
rect 10002 14870 10004 14922
rect 9948 14868 10004 14870
rect 10052 14922 10108 14924
rect 10052 14870 10054 14922
rect 10054 14870 10106 14922
rect 10106 14870 10108 14922
rect 10052 14868 10108 14870
rect 10156 14922 10212 14924
rect 10156 14870 10158 14922
rect 10158 14870 10210 14922
rect 10210 14870 10212 14922
rect 10156 14868 10212 14870
rect 11116 14364 11172 14420
rect 10948 13634 11004 13636
rect 10948 13582 10950 13634
rect 10950 13582 11002 13634
rect 11002 13582 11004 13634
rect 10948 13580 11004 13582
rect 10108 13468 10164 13524
rect 9948 13354 10004 13356
rect 9948 13302 9950 13354
rect 9950 13302 10002 13354
rect 10002 13302 10004 13354
rect 9948 13300 10004 13302
rect 10052 13354 10108 13356
rect 10052 13302 10054 13354
rect 10054 13302 10106 13354
rect 10106 13302 10108 13354
rect 10052 13300 10108 13302
rect 10156 13354 10212 13356
rect 10156 13302 10158 13354
rect 10158 13302 10210 13354
rect 10210 13302 10212 13354
rect 10156 13300 10212 13302
rect 9996 12348 10052 12404
rect 10668 12348 10724 12404
rect 10500 12236 10556 12292
rect 8092 12012 8148 12068
rect 9660 12178 9716 12180
rect 9660 12126 9662 12178
rect 9662 12126 9714 12178
rect 9714 12126 9716 12178
rect 9660 12124 9716 12126
rect 10332 12012 10388 12068
rect 7980 11228 8036 11284
rect 8428 11228 8484 11284
rect 7756 10780 7812 10836
rect 7308 9996 7364 10052
rect 7532 9996 7588 10052
rect 7644 10220 7700 10276
rect 7420 9884 7476 9940
rect 8652 9772 8708 9828
rect 7036 9434 7092 9436
rect 7036 9382 7038 9434
rect 7038 9382 7090 9434
rect 7090 9382 7092 9434
rect 7036 9380 7092 9382
rect 7140 9434 7196 9436
rect 7140 9382 7142 9434
rect 7142 9382 7194 9434
rect 7194 9382 7196 9434
rect 7140 9380 7196 9382
rect 7244 9434 7300 9436
rect 7244 9382 7246 9434
rect 7246 9382 7298 9434
rect 7298 9382 7300 9434
rect 7244 9380 7300 9382
rect 7644 8930 7700 8932
rect 7644 8878 7646 8930
rect 7646 8878 7698 8930
rect 7698 8878 7700 8930
rect 7644 8876 7700 8878
rect 7756 8764 7812 8820
rect 6860 8316 6916 8372
rect 7532 8316 7588 8372
rect 7036 7866 7092 7868
rect 7036 7814 7038 7866
rect 7038 7814 7090 7866
rect 7090 7814 7092 7866
rect 7036 7812 7092 7814
rect 7140 7866 7196 7868
rect 7140 7814 7142 7866
rect 7142 7814 7194 7866
rect 7194 7814 7196 7866
rect 7140 7812 7196 7814
rect 7244 7866 7300 7868
rect 7244 7814 7246 7866
rect 7246 7814 7298 7866
rect 7298 7814 7300 7866
rect 7244 7812 7300 7814
rect 4124 7082 4180 7084
rect 4124 7030 4126 7082
rect 4126 7030 4178 7082
rect 4178 7030 4180 7082
rect 4124 7028 4180 7030
rect 4228 7082 4284 7084
rect 4228 7030 4230 7082
rect 4230 7030 4282 7082
rect 4282 7030 4284 7082
rect 4228 7028 4284 7030
rect 4332 7082 4388 7084
rect 4332 7030 4334 7082
rect 4334 7030 4386 7082
rect 4386 7030 4388 7082
rect 4332 7028 4388 7030
rect 9660 11394 9716 11396
rect 9660 11342 9662 11394
rect 9662 11342 9714 11394
rect 9714 11342 9716 11394
rect 9660 11340 9716 11342
rect 9948 11786 10004 11788
rect 9948 11734 9950 11786
rect 9950 11734 10002 11786
rect 10002 11734 10004 11786
rect 9948 11732 10004 11734
rect 10052 11786 10108 11788
rect 10052 11734 10054 11786
rect 10054 11734 10106 11786
rect 10106 11734 10108 11786
rect 10052 11732 10108 11734
rect 10156 11786 10212 11788
rect 10156 11734 10158 11786
rect 10158 11734 10210 11786
rect 10210 11734 10212 11786
rect 10156 11732 10212 11734
rect 9948 10218 10004 10220
rect 9948 10166 9950 10218
rect 9950 10166 10002 10218
rect 10002 10166 10004 10218
rect 9948 10164 10004 10166
rect 10052 10218 10108 10220
rect 10052 10166 10054 10218
rect 10054 10166 10106 10218
rect 10106 10166 10108 10218
rect 10052 10164 10108 10166
rect 10156 10218 10212 10220
rect 10156 10166 10158 10218
rect 10158 10166 10210 10218
rect 10210 10166 10212 10218
rect 10156 10164 10212 10166
rect 8092 8540 8148 8596
rect 9884 9884 9940 9940
rect 10220 9772 10276 9828
rect 11396 13746 11452 13748
rect 11396 13694 11398 13746
rect 11398 13694 11450 13746
rect 11450 13694 11452 13746
rect 11396 13692 11452 13694
rect 11116 12348 11172 12404
rect 11788 13580 11844 13636
rect 11900 12236 11956 12292
rect 11004 12178 11060 12180
rect 11004 12126 11006 12178
rect 11006 12126 11058 12178
rect 11058 12126 11060 12178
rect 11004 12124 11060 12126
rect 13020 14530 13076 14532
rect 13020 14478 13022 14530
rect 13022 14478 13074 14530
rect 13074 14478 13076 14530
rect 13020 14476 13076 14478
rect 13468 14418 13524 14420
rect 13468 14366 13470 14418
rect 13470 14366 13522 14418
rect 13522 14366 13524 14418
rect 13468 14364 13524 14366
rect 12860 14138 12916 14140
rect 12860 14086 12862 14138
rect 12862 14086 12914 14138
rect 12914 14086 12916 14138
rect 12860 14084 12916 14086
rect 12964 14138 13020 14140
rect 12964 14086 12966 14138
rect 12966 14086 13018 14138
rect 13018 14086 13020 14138
rect 12964 14084 13020 14086
rect 13068 14138 13124 14140
rect 13068 14086 13070 14138
rect 13070 14086 13122 14138
rect 13122 14086 13124 14138
rect 13068 14084 13124 14086
rect 13804 14364 13860 14420
rect 13356 13132 13412 13188
rect 12860 12570 12916 12572
rect 12860 12518 12862 12570
rect 12862 12518 12914 12570
rect 12914 12518 12916 12570
rect 12860 12516 12916 12518
rect 12964 12570 13020 12572
rect 12964 12518 12966 12570
rect 12966 12518 13018 12570
rect 13018 12518 13020 12570
rect 12964 12516 13020 12518
rect 13068 12570 13124 12572
rect 13068 12518 13070 12570
rect 13070 12518 13122 12570
rect 13122 12518 13124 12570
rect 13068 12516 13124 12518
rect 13356 12402 13412 12404
rect 13356 12350 13358 12402
rect 13358 12350 13410 12402
rect 13410 12350 13412 12402
rect 13356 12348 13412 12350
rect 12012 12012 12068 12068
rect 11246 11676 11302 11732
rect 10892 11394 10948 11396
rect 10892 11342 10894 11394
rect 10894 11342 10946 11394
rect 10946 11342 10948 11394
rect 10892 11340 10948 11342
rect 12684 11676 12740 11732
rect 12348 9884 12404 9940
rect 12796 11116 12852 11172
rect 12860 11002 12916 11004
rect 12860 10950 12862 11002
rect 12862 10950 12914 11002
rect 12914 10950 12916 11002
rect 12860 10948 12916 10950
rect 12964 11002 13020 11004
rect 12964 10950 12966 11002
rect 12966 10950 13018 11002
rect 13018 10950 13020 11002
rect 12964 10948 13020 10950
rect 13068 11002 13124 11004
rect 13068 10950 13070 11002
rect 13070 10950 13122 11002
rect 13122 10950 13124 11002
rect 13068 10948 13124 10950
rect 13636 11116 13692 11172
rect 13636 9884 13692 9940
rect 10556 8818 10612 8820
rect 10556 8766 10558 8818
rect 10558 8766 10610 8818
rect 10610 8766 10612 8818
rect 10556 8764 10612 8766
rect 9948 8650 10004 8652
rect 9948 8598 9950 8650
rect 9950 8598 10002 8650
rect 10002 8598 10004 8650
rect 9948 8596 10004 8598
rect 10052 8650 10108 8652
rect 10052 8598 10054 8650
rect 10054 8598 10106 8650
rect 10106 8598 10108 8650
rect 10052 8596 10108 8598
rect 10156 8650 10212 8652
rect 10156 8598 10158 8650
rect 10158 8598 10210 8650
rect 10210 8598 10212 8650
rect 10156 8596 10212 8598
rect 9772 8316 9828 8372
rect 9548 7532 9604 7588
rect 7868 7362 7924 7364
rect 7868 7310 7870 7362
rect 7870 7310 7922 7362
rect 7922 7310 7924 7362
rect 7868 7308 7924 7310
rect 7036 6298 7092 6300
rect 7036 6246 7038 6298
rect 7038 6246 7090 6298
rect 7090 6246 7092 6298
rect 7036 6244 7092 6246
rect 7140 6298 7196 6300
rect 7140 6246 7142 6298
rect 7142 6246 7194 6298
rect 7194 6246 7196 6298
rect 7140 6244 7196 6246
rect 7244 6298 7300 6300
rect 7244 6246 7246 6298
rect 7246 6246 7298 6298
rect 7298 6246 7300 6298
rect 7244 6244 7300 6246
rect 4124 5514 4180 5516
rect 4124 5462 4126 5514
rect 4126 5462 4178 5514
rect 4178 5462 4180 5514
rect 4124 5460 4180 5462
rect 4228 5514 4284 5516
rect 4228 5462 4230 5514
rect 4230 5462 4282 5514
rect 4282 5462 4284 5514
rect 4228 5460 4284 5462
rect 4332 5514 4388 5516
rect 4332 5462 4334 5514
rect 4334 5462 4386 5514
rect 4386 5462 4388 5514
rect 4332 5460 4388 5462
rect 12860 9434 12916 9436
rect 12860 9382 12862 9434
rect 12862 9382 12914 9434
rect 12914 9382 12916 9434
rect 12860 9380 12916 9382
rect 12964 9434 13020 9436
rect 12964 9382 12966 9434
rect 12966 9382 13018 9434
rect 13018 9382 13020 9434
rect 12964 9380 13020 9382
rect 13068 9434 13124 9436
rect 13068 9382 13070 9434
rect 13070 9382 13122 9434
rect 13122 9382 13124 9434
rect 13068 9380 13124 9382
rect 12908 9154 12964 9156
rect 12908 9102 12910 9154
rect 12910 9102 12962 9154
rect 12962 9102 12964 9154
rect 12908 9100 12964 9102
rect 13244 9100 13300 9156
rect 12348 8316 12404 8372
rect 11116 7980 11172 8036
rect 11676 7980 11732 8036
rect 11284 7308 11340 7364
rect 9948 7082 10004 7084
rect 9948 7030 9950 7082
rect 9950 7030 10002 7082
rect 10002 7030 10004 7082
rect 9948 7028 10004 7030
rect 10052 7082 10108 7084
rect 10052 7030 10054 7082
rect 10054 7030 10106 7082
rect 10106 7030 10108 7082
rect 10052 7028 10108 7030
rect 10156 7082 10212 7084
rect 10156 7030 10158 7082
rect 10158 7030 10210 7082
rect 10210 7030 10212 7082
rect 10156 7028 10212 7030
rect 10220 6690 10276 6692
rect 10220 6638 10222 6690
rect 10222 6638 10274 6690
rect 10274 6638 10276 6690
rect 10220 6636 10276 6638
rect 12860 7866 12916 7868
rect 12860 7814 12862 7866
rect 12862 7814 12914 7866
rect 12914 7814 12916 7866
rect 12860 7812 12916 7814
rect 12964 7866 13020 7868
rect 12964 7814 12966 7866
rect 12966 7814 13018 7866
rect 13018 7814 13020 7866
rect 12964 7812 13020 7814
rect 13068 7866 13124 7868
rect 13068 7814 13070 7866
rect 13070 7814 13122 7866
rect 13122 7814 13124 7866
rect 13068 7812 13124 7814
rect 11844 6690 11900 6692
rect 11844 6638 11846 6690
rect 11846 6638 11898 6690
rect 11898 6638 11900 6690
rect 11844 6636 11900 6638
rect 11228 5906 11284 5908
rect 11228 5854 11230 5906
rect 11230 5854 11282 5906
rect 11282 5854 11284 5906
rect 11228 5852 11284 5854
rect 11770 5906 11826 5908
rect 11770 5854 11772 5906
rect 11772 5854 11824 5906
rect 11824 5854 11826 5906
rect 11770 5852 11826 5854
rect 9948 5514 10004 5516
rect 9948 5462 9950 5514
rect 9950 5462 10002 5514
rect 10002 5462 10004 5514
rect 9948 5460 10004 5462
rect 10052 5514 10108 5516
rect 10052 5462 10054 5514
rect 10054 5462 10106 5514
rect 10106 5462 10108 5514
rect 10052 5460 10108 5462
rect 10156 5514 10212 5516
rect 10156 5462 10158 5514
rect 10158 5462 10210 5514
rect 10210 5462 10212 5514
rect 10156 5460 10212 5462
rect 12590 6578 12646 6580
rect 12590 6526 12592 6578
rect 12592 6526 12644 6578
rect 12644 6526 12646 6578
rect 12590 6524 12646 6526
rect 12860 6298 12916 6300
rect 12860 6246 12862 6298
rect 12862 6246 12914 6298
rect 12914 6246 12916 6298
rect 12860 6244 12916 6246
rect 12964 6298 13020 6300
rect 12964 6246 12966 6298
rect 12966 6246 13018 6298
rect 13018 6246 13020 6298
rect 12964 6244 13020 6246
rect 13068 6298 13124 6300
rect 13068 6246 13070 6298
rect 13070 6246 13122 6298
rect 13122 6246 13124 6298
rect 13068 6244 13124 6246
rect 12684 6018 12740 6020
rect 12684 5966 12686 6018
rect 12686 5966 12738 6018
rect 12738 5966 12740 6018
rect 12684 5964 12740 5966
rect 14382 14530 14438 14532
rect 14382 14478 14384 14530
rect 14384 14478 14436 14530
rect 14436 14478 14438 14530
rect 14382 14476 14438 14478
rect 13916 11900 13972 11956
rect 15772 16490 15828 16492
rect 15772 16438 15774 16490
rect 15774 16438 15826 16490
rect 15826 16438 15828 16490
rect 15772 16436 15828 16438
rect 15876 16490 15932 16492
rect 15876 16438 15878 16490
rect 15878 16438 15930 16490
rect 15930 16438 15932 16490
rect 15876 16436 15932 16438
rect 15980 16490 16036 16492
rect 15980 16438 15982 16490
rect 15982 16438 16034 16490
rect 16034 16438 16036 16490
rect 15980 16436 16036 16438
rect 19516 19122 19572 19124
rect 19516 19070 19518 19122
rect 19518 19070 19570 19122
rect 19570 19070 19572 19122
rect 19516 19068 19572 19070
rect 20188 20018 20244 20020
rect 20188 19966 20190 20018
rect 20190 19966 20242 20018
rect 20242 19966 20244 20018
rect 20860 21586 20916 21588
rect 20860 21534 20862 21586
rect 20862 21534 20914 21586
rect 20914 21534 20916 21586
rect 20860 21532 20916 21534
rect 21084 20972 21140 21028
rect 20524 20130 20580 20132
rect 20524 20078 20526 20130
rect 20526 20078 20578 20130
rect 20578 20078 20580 20130
rect 20524 20076 20580 20078
rect 20636 20300 20692 20356
rect 20188 19964 20244 19966
rect 21532 21644 21588 21700
rect 21364 21026 21420 21028
rect 21364 20974 21366 21026
rect 21366 20974 21418 21026
rect 21418 20974 21420 21026
rect 21364 20972 21420 20974
rect 21596 21194 21652 21196
rect 21596 21142 21598 21194
rect 21598 21142 21650 21194
rect 21650 21142 21652 21194
rect 21596 21140 21652 21142
rect 21700 21194 21756 21196
rect 21700 21142 21702 21194
rect 21702 21142 21754 21194
rect 21754 21142 21756 21194
rect 21700 21140 21756 21142
rect 21804 21194 21860 21196
rect 21804 21142 21806 21194
rect 21806 21142 21858 21194
rect 21858 21142 21860 21194
rect 21804 21140 21860 21142
rect 21980 21196 22036 21252
rect 21868 20802 21924 20804
rect 21868 20750 21870 20802
rect 21870 20750 21922 20802
rect 21922 20750 21924 20802
rect 21868 20748 21924 20750
rect 21644 20300 21700 20356
rect 24508 21978 24564 21980
rect 24508 21926 24510 21978
rect 24510 21926 24562 21978
rect 24562 21926 24564 21978
rect 24508 21924 24564 21926
rect 24612 21978 24668 21980
rect 24612 21926 24614 21978
rect 24614 21926 24666 21978
rect 24666 21926 24668 21978
rect 24612 21924 24668 21926
rect 24716 21978 24772 21980
rect 24716 21926 24718 21978
rect 24718 21926 24770 21978
rect 24770 21926 24772 21978
rect 24716 21924 24772 21926
rect 23080 20802 23136 20804
rect 23080 20750 23082 20802
rect 23082 20750 23134 20802
rect 23134 20750 23136 20802
rect 23080 20748 23136 20750
rect 22876 20300 22932 20356
rect 23548 20076 23604 20132
rect 22988 19964 23044 20020
rect 22652 19852 22708 19908
rect 21596 19626 21652 19628
rect 21596 19574 21598 19626
rect 21598 19574 21650 19626
rect 21650 19574 21652 19626
rect 21596 19572 21652 19574
rect 21700 19626 21756 19628
rect 21700 19574 21702 19626
rect 21702 19574 21754 19626
rect 21754 19574 21756 19626
rect 21700 19572 21756 19574
rect 21804 19626 21860 19628
rect 21804 19574 21806 19626
rect 21806 19574 21858 19626
rect 21858 19574 21860 19626
rect 21804 19572 21860 19574
rect 19404 17500 19460 17556
rect 18684 17274 18740 17276
rect 18684 17222 18686 17274
rect 18686 17222 18738 17274
rect 18738 17222 18740 17274
rect 18684 17220 18740 17222
rect 18788 17274 18844 17276
rect 18788 17222 18790 17274
rect 18790 17222 18842 17274
rect 18842 17222 18844 17274
rect 18788 17220 18844 17222
rect 18892 17274 18948 17276
rect 18892 17222 18894 17274
rect 18894 17222 18946 17274
rect 18946 17222 18948 17274
rect 18892 17220 18948 17222
rect 18508 17052 18564 17108
rect 14924 14364 14980 14420
rect 15820 15090 15876 15092
rect 15820 15038 15822 15090
rect 15822 15038 15874 15090
rect 15874 15038 15876 15090
rect 15820 15036 15876 15038
rect 15772 14922 15828 14924
rect 15772 14870 15774 14922
rect 15774 14870 15826 14922
rect 15826 14870 15828 14922
rect 15772 14868 15828 14870
rect 15876 14922 15932 14924
rect 15876 14870 15878 14922
rect 15878 14870 15930 14922
rect 15930 14870 15932 14922
rect 15876 14868 15932 14870
rect 15980 14922 16036 14924
rect 15980 14870 15982 14922
rect 15982 14870 16034 14922
rect 16034 14870 16036 14922
rect 15980 14868 16036 14870
rect 20188 18396 20244 18452
rect 20636 19234 20692 19236
rect 20636 19182 20638 19234
rect 20638 19182 20690 19234
rect 20690 19182 20692 19234
rect 20636 19180 20692 19182
rect 20860 19068 20916 19124
rect 22876 19628 22932 19684
rect 21420 19190 21476 19236
rect 21420 19180 21422 19190
rect 21422 19180 21474 19190
rect 21474 19180 21476 19190
rect 21756 19234 21812 19236
rect 21756 19182 21758 19234
rect 21758 19182 21810 19234
rect 21810 19182 21812 19234
rect 21756 19180 21812 19182
rect 20076 17554 20132 17556
rect 20076 17502 20078 17554
rect 20078 17502 20130 17554
rect 20130 17502 20132 17554
rect 20076 17500 20132 17502
rect 20188 17052 20244 17108
rect 22036 18338 22092 18340
rect 22036 18286 22038 18338
rect 22038 18286 22090 18338
rect 22090 18286 22092 18338
rect 22036 18284 22092 18286
rect 23996 19628 24052 19684
rect 23436 19516 23492 19572
rect 23231 19234 23287 19236
rect 23231 19182 23233 19234
rect 23233 19182 23285 19234
rect 23285 19182 23287 19234
rect 23231 19180 23287 19182
rect 23100 18396 23156 18452
rect 24508 20410 24564 20412
rect 24508 20358 24510 20410
rect 24510 20358 24562 20410
rect 24562 20358 24564 20410
rect 24508 20356 24564 20358
rect 24612 20410 24668 20412
rect 24612 20358 24614 20410
rect 24614 20358 24666 20410
rect 24666 20358 24668 20410
rect 24612 20356 24668 20358
rect 24716 20410 24772 20412
rect 24716 20358 24718 20410
rect 24718 20358 24770 20410
rect 24770 20358 24772 20410
rect 24716 20356 24772 20358
rect 24892 19964 24948 20020
rect 24508 18842 24564 18844
rect 24508 18790 24510 18842
rect 24510 18790 24562 18842
rect 24562 18790 24564 18842
rect 24508 18788 24564 18790
rect 24612 18842 24668 18844
rect 24612 18790 24614 18842
rect 24614 18790 24666 18842
rect 24666 18790 24668 18842
rect 24612 18788 24668 18790
rect 24716 18842 24772 18844
rect 24716 18790 24718 18842
rect 24718 18790 24770 18842
rect 24770 18790 24772 18842
rect 24716 18788 24772 18790
rect 22764 18284 22820 18340
rect 21596 18058 21652 18060
rect 21596 18006 21598 18058
rect 21598 18006 21650 18058
rect 21650 18006 21652 18058
rect 21596 18004 21652 18006
rect 21700 18058 21756 18060
rect 21700 18006 21702 18058
rect 21702 18006 21754 18058
rect 21754 18006 21756 18058
rect 21700 18004 21756 18006
rect 21804 18058 21860 18060
rect 21804 18006 21806 18058
rect 21806 18006 21858 18058
rect 21858 18006 21860 18058
rect 22428 18060 22484 18116
rect 21804 18004 21860 18006
rect 22764 17948 22820 18004
rect 22092 17666 22148 17668
rect 22092 17614 22094 17666
rect 22094 17614 22146 17666
rect 22146 17614 22148 17666
rect 22092 17612 22148 17614
rect 22204 17500 22260 17556
rect 19740 16828 19796 16884
rect 19628 16604 19684 16660
rect 19292 16098 19348 16100
rect 19292 16046 19294 16098
rect 19294 16046 19346 16098
rect 19346 16046 19348 16098
rect 19292 16044 19348 16046
rect 20412 16857 20414 16884
rect 20414 16857 20466 16884
rect 20466 16857 20468 16884
rect 20412 16828 20468 16857
rect 20076 16604 20132 16660
rect 22968 17500 23024 17556
rect 23100 16940 23156 16996
rect 21596 16490 21652 16492
rect 21596 16438 21598 16490
rect 21598 16438 21650 16490
rect 21650 16438 21652 16490
rect 21596 16436 21652 16438
rect 21700 16490 21756 16492
rect 21700 16438 21702 16490
rect 21702 16438 21754 16490
rect 21754 16438 21756 16490
rect 21700 16436 21756 16438
rect 21804 16490 21860 16492
rect 21804 16438 21806 16490
rect 21806 16438 21858 16490
rect 21858 16438 21860 16490
rect 21804 16436 21860 16438
rect 20636 16098 20692 16100
rect 19180 15932 19236 15988
rect 18684 15706 18740 15708
rect 18684 15654 18686 15706
rect 18686 15654 18738 15706
rect 18738 15654 18740 15706
rect 18684 15652 18740 15654
rect 18788 15706 18844 15708
rect 18788 15654 18790 15706
rect 18790 15654 18842 15706
rect 18842 15654 18844 15706
rect 18788 15652 18844 15654
rect 18892 15706 18948 15708
rect 18892 15654 18894 15706
rect 18894 15654 18946 15706
rect 18946 15654 18948 15706
rect 18892 15652 18948 15654
rect 17052 15036 17108 15092
rect 14588 13020 14644 13076
rect 14830 12850 14886 12852
rect 14830 12798 14832 12850
rect 14832 12798 14884 12850
rect 14884 12798 14886 12850
rect 14830 12796 14886 12798
rect 18508 14924 18564 14980
rect 15772 13354 15828 13356
rect 15772 13302 15774 13354
rect 15774 13302 15826 13354
rect 15826 13302 15828 13354
rect 15772 13300 15828 13302
rect 15876 13354 15932 13356
rect 15876 13302 15878 13354
rect 15878 13302 15930 13354
rect 15930 13302 15932 13354
rect 15876 13300 15932 13302
rect 15980 13354 16036 13356
rect 15980 13302 15982 13354
rect 15982 13302 16034 13354
rect 16034 13302 16036 13354
rect 15980 13300 16036 13302
rect 18684 14138 18740 14140
rect 18684 14086 18686 14138
rect 18686 14086 18738 14138
rect 18738 14086 18740 14138
rect 18684 14084 18740 14086
rect 18788 14138 18844 14140
rect 18788 14086 18790 14138
rect 18790 14086 18842 14138
rect 18842 14086 18844 14138
rect 18788 14084 18844 14086
rect 18892 14138 18948 14140
rect 18892 14086 18894 14138
rect 18894 14086 18946 14138
rect 18946 14086 18948 14138
rect 18892 14084 18948 14086
rect 16716 13244 16772 13300
rect 17724 13244 17780 13300
rect 15372 13074 15428 13076
rect 15372 13022 15374 13074
rect 15374 13022 15426 13074
rect 15426 13022 15428 13074
rect 15372 13020 15428 13022
rect 15036 12124 15092 12180
rect 15596 12796 15652 12852
rect 15932 12402 15988 12404
rect 15932 12350 15934 12402
rect 15934 12350 15986 12402
rect 15986 12350 15988 12402
rect 15932 12348 15988 12350
rect 17276 12348 17332 12404
rect 14700 11954 14756 11956
rect 14700 11902 14702 11954
rect 14702 11902 14754 11954
rect 14754 11902 14756 11954
rect 14700 11900 14756 11902
rect 15772 11786 15828 11788
rect 15772 11734 15774 11786
rect 15774 11734 15826 11786
rect 15826 11734 15828 11786
rect 15772 11732 15828 11734
rect 15876 11786 15932 11788
rect 15876 11734 15878 11786
rect 15878 11734 15930 11786
rect 15930 11734 15932 11786
rect 15876 11732 15932 11734
rect 15980 11786 16036 11788
rect 15980 11734 15982 11786
rect 15982 11734 16034 11786
rect 16034 11734 16036 11786
rect 15980 11732 16036 11734
rect 14140 10610 14196 10612
rect 14140 10558 14142 10610
rect 14142 10558 14194 10610
rect 14194 10558 14196 10610
rect 14140 10556 14196 10558
rect 15260 11228 15316 11284
rect 15260 10556 15316 10612
rect 14140 9826 14196 9828
rect 14140 9774 14142 9826
rect 14142 9774 14194 9826
rect 14194 9774 14196 9826
rect 14140 9772 14196 9774
rect 16044 11282 16100 11284
rect 16044 11230 16046 11282
rect 16046 11230 16098 11282
rect 16098 11230 16100 11282
rect 16044 11228 16100 11230
rect 16268 10834 16324 10836
rect 16268 10782 16270 10834
rect 16270 10782 16322 10834
rect 16322 10782 16324 10834
rect 16268 10780 16324 10782
rect 19964 15314 20020 15316
rect 19964 15262 19966 15314
rect 19966 15262 20018 15314
rect 20018 15262 20020 15314
rect 19964 15260 20020 15262
rect 20188 15372 20244 15428
rect 20636 16046 20638 16098
rect 20638 16046 20690 16098
rect 20690 16046 20692 16098
rect 20636 16044 20692 16046
rect 21084 16044 21140 16100
rect 20076 15148 20132 15204
rect 20356 14754 20412 14756
rect 20356 14702 20358 14754
rect 20358 14702 20410 14754
rect 20410 14702 20412 14754
rect 20356 14700 20412 14702
rect 20860 15314 20916 15316
rect 20860 15262 20862 15314
rect 20862 15262 20914 15314
rect 20914 15262 20916 15314
rect 20860 15260 20916 15262
rect 20524 14700 20580 14756
rect 21756 16044 21812 16100
rect 21252 15426 21308 15428
rect 21252 15374 21254 15426
rect 21254 15374 21306 15426
rect 21306 15374 21308 15426
rect 21252 15372 21308 15374
rect 21980 15820 22036 15876
rect 22428 16044 22484 16100
rect 21756 15314 21812 15316
rect 21756 15262 21758 15314
rect 21758 15262 21810 15314
rect 21810 15262 21812 15314
rect 21756 15260 21812 15262
rect 22540 15260 22596 15316
rect 23996 18450 24052 18452
rect 23996 18398 23998 18450
rect 23998 18398 24050 18450
rect 24050 18398 24052 18450
rect 23996 18396 24052 18398
rect 23660 16882 23716 16884
rect 23660 16830 23662 16882
rect 23662 16830 23714 16882
rect 23714 16830 23716 16882
rect 23660 16828 23716 16830
rect 22783 16098 22839 16100
rect 22783 16046 22785 16098
rect 22785 16046 22837 16098
rect 22837 16046 22839 16098
rect 22783 16044 22839 16046
rect 22652 15148 22708 15204
rect 22764 15820 22820 15876
rect 21596 14922 21652 14924
rect 21596 14870 21598 14922
rect 21598 14870 21650 14922
rect 21650 14870 21652 14922
rect 21596 14868 21652 14870
rect 21700 14922 21756 14924
rect 21700 14870 21702 14922
rect 21702 14870 21754 14922
rect 21754 14870 21756 14922
rect 21700 14868 21756 14870
rect 21804 14922 21860 14924
rect 21804 14870 21806 14922
rect 21806 14870 21858 14922
rect 21858 14870 21860 14922
rect 21804 14868 21860 14870
rect 21420 14700 21476 14756
rect 20860 13746 20916 13748
rect 20860 13694 20862 13746
rect 20862 13694 20914 13746
rect 20914 13694 20916 13746
rect 20860 13692 20916 13694
rect 20636 13580 20692 13636
rect 19404 13356 19460 13412
rect 18684 12570 18740 12572
rect 18684 12518 18686 12570
rect 18686 12518 18738 12570
rect 18738 12518 18740 12570
rect 18684 12516 18740 12518
rect 18788 12570 18844 12572
rect 18788 12518 18790 12570
rect 18790 12518 18842 12570
rect 18842 12518 18844 12570
rect 18788 12516 18844 12518
rect 18892 12570 18948 12572
rect 18892 12518 18894 12570
rect 18894 12518 18946 12570
rect 18946 12518 18948 12570
rect 18892 12516 18948 12518
rect 21084 12796 21140 12852
rect 21308 13746 21364 13748
rect 21308 13694 21310 13746
rect 21310 13694 21362 13746
rect 21362 13694 21364 13746
rect 21308 13692 21364 13694
rect 21644 13580 21700 13636
rect 22204 13580 22260 13636
rect 21420 13468 21476 13524
rect 21596 13354 21652 13356
rect 21596 13302 21598 13354
rect 21598 13302 21650 13354
rect 21650 13302 21652 13354
rect 21596 13300 21652 13302
rect 21700 13354 21756 13356
rect 21700 13302 21702 13354
rect 21702 13302 21754 13354
rect 21754 13302 21756 13354
rect 21700 13300 21756 13302
rect 21804 13354 21860 13356
rect 21804 13302 21806 13354
rect 21806 13302 21858 13354
rect 21858 13302 21860 13354
rect 21804 13300 21860 13302
rect 23548 15314 23604 15316
rect 23548 15262 23550 15314
rect 23550 15262 23602 15314
rect 23602 15262 23604 15314
rect 23548 15260 23604 15262
rect 22988 15202 23044 15204
rect 22988 15150 22990 15202
rect 22990 15150 23042 15202
rect 23042 15150 23044 15202
rect 22988 15148 23044 15150
rect 23212 15148 23268 15204
rect 24508 17274 24564 17276
rect 24508 17222 24510 17274
rect 24510 17222 24562 17274
rect 24562 17222 24564 17274
rect 24508 17220 24564 17222
rect 24612 17274 24668 17276
rect 24612 17222 24614 17274
rect 24614 17222 24666 17274
rect 24666 17222 24668 17274
rect 24612 17220 24668 17222
rect 24716 17274 24772 17276
rect 24716 17222 24718 17274
rect 24718 17222 24770 17274
rect 24770 17222 24772 17274
rect 24716 17220 24772 17222
rect 24276 15986 24332 15988
rect 24276 15934 24278 15986
rect 24278 15934 24330 15986
rect 24330 15934 24332 15986
rect 24276 15932 24332 15934
rect 25004 16828 25060 16884
rect 24508 15706 24564 15708
rect 24508 15654 24510 15706
rect 24510 15654 24562 15706
rect 24562 15654 24564 15706
rect 24508 15652 24564 15654
rect 24612 15706 24668 15708
rect 24612 15654 24614 15706
rect 24614 15654 24666 15706
rect 24666 15654 24668 15706
rect 24612 15652 24668 15654
rect 24716 15706 24772 15708
rect 24716 15654 24718 15706
rect 24718 15654 24770 15706
rect 24770 15654 24772 15706
rect 24716 15652 24772 15654
rect 24108 15148 24164 15204
rect 23604 13970 23660 13972
rect 23604 13918 23606 13970
rect 23606 13918 23658 13970
rect 23658 13918 23660 13970
rect 23604 13916 23660 13918
rect 23772 13916 23828 13972
rect 23100 13746 23156 13748
rect 23100 13694 23102 13746
rect 23102 13694 23154 13746
rect 23154 13694 23156 13746
rect 23100 13692 23156 13694
rect 24508 14138 24564 14140
rect 24508 14086 24510 14138
rect 24510 14086 24562 14138
rect 24562 14086 24564 14138
rect 24508 14084 24564 14086
rect 24612 14138 24668 14140
rect 24612 14086 24614 14138
rect 24614 14086 24666 14138
rect 24666 14086 24668 14138
rect 24612 14084 24668 14086
rect 24716 14138 24772 14140
rect 24716 14086 24718 14138
rect 24718 14086 24770 14138
rect 24770 14086 24772 14138
rect 24716 14084 24772 14086
rect 23436 12962 23492 12964
rect 23436 12910 23438 12962
rect 23438 12910 23490 12962
rect 23490 12910 23492 12962
rect 23436 12908 23492 12910
rect 23996 12962 24052 12964
rect 23996 12910 23998 12962
rect 23998 12910 24050 12962
rect 24050 12910 24052 12962
rect 23996 12908 24052 12910
rect 22559 12796 22615 12852
rect 17948 10780 18004 10836
rect 18684 11002 18740 11004
rect 18684 10950 18686 11002
rect 18686 10950 18738 11002
rect 18738 10950 18740 11002
rect 18684 10948 18740 10950
rect 18788 11002 18844 11004
rect 18788 10950 18790 11002
rect 18790 10950 18842 11002
rect 18842 10950 18844 11002
rect 18788 10948 18844 10950
rect 18892 11002 18948 11004
rect 18892 10950 18894 11002
rect 18894 10950 18946 11002
rect 18946 10950 18948 11002
rect 18892 10948 18948 10950
rect 15772 10218 15828 10220
rect 15772 10166 15774 10218
rect 15774 10166 15826 10218
rect 15826 10166 15828 10218
rect 15772 10164 15828 10166
rect 15876 10218 15932 10220
rect 15876 10166 15878 10218
rect 15878 10166 15930 10218
rect 15930 10166 15932 10218
rect 15876 10164 15932 10166
rect 15980 10218 16036 10220
rect 15980 10166 15982 10218
rect 15982 10166 16034 10218
rect 16034 10166 16036 10218
rect 15980 10164 16036 10166
rect 15484 9826 15540 9828
rect 13804 9100 13860 9156
rect 15484 9774 15486 9826
rect 15486 9774 15538 9826
rect 15538 9774 15540 9826
rect 15484 9772 15540 9774
rect 16492 9826 16548 9828
rect 16492 9774 16494 9826
rect 16494 9774 16546 9826
rect 16546 9774 16548 9826
rect 16492 9772 16548 9774
rect 13748 8876 13804 8932
rect 13468 8316 13524 8372
rect 16604 9266 16660 9268
rect 16604 9214 16606 9266
rect 16606 9214 16658 9266
rect 16658 9214 16660 9266
rect 16604 9212 16660 9214
rect 18396 9212 18452 9268
rect 15772 8650 15828 8652
rect 15772 8598 15774 8650
rect 15774 8598 15826 8650
rect 15826 8598 15828 8650
rect 15772 8596 15828 8598
rect 15876 8650 15932 8652
rect 15876 8598 15878 8650
rect 15878 8598 15930 8650
rect 15930 8598 15932 8650
rect 15876 8596 15932 8598
rect 15980 8650 16036 8652
rect 15980 8598 15982 8650
rect 15982 8598 16034 8650
rect 16034 8598 16036 8650
rect 15980 8596 16036 8598
rect 19852 11788 19908 11844
rect 22092 12012 22148 12068
rect 21596 11786 21652 11788
rect 21596 11734 21598 11786
rect 21598 11734 21650 11786
rect 21650 11734 21652 11786
rect 21596 11732 21652 11734
rect 21700 11786 21756 11788
rect 21700 11734 21702 11786
rect 21702 11734 21754 11786
rect 21754 11734 21756 11786
rect 21700 11732 21756 11734
rect 21804 11786 21860 11788
rect 21804 11734 21806 11786
rect 21806 11734 21858 11786
rect 21858 11734 21860 11786
rect 21804 11732 21860 11734
rect 21756 11452 21812 11508
rect 22876 11564 22932 11620
rect 22988 12124 23044 12180
rect 23212 12236 23268 12292
rect 24052 12236 24108 12292
rect 22652 11452 22708 11508
rect 23324 11506 23380 11508
rect 23324 11454 23326 11506
rect 23326 11454 23378 11506
rect 23378 11454 23380 11506
rect 23324 11452 23380 11454
rect 23884 12178 23940 12180
rect 23884 12126 23886 12178
rect 23886 12126 23938 12178
rect 23938 12126 23940 12178
rect 23884 12124 23940 12126
rect 24508 12570 24564 12572
rect 24508 12518 24510 12570
rect 24510 12518 24562 12570
rect 24562 12518 24564 12570
rect 24508 12516 24564 12518
rect 24612 12570 24668 12572
rect 24612 12518 24614 12570
rect 24614 12518 24666 12570
rect 24666 12518 24668 12570
rect 24612 12516 24668 12518
rect 24716 12570 24772 12572
rect 24716 12518 24718 12570
rect 24718 12518 24770 12570
rect 24770 12518 24772 12570
rect 24716 12516 24772 12518
rect 24276 11900 24332 11956
rect 23660 11564 23716 11620
rect 21596 10218 21652 10220
rect 21596 10166 21598 10218
rect 21598 10166 21650 10218
rect 21650 10166 21652 10218
rect 21596 10164 21652 10166
rect 21700 10218 21756 10220
rect 21700 10166 21702 10218
rect 21702 10166 21754 10218
rect 21754 10166 21756 10218
rect 21700 10164 21756 10166
rect 21804 10218 21860 10220
rect 21804 10166 21806 10218
rect 21806 10166 21858 10218
rect 21858 10166 21860 10218
rect 21804 10164 21860 10166
rect 24508 11002 24564 11004
rect 24508 10950 24510 11002
rect 24510 10950 24562 11002
rect 24562 10950 24564 11002
rect 24508 10948 24564 10950
rect 24612 11002 24668 11004
rect 24612 10950 24614 11002
rect 24614 10950 24666 11002
rect 24666 10950 24668 11002
rect 24612 10948 24668 10950
rect 24716 11002 24772 11004
rect 24716 10950 24718 11002
rect 24718 10950 24770 11002
rect 24770 10950 24772 11002
rect 24716 10948 24772 10950
rect 22260 10108 22316 10164
rect 21420 9884 21476 9940
rect 21980 9938 22036 9940
rect 21980 9886 21982 9938
rect 21982 9886 22034 9938
rect 22034 9886 22036 9938
rect 21980 9884 22036 9886
rect 19180 9548 19236 9604
rect 18684 9434 18740 9436
rect 18684 9382 18686 9434
rect 18686 9382 18738 9434
rect 18738 9382 18740 9434
rect 18684 9380 18740 9382
rect 18788 9434 18844 9436
rect 18788 9382 18790 9434
rect 18790 9382 18842 9434
rect 18842 9382 18844 9434
rect 18788 9380 18844 9382
rect 18892 9434 18948 9436
rect 18892 9382 18894 9434
rect 18894 9382 18946 9434
rect 18946 9382 18948 9434
rect 18892 9380 18948 9382
rect 14364 8316 14420 8372
rect 14924 8316 14980 8372
rect 15708 8370 15764 8372
rect 15708 8318 15710 8370
rect 15710 8318 15762 8370
rect 15762 8318 15764 8370
rect 15708 8316 15764 8318
rect 21196 9548 21252 9604
rect 23343 9548 23399 9604
rect 21596 8650 21652 8652
rect 21596 8598 21598 8650
rect 21598 8598 21650 8650
rect 21650 8598 21652 8650
rect 21596 8596 21652 8598
rect 21700 8650 21756 8652
rect 21700 8598 21702 8650
rect 21702 8598 21754 8650
rect 21754 8598 21756 8650
rect 21700 8596 21756 8598
rect 21804 8650 21860 8652
rect 21804 8598 21806 8650
rect 21806 8598 21858 8650
rect 21858 8598 21860 8650
rect 21804 8596 21860 8598
rect 13636 7532 13692 7588
rect 16156 7698 16212 7700
rect 16156 7646 16158 7698
rect 16158 7646 16210 7698
rect 16210 7646 16212 7698
rect 16156 7644 16212 7646
rect 17612 7644 17668 7700
rect 18684 7866 18740 7868
rect 18684 7814 18686 7866
rect 18686 7814 18738 7866
rect 18738 7814 18740 7866
rect 18684 7812 18740 7814
rect 18788 7866 18844 7868
rect 18788 7814 18790 7866
rect 18790 7814 18842 7866
rect 18842 7814 18844 7866
rect 18788 7812 18844 7814
rect 18892 7866 18948 7868
rect 18892 7814 18894 7866
rect 18894 7814 18946 7866
rect 18946 7814 18948 7866
rect 18892 7812 18948 7814
rect 15772 7082 15828 7084
rect 15772 7030 15774 7082
rect 15774 7030 15826 7082
rect 15826 7030 15828 7082
rect 15772 7028 15828 7030
rect 15876 7082 15932 7084
rect 15876 7030 15878 7082
rect 15878 7030 15930 7082
rect 15930 7030 15932 7082
rect 15876 7028 15932 7030
rect 15980 7082 16036 7084
rect 15980 7030 15982 7082
rect 15982 7030 16034 7082
rect 16034 7030 16036 7082
rect 15980 7028 16036 7030
rect 13356 6524 13412 6580
rect 13244 6018 13300 6020
rect 13244 5966 13246 6018
rect 13246 5966 13298 6018
rect 13298 5966 13300 6018
rect 13244 5964 13300 5966
rect 14700 6748 14756 6804
rect 15820 6802 15876 6804
rect 15820 6750 15822 6802
rect 15822 6750 15874 6802
rect 15874 6750 15876 6802
rect 15820 6748 15876 6750
rect 18732 7474 18788 7476
rect 18732 7422 18734 7474
rect 18734 7422 18786 7474
rect 18786 7422 18788 7474
rect 18732 7420 18788 7422
rect 16716 6412 16772 6468
rect 18284 6412 18340 6468
rect 15772 5514 15828 5516
rect 15772 5462 15774 5514
rect 15774 5462 15826 5514
rect 15826 5462 15828 5514
rect 15772 5460 15828 5462
rect 15876 5514 15932 5516
rect 15876 5462 15878 5514
rect 15878 5462 15930 5514
rect 15930 5462 15932 5514
rect 15876 5460 15932 5462
rect 15980 5514 16036 5516
rect 15980 5462 15982 5514
rect 15982 5462 16034 5514
rect 16034 5462 16036 5514
rect 15980 5460 16036 5462
rect 19964 8243 20020 8260
rect 19964 8204 19966 8243
rect 19966 8204 20018 8243
rect 20018 8204 20020 8243
rect 22092 8204 22148 8260
rect 21644 7644 21700 7700
rect 19852 7420 19908 7476
rect 21980 7532 22036 7588
rect 21596 7082 21652 7084
rect 21596 7030 21598 7082
rect 21598 7030 21650 7082
rect 21650 7030 21652 7082
rect 21596 7028 21652 7030
rect 21700 7082 21756 7084
rect 21700 7030 21702 7082
rect 21702 7030 21754 7082
rect 21754 7030 21756 7082
rect 21700 7028 21756 7030
rect 21804 7082 21860 7084
rect 21804 7030 21806 7082
rect 21806 7030 21858 7082
rect 21858 7030 21860 7082
rect 21804 7028 21860 7030
rect 18956 6412 19012 6468
rect 18684 6298 18740 6300
rect 18684 6246 18686 6298
rect 18686 6246 18738 6298
rect 18738 6246 18740 6298
rect 18684 6244 18740 6246
rect 18788 6298 18844 6300
rect 18788 6246 18790 6298
rect 18790 6246 18842 6298
rect 18842 6246 18844 6298
rect 18788 6244 18844 6246
rect 18892 6298 18948 6300
rect 18892 6246 18894 6298
rect 18894 6246 18946 6298
rect 18946 6246 18948 6298
rect 18892 6244 18948 6246
rect 18751 6076 18807 6132
rect 19628 5964 19684 6020
rect 18284 5068 18340 5124
rect 20300 6076 20356 6132
rect 7036 4730 7092 4732
rect 7036 4678 7038 4730
rect 7038 4678 7090 4730
rect 7090 4678 7092 4730
rect 7036 4676 7092 4678
rect 7140 4730 7196 4732
rect 7140 4678 7142 4730
rect 7142 4678 7194 4730
rect 7194 4678 7196 4730
rect 7140 4676 7196 4678
rect 7244 4730 7300 4732
rect 7244 4678 7246 4730
rect 7246 4678 7298 4730
rect 7298 4678 7300 4730
rect 7244 4676 7300 4678
rect 12860 4730 12916 4732
rect 12860 4678 12862 4730
rect 12862 4678 12914 4730
rect 12914 4678 12916 4730
rect 12860 4676 12916 4678
rect 12964 4730 13020 4732
rect 12964 4678 12966 4730
rect 12966 4678 13018 4730
rect 13018 4678 13020 4730
rect 12964 4676 13020 4678
rect 13068 4730 13124 4732
rect 13068 4678 13070 4730
rect 13070 4678 13122 4730
rect 13122 4678 13124 4730
rect 13068 4676 13124 4678
rect 18684 4730 18740 4732
rect 18684 4678 18686 4730
rect 18686 4678 18738 4730
rect 18738 4678 18740 4730
rect 18684 4676 18740 4678
rect 18788 4730 18844 4732
rect 18788 4678 18790 4730
rect 18790 4678 18842 4730
rect 18842 4678 18844 4730
rect 18788 4676 18844 4678
rect 18892 4730 18948 4732
rect 18892 4678 18894 4730
rect 18894 4678 18946 4730
rect 18946 4678 18948 4730
rect 18892 4676 18948 4678
rect 20188 5740 20244 5796
rect 20300 5628 20356 5684
rect 20804 6076 20860 6132
rect 20972 5852 21028 5908
rect 21420 5906 21476 5908
rect 21420 5854 21422 5906
rect 21422 5854 21474 5906
rect 21474 5854 21476 5906
rect 21420 5852 21476 5854
rect 21196 5740 21252 5796
rect 21756 5794 21812 5796
rect 21756 5742 21758 5794
rect 21758 5742 21810 5794
rect 21810 5742 21812 5794
rect 21756 5740 21812 5742
rect 21980 6412 22036 6468
rect 21084 5628 21140 5684
rect 22092 5964 22148 6020
rect 23772 10108 23828 10164
rect 23548 9548 23604 9604
rect 23884 9548 23940 9604
rect 24508 9434 24564 9436
rect 24508 9382 24510 9434
rect 24510 9382 24562 9434
rect 24562 9382 24564 9434
rect 24508 9380 24564 9382
rect 24612 9434 24668 9436
rect 24612 9382 24614 9434
rect 24614 9382 24666 9434
rect 24666 9382 24668 9434
rect 24612 9380 24668 9382
rect 24716 9434 24772 9436
rect 24716 9382 24718 9434
rect 24718 9382 24770 9434
rect 24770 9382 24772 9434
rect 24716 9380 24772 9382
rect 22428 7532 22484 7588
rect 23100 8370 23156 8372
rect 23100 8318 23102 8370
rect 23102 8318 23154 8370
rect 23154 8318 23156 8370
rect 23100 8316 23156 8318
rect 23100 7644 23156 7700
rect 22652 6188 22708 6244
rect 22204 5852 22260 5908
rect 24892 8316 24948 8372
rect 23343 7644 23399 7700
rect 23772 7644 23828 7700
rect 24508 7866 24564 7868
rect 24508 7814 24510 7866
rect 24510 7814 24562 7866
rect 24562 7814 24564 7866
rect 24508 7812 24564 7814
rect 24612 7866 24668 7868
rect 24612 7814 24614 7866
rect 24614 7814 24666 7866
rect 24666 7814 24668 7866
rect 24612 7812 24668 7814
rect 24716 7866 24772 7868
rect 24716 7814 24718 7866
rect 24718 7814 24770 7866
rect 24770 7814 24772 7866
rect 24716 7812 24772 7814
rect 23212 6860 23268 6916
rect 23884 6860 23940 6916
rect 22876 6466 22932 6468
rect 22876 6414 22878 6466
rect 22878 6414 22930 6466
rect 22930 6414 22932 6466
rect 22876 6412 22932 6414
rect 22559 5964 22615 6020
rect 23436 5906 23492 5908
rect 23436 5854 23438 5906
rect 23438 5854 23490 5906
rect 23490 5854 23492 5906
rect 23436 5852 23492 5854
rect 21980 5628 22036 5684
rect 21596 5514 21652 5516
rect 21596 5462 21598 5514
rect 21598 5462 21650 5514
rect 21650 5462 21652 5514
rect 21596 5460 21652 5462
rect 21700 5514 21756 5516
rect 21700 5462 21702 5514
rect 21702 5462 21754 5514
rect 21754 5462 21756 5514
rect 21700 5460 21756 5462
rect 21804 5514 21860 5516
rect 21804 5462 21806 5514
rect 21806 5462 21858 5514
rect 21858 5462 21860 5514
rect 21804 5460 21860 5462
rect 20972 5180 21028 5236
rect 19404 4508 19460 4564
rect 22428 5292 22484 5348
rect 21308 5068 21364 5124
rect 21532 5068 21588 5124
rect 22092 4338 22148 4340
rect 22092 4286 22094 4338
rect 22094 4286 22146 4338
rect 22146 4286 22148 4338
rect 22092 4284 22148 4286
rect 22540 5122 22596 5124
rect 22540 5070 22542 5122
rect 22542 5070 22594 5122
rect 22594 5070 22596 5122
rect 22540 5068 22596 5070
rect 23324 5234 23380 5236
rect 23324 5182 23326 5234
rect 23326 5182 23378 5234
rect 23378 5182 23380 5234
rect 23324 5180 23380 5182
rect 23660 5122 23716 5124
rect 23660 5070 23662 5122
rect 23662 5070 23714 5122
rect 23714 5070 23716 5122
rect 23660 5068 23716 5070
rect 4124 3946 4180 3948
rect 4124 3894 4126 3946
rect 4126 3894 4178 3946
rect 4178 3894 4180 3946
rect 4124 3892 4180 3894
rect 4228 3946 4284 3948
rect 4228 3894 4230 3946
rect 4230 3894 4282 3946
rect 4282 3894 4284 3946
rect 4228 3892 4284 3894
rect 4332 3946 4388 3948
rect 4332 3894 4334 3946
rect 4334 3894 4386 3946
rect 4386 3894 4388 3946
rect 4332 3892 4388 3894
rect 9948 3946 10004 3948
rect 9948 3894 9950 3946
rect 9950 3894 10002 3946
rect 10002 3894 10004 3946
rect 9948 3892 10004 3894
rect 10052 3946 10108 3948
rect 10052 3894 10054 3946
rect 10054 3894 10106 3946
rect 10106 3894 10108 3946
rect 10052 3892 10108 3894
rect 10156 3946 10212 3948
rect 10156 3894 10158 3946
rect 10158 3894 10210 3946
rect 10210 3894 10212 3946
rect 10156 3892 10212 3894
rect 15772 3946 15828 3948
rect 15772 3894 15774 3946
rect 15774 3894 15826 3946
rect 15826 3894 15828 3946
rect 15772 3892 15828 3894
rect 15876 3946 15932 3948
rect 15876 3894 15878 3946
rect 15878 3894 15930 3946
rect 15930 3894 15932 3946
rect 15876 3892 15932 3894
rect 15980 3946 16036 3948
rect 15980 3894 15982 3946
rect 15982 3894 16034 3946
rect 16034 3894 16036 3946
rect 15980 3892 16036 3894
rect 21596 3946 21652 3948
rect 21596 3894 21598 3946
rect 21598 3894 21650 3946
rect 21650 3894 21652 3946
rect 21596 3892 21652 3894
rect 21700 3946 21756 3948
rect 21700 3894 21702 3946
rect 21702 3894 21754 3946
rect 21754 3894 21756 3946
rect 21700 3892 21756 3894
rect 21804 3946 21860 3948
rect 21804 3894 21806 3946
rect 21806 3894 21858 3946
rect 21858 3894 21860 3946
rect 21804 3892 21860 3894
rect 23192 3948 23248 4004
rect 23996 5852 24052 5908
rect 24508 6298 24564 6300
rect 24220 5852 24276 5908
rect 23996 5292 24052 5348
rect 23996 3948 24052 4004
rect 24332 6188 24388 6244
rect 24508 6246 24510 6298
rect 24510 6246 24562 6298
rect 24562 6246 24564 6298
rect 24508 6244 24564 6246
rect 24612 6298 24668 6300
rect 24612 6246 24614 6298
rect 24614 6246 24666 6298
rect 24666 6246 24668 6298
rect 24612 6244 24668 6246
rect 24716 6298 24772 6300
rect 24716 6246 24718 6298
rect 24718 6246 24770 6298
rect 24770 6246 24772 6298
rect 24716 6244 24772 6246
rect 25004 5180 25060 5236
rect 24508 4730 24564 4732
rect 24508 4678 24510 4730
rect 24510 4678 24562 4730
rect 24562 4678 24564 4730
rect 24508 4676 24564 4678
rect 24612 4730 24668 4732
rect 24612 4678 24614 4730
rect 24614 4678 24666 4730
rect 24666 4678 24668 4730
rect 24612 4676 24668 4678
rect 24716 4730 24772 4732
rect 24716 4678 24718 4730
rect 24718 4678 24770 4730
rect 24770 4678 24772 4730
rect 24716 4676 24772 4678
rect 24332 3836 24388 3892
rect 7036 3162 7092 3164
rect 7036 3110 7038 3162
rect 7038 3110 7090 3162
rect 7090 3110 7092 3162
rect 7036 3108 7092 3110
rect 7140 3162 7196 3164
rect 7140 3110 7142 3162
rect 7142 3110 7194 3162
rect 7194 3110 7196 3162
rect 7140 3108 7196 3110
rect 7244 3162 7300 3164
rect 7244 3110 7246 3162
rect 7246 3110 7298 3162
rect 7298 3110 7300 3162
rect 7244 3108 7300 3110
rect 12860 3162 12916 3164
rect 12860 3110 12862 3162
rect 12862 3110 12914 3162
rect 12914 3110 12916 3162
rect 12860 3108 12916 3110
rect 12964 3162 13020 3164
rect 12964 3110 12966 3162
rect 12966 3110 13018 3162
rect 13018 3110 13020 3162
rect 12964 3108 13020 3110
rect 13068 3162 13124 3164
rect 13068 3110 13070 3162
rect 13070 3110 13122 3162
rect 13122 3110 13124 3162
rect 13068 3108 13124 3110
rect 18684 3162 18740 3164
rect 18684 3110 18686 3162
rect 18686 3110 18738 3162
rect 18738 3110 18740 3162
rect 18684 3108 18740 3110
rect 18788 3162 18844 3164
rect 18788 3110 18790 3162
rect 18790 3110 18842 3162
rect 18842 3110 18844 3162
rect 18788 3108 18844 3110
rect 18892 3162 18948 3164
rect 18892 3110 18894 3162
rect 18894 3110 18946 3162
rect 18946 3110 18948 3162
rect 18892 3108 18948 3110
rect 24508 3162 24564 3164
rect 24508 3110 24510 3162
rect 24510 3110 24562 3162
rect 24562 3110 24564 3162
rect 24508 3108 24564 3110
rect 24612 3162 24668 3164
rect 24612 3110 24614 3162
rect 24614 3110 24666 3162
rect 24666 3110 24668 3162
rect 24612 3108 24668 3110
rect 24716 3162 24772 3164
rect 24716 3110 24718 3162
rect 24718 3110 24770 3162
rect 24770 3110 24772 3162
rect 24716 3108 24772 3110
rect 21532 1820 21588 1876
<< metal3 >>
rect 25200 24052 26000 24080
rect 22866 23996 22876 24052
rect 22932 23996 26000 24052
rect 25200 23968 26000 23996
rect 4114 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4398 22764
rect 9938 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10222 22764
rect 15762 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16046 22764
rect 21586 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21870 22764
rect 21298 22540 21308 22596
rect 21364 22540 22540 22596
rect 22596 22540 22606 22596
rect 10098 22316 10108 22372
rect 10164 22316 11564 22372
rect 11620 22316 11630 22372
rect 12786 22316 12796 22372
rect 12852 22316 13580 22372
rect 13636 22316 13972 22372
rect 14028 22316 14038 22372
rect 19562 22204 19572 22260
rect 19628 22204 19740 22260
rect 19796 22204 24948 22260
rect 7186 22092 7196 22148
rect 7252 22092 8428 22148
rect 8484 22092 9324 22148
rect 9380 22092 9390 22148
rect 24892 22036 24948 22204
rect 25200 22036 26000 22064
rect 24892 21980 26000 22036
rect 7026 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7310 21980
rect 12850 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13134 21980
rect 18674 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18958 21980
rect 24498 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24782 21980
rect 25200 21952 26000 21980
rect 20066 21868 20076 21924
rect 20132 21868 22036 21924
rect 17826 21644 17836 21700
rect 17892 21644 21532 21700
rect 21588 21644 21598 21700
rect 7410 21532 7420 21588
rect 7476 21532 8204 21588
rect 8260 21532 8270 21588
rect 17266 21532 17276 21588
rect 17332 21532 20860 21588
rect 20916 21532 20926 21588
rect 5506 21420 5516 21476
rect 5572 21420 7980 21476
rect 8036 21420 8046 21476
rect 11330 21420 11340 21476
rect 11396 21420 13916 21476
rect 13972 21420 13982 21476
rect 21980 21252 22036 21868
rect 21970 21196 21980 21252
rect 22036 21196 22046 21252
rect 4114 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4398 21196
rect 9938 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10222 21196
rect 15762 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16046 21196
rect 21586 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21870 21196
rect 10322 21084 10332 21140
rect 10388 21084 11340 21140
rect 11396 21084 14812 21140
rect 14868 21084 14878 21140
rect 20290 20972 20300 21028
rect 20356 20972 21084 21028
rect 21140 20972 21364 21028
rect 21420 20972 21430 21028
rect 7970 20860 7980 20916
rect 8036 20860 10332 20916
rect 10388 20860 10398 20916
rect 10882 20860 10892 20916
rect 10948 20860 12236 20916
rect 12292 20860 12302 20916
rect 14802 20860 14812 20916
rect 14868 20860 17836 20916
rect 17892 20860 17902 20916
rect 8082 20748 8092 20804
rect 8148 20748 9212 20804
rect 9268 20748 9278 20804
rect 9650 20748 9660 20804
rect 9716 20748 10556 20804
rect 10612 20748 10622 20804
rect 11666 20748 11676 20804
rect 11732 20748 12124 20804
rect 12180 20748 12190 20804
rect 14690 20748 14700 20804
rect 14756 20748 15148 20804
rect 15204 20748 17052 20804
rect 17108 20748 17118 20804
rect 18946 20748 18956 20804
rect 19012 20748 20076 20804
rect 20132 20748 20412 20804
rect 20468 20748 21868 20804
rect 21924 20748 23080 20804
rect 23136 20748 23146 20804
rect 8978 20524 8988 20580
rect 9044 20524 10444 20580
rect 10500 20524 10510 20580
rect 7026 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7310 20412
rect 12850 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13134 20412
rect 18674 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18958 20412
rect 24498 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24782 20412
rect 19170 20300 19180 20356
rect 19236 20300 20636 20356
rect 20692 20300 21644 20356
rect 21700 20300 21710 20356
rect 22642 20300 22652 20356
rect 22708 20300 22876 20356
rect 22932 20300 22942 20356
rect 4666 20188 4676 20244
rect 4732 20188 5516 20244
rect 5572 20188 6300 20244
rect 6356 20188 8764 20244
rect 8820 20188 8830 20244
rect 11452 20188 11564 20244
rect 11620 20188 11630 20244
rect 18386 20188 18396 20244
rect 18452 20188 19740 20244
rect 19796 20188 19806 20244
rect 11452 20132 11508 20188
rect 9874 20076 9884 20132
rect 9940 20076 13804 20132
rect 13860 20076 14140 20132
rect 14196 20076 15148 20132
rect 15204 20076 15214 20132
rect 20514 20076 20524 20132
rect 20580 20076 23548 20132
rect 23604 20076 23614 20132
rect 25200 20020 26000 20048
rect 9202 19964 9212 20020
rect 9268 19964 9660 20020
rect 9716 19964 9726 20020
rect 10658 19964 10668 20020
rect 10724 19964 12348 20020
rect 12404 19964 12414 20020
rect 19394 19964 19404 20020
rect 19460 19964 20188 20020
rect 20244 19964 20254 20020
rect 22876 19964 22988 20020
rect 23044 19964 23054 20020
rect 24882 19964 24892 20020
rect 24948 19964 26000 20020
rect 6178 19852 6188 19908
rect 6244 19852 11732 19908
rect 11788 19852 11798 19908
rect 22614 19852 22652 19908
rect 22708 19852 22718 19908
rect 22876 19684 22932 19964
rect 25200 19936 26000 19964
rect 22866 19628 22876 19684
rect 22932 19628 22942 19684
rect 23436 19628 23996 19684
rect 24052 19628 24062 19684
rect 4114 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4398 19628
rect 9938 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10222 19628
rect 15762 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16046 19628
rect 21586 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21870 19628
rect 23436 19572 23492 19628
rect 23426 19516 23436 19572
rect 23492 19516 23502 19572
rect 9650 19292 9660 19348
rect 9716 19292 12068 19348
rect 12124 19292 13580 19348
rect 13636 19292 13646 19348
rect 9482 19180 9492 19236
rect 9548 19180 10220 19236
rect 10276 19180 10836 19236
rect 10892 19180 10902 19236
rect 11386 19180 11396 19236
rect 11452 19180 11900 19236
rect 11956 19180 11966 19236
rect 13682 19180 13692 19236
rect 13748 19180 15484 19236
rect 15540 19180 15550 19236
rect 20626 19180 20636 19236
rect 20692 19180 21420 19236
rect 21476 19180 21486 19236
rect 21746 19180 21756 19236
rect 21812 19180 23231 19236
rect 23287 19180 23297 19236
rect 21756 19124 21812 19180
rect 8978 19068 8988 19124
rect 9044 19068 9212 19124
rect 9268 19068 11004 19124
rect 11060 19068 11070 19124
rect 19506 19068 19516 19124
rect 19572 19068 20860 19124
rect 20916 19068 21812 19124
rect 4722 18844 4732 18900
rect 4788 18844 5068 18900
rect 5124 18844 5134 18900
rect 7026 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7310 18844
rect 12850 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13134 18844
rect 18674 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18958 18844
rect 24498 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24782 18844
rect 2818 18620 2828 18676
rect 2884 18620 6748 18676
rect 6804 18620 6814 18676
rect 9986 18508 9996 18564
rect 10052 18508 11116 18564
rect 11172 18508 12348 18564
rect 12404 18508 12414 18564
rect 4274 18396 4284 18452
rect 4340 18396 5292 18452
rect 5348 18396 5358 18452
rect 12002 18396 12012 18452
rect 12068 18396 12460 18452
rect 12516 18396 12908 18452
rect 12964 18396 12974 18452
rect 18162 18396 18172 18452
rect 18228 18396 20188 18452
rect 20244 18396 20254 18452
rect 23090 18396 23100 18452
rect 23156 18396 23996 18452
rect 24052 18396 24062 18452
rect 5058 18284 5068 18340
rect 5124 18284 6728 18340
rect 6784 18284 6794 18340
rect 22026 18284 22036 18340
rect 22092 18284 22764 18340
rect 22820 18284 22830 18340
rect 8082 18172 8092 18228
rect 8148 18172 12124 18228
rect 12180 18172 12572 18228
rect 12628 18172 12638 18228
rect 22418 18060 22428 18116
rect 22484 18060 22494 18116
rect 4114 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4398 18060
rect 9938 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10222 18060
rect 15762 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16046 18060
rect 21586 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21870 18060
rect 6514 17948 6524 18004
rect 6580 17948 8148 18004
rect 7494 17836 7532 17892
rect 7588 17836 7598 17892
rect 7858 17836 7868 17892
rect 7924 17836 7934 17892
rect 7868 17668 7924 17836
rect 8092 17780 8148 17948
rect 22428 17892 22484 18060
rect 25200 18004 26000 18032
rect 22754 17948 22764 18004
rect 22820 17948 26000 18004
rect 25200 17920 26000 17948
rect 8642 17836 8652 17892
rect 8708 17836 11116 17892
rect 11172 17836 11844 17892
rect 11900 17836 11910 17892
rect 22092 17836 22484 17892
rect 8092 17724 10556 17780
rect 10612 17724 10622 17780
rect 14578 17724 14588 17780
rect 14644 17724 15148 17780
rect 15204 17724 15214 17780
rect 22092 17668 22148 17836
rect 4162 17612 4172 17668
rect 4228 17612 4676 17668
rect 4732 17612 4742 17668
rect 6290 17612 6300 17668
rect 6356 17612 8316 17668
rect 8372 17612 8382 17668
rect 8474 17612 8484 17668
rect 8540 17612 9212 17668
rect 9268 17612 9278 17668
rect 11554 17612 11564 17668
rect 11620 17612 12236 17668
rect 12292 17612 12302 17668
rect 22082 17612 22092 17668
rect 22148 17612 22158 17668
rect 4946 17500 4956 17556
rect 5012 17500 8596 17556
rect 8540 17444 8596 17500
rect 6010 17388 6020 17444
rect 6076 17388 6412 17444
rect 6468 17388 8428 17444
rect 8530 17388 8540 17444
rect 8596 17388 8606 17444
rect 8372 17332 8428 17388
rect 8764 17332 8820 17612
rect 19394 17500 19404 17556
rect 19460 17500 20076 17556
rect 20132 17500 22204 17556
rect 22260 17500 22968 17556
rect 23024 17500 23034 17556
rect 4274 17276 4284 17332
rect 4340 17276 6468 17332
rect 7410 17276 7420 17332
rect 7476 17276 8092 17332
rect 8148 17276 8158 17332
rect 8372 17276 8820 17332
rect 6412 17220 6468 17276
rect 7026 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7310 17276
rect 12850 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13134 17276
rect 18674 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18958 17276
rect 24498 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24782 17276
rect 4620 17164 5852 17220
rect 5908 17164 5918 17220
rect 6402 17164 6412 17220
rect 6468 17164 6478 17220
rect 8306 17164 8316 17220
rect 8372 17164 8652 17220
rect 8708 17164 8718 17220
rect 4620 17108 4676 17164
rect 3714 17052 3724 17108
rect 3780 17052 4620 17108
rect 4676 17052 4686 17108
rect 5058 17052 5068 17108
rect 5124 17052 8204 17108
rect 8260 17052 8270 17108
rect 8428 17052 8988 17108
rect 9044 17052 10276 17108
rect 18498 17052 18508 17108
rect 18564 17052 20188 17108
rect 20244 17052 20254 17108
rect 8428 16996 8484 17052
rect 10220 16996 10276 17052
rect 3266 16940 3276 16996
rect 3332 16940 4060 16996
rect 4116 16940 4126 16996
rect 4386 16940 4396 16996
rect 4452 16940 6300 16996
rect 6356 16940 6366 16996
rect 8306 16940 8316 16996
rect 8372 16940 8484 16996
rect 8540 16940 8876 16996
rect 8932 16940 9884 16996
rect 9940 16940 9950 16996
rect 10210 16940 10220 16996
rect 10276 16940 23100 16996
rect 23156 16940 23166 16996
rect 8540 16884 8596 16940
rect 2370 16828 2380 16884
rect 2436 16828 3388 16884
rect 3444 16828 3454 16884
rect 4946 16828 4956 16884
rect 5012 16828 5022 16884
rect 6850 16828 6860 16884
rect 6916 16828 7868 16884
rect 7924 16828 7934 16884
rect 8194 16828 8204 16884
rect 8260 16828 8596 16884
rect 8754 16828 8764 16884
rect 8820 16828 9548 16884
rect 9604 16828 9614 16884
rect 12114 16828 12124 16884
rect 12180 16828 12908 16884
rect 12964 16828 12974 16884
rect 13402 16828 13412 16884
rect 13468 16828 14252 16884
rect 14308 16828 14700 16884
rect 14756 16828 14766 16884
rect 19730 16828 19740 16884
rect 19796 16828 20412 16884
rect 20468 16828 20478 16884
rect 23650 16828 23660 16884
rect 23716 16828 25004 16884
rect 25060 16828 25070 16884
rect 4956 16772 5012 16828
rect 3602 16716 3612 16772
rect 3668 16716 5012 16772
rect 6738 16716 6748 16772
rect 6804 16716 8428 16772
rect 7522 16604 7532 16660
rect 7588 16604 7644 16660
rect 7700 16604 7710 16660
rect 8372 16604 8428 16716
rect 8484 16604 8494 16660
rect 19618 16604 19628 16660
rect 19684 16604 20076 16660
rect 20132 16604 20142 16660
rect 4114 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4398 16492
rect 9938 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10222 16492
rect 15762 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16046 16492
rect 21586 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21870 16492
rect 3042 16156 3052 16212
rect 3108 16156 3612 16212
rect 3668 16156 3678 16212
rect 4386 16156 4396 16212
rect 4452 16156 5684 16212
rect 11778 16156 11788 16212
rect 11844 16156 11854 16212
rect 2818 16044 2828 16100
rect 2884 16044 3500 16100
rect 3556 16044 4562 16100
rect 4618 16044 4628 16100
rect 5628 15988 5684 16156
rect 11788 16100 11844 16156
rect 7970 16044 7980 16100
rect 8036 16044 11452 16100
rect 11508 16044 12236 16100
rect 12292 16044 12302 16100
rect 12506 16044 12516 16100
rect 12572 16044 14364 16100
rect 14420 16044 14430 16100
rect 19282 16044 19292 16100
rect 19348 16044 20636 16100
rect 20692 16044 21084 16100
rect 21140 16044 21150 16100
rect 21746 16044 21756 16100
rect 21812 16044 22428 16100
rect 22484 16044 22783 16100
rect 22839 16044 22849 16100
rect 25200 15988 26000 16016
rect 5618 15932 5628 15988
rect 5684 15932 6636 15988
rect 6692 15932 7644 15988
rect 7700 15932 7710 15988
rect 11722 15932 11732 15988
rect 11788 15932 19180 15988
rect 19236 15932 19246 15988
rect 24266 15932 24276 15988
rect 24332 15932 26000 15988
rect 25200 15904 26000 15932
rect 4274 15820 4284 15876
rect 4340 15820 6300 15876
rect 6356 15820 9660 15876
rect 9716 15820 10556 15876
rect 10612 15820 10622 15876
rect 21970 15820 21980 15876
rect 22036 15820 22764 15876
rect 22820 15820 22830 15876
rect 3154 15708 3164 15764
rect 3220 15708 3836 15764
rect 3892 15708 3902 15764
rect 7026 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7310 15708
rect 12850 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13134 15708
rect 18674 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18958 15708
rect 24498 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24782 15708
rect 8866 15484 8876 15540
rect 8932 15484 10220 15540
rect 10276 15484 10286 15540
rect 12338 15484 12348 15540
rect 12404 15484 13580 15540
rect 13636 15484 13646 15540
rect 3938 15372 3948 15428
rect 4004 15372 4508 15428
rect 4564 15372 4574 15428
rect 5730 15372 5740 15428
rect 5796 15372 7532 15428
rect 7588 15372 7598 15428
rect 20178 15372 20188 15428
rect 20244 15372 21252 15428
rect 21308 15372 21318 15428
rect 7410 15260 7420 15316
rect 7476 15260 7980 15316
rect 8036 15260 8046 15316
rect 9762 15260 9772 15316
rect 9828 15260 10332 15316
rect 10388 15260 10398 15316
rect 10668 15260 10780 15316
rect 10836 15260 11228 15316
rect 11284 15260 11294 15316
rect 19954 15260 19964 15316
rect 20020 15260 20860 15316
rect 20916 15260 21756 15316
rect 21812 15260 21822 15316
rect 22530 15260 22540 15316
rect 22596 15260 23548 15316
rect 23604 15260 23614 15316
rect 10668 15204 10724 15260
rect 7244 15148 7254 15204
rect 7310 15148 10052 15204
rect 10108 15148 10724 15204
rect 10882 15148 10892 15204
rect 10948 15148 12012 15204
rect 12068 15148 12078 15204
rect 18508 15148 20076 15204
rect 20132 15148 20142 15204
rect 22642 15148 22652 15204
rect 22708 15148 22988 15204
rect 23044 15148 23054 15204
rect 23202 15148 23212 15204
rect 23268 15148 24108 15204
rect 24164 15148 24174 15204
rect 4722 15036 4732 15092
rect 4788 15036 6412 15092
rect 6468 15036 6860 15092
rect 6916 15036 6926 15092
rect 7382 15036 7420 15092
rect 7476 15036 7486 15092
rect 15810 15036 15820 15092
rect 15876 15036 17052 15092
rect 17108 15036 17118 15092
rect 18508 14980 18564 15148
rect 18498 14924 18508 14980
rect 18564 14924 18574 14980
rect 4114 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4398 14924
rect 9938 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10222 14924
rect 15762 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16046 14924
rect 21586 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21870 14924
rect 20346 14700 20356 14756
rect 20412 14700 20524 14756
rect 20580 14700 21420 14756
rect 21476 14700 21486 14756
rect 5786 14476 5796 14532
rect 5852 14476 6524 14532
rect 6580 14476 6590 14532
rect 7858 14476 7868 14532
rect 7924 14476 8260 14532
rect 8316 14476 8326 14532
rect 13010 14476 13020 14532
rect 13076 14476 14382 14532
rect 14438 14476 14448 14532
rect 8754 14364 8764 14420
rect 8820 14364 11116 14420
rect 11172 14364 11182 14420
rect 13458 14364 13468 14420
rect 13524 14364 13804 14420
rect 13860 14364 14924 14420
rect 14980 14364 14990 14420
rect 3490 14252 3500 14308
rect 3556 14252 4900 14308
rect 4956 14252 9100 14308
rect 9156 14252 9166 14308
rect 7026 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7310 14140
rect 12850 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13134 14140
rect 18674 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18958 14140
rect 24498 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24782 14140
rect 25200 13972 26000 14000
rect 23594 13916 23604 13972
rect 23660 13916 23772 13972
rect 23828 13916 26000 13972
rect 25200 13888 26000 13916
rect 4834 13804 4844 13860
rect 4900 13804 6972 13860
rect 7028 13804 7038 13860
rect 7522 13804 7532 13860
rect 7588 13804 7980 13860
rect 8036 13804 8316 13860
rect 8372 13804 8382 13860
rect 2818 13692 2828 13748
rect 2884 13692 4508 13748
rect 4564 13692 4574 13748
rect 6514 13692 6524 13748
rect 6580 13692 7756 13748
rect 7812 13692 9212 13748
rect 9268 13692 11396 13748
rect 11452 13692 11462 13748
rect 20850 13692 20860 13748
rect 20916 13692 21308 13748
rect 21364 13692 23100 13748
rect 23156 13692 23166 13748
rect 4610 13580 4620 13636
rect 4676 13580 10948 13636
rect 11004 13580 11788 13636
rect 11844 13580 11854 13636
rect 20626 13580 20636 13636
rect 20692 13580 21644 13636
rect 21700 13580 22204 13636
rect 22260 13580 22270 13636
rect 1586 13468 1596 13524
rect 1652 13468 4900 13524
rect 4956 13468 6524 13524
rect 6580 13468 6590 13524
rect 7634 13468 7644 13524
rect 7700 13468 8540 13524
rect 8596 13468 8606 13524
rect 9772 13468 10108 13524
rect 10164 13468 10174 13524
rect 19404 13468 21420 13524
rect 21476 13468 21486 13524
rect 9772 13412 9828 13468
rect 19404 13412 19460 13468
rect 6066 13356 6076 13412
rect 6132 13356 9828 13412
rect 19394 13356 19404 13412
rect 19460 13356 19470 13412
rect 4114 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4398 13356
rect 9938 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10222 13356
rect 15762 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16046 13356
rect 21586 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21870 13356
rect 6738 13244 6748 13300
rect 6804 13244 8126 13300
rect 8182 13244 8192 13300
rect 16706 13244 16716 13300
rect 16772 13244 17724 13300
rect 17780 13244 17790 13300
rect 16716 13188 16772 13244
rect 5740 13132 6860 13188
rect 6916 13132 7420 13188
rect 7476 13132 7486 13188
rect 13346 13132 13356 13188
rect 13412 13132 16772 13188
rect 3714 13020 3724 13076
rect 3780 13020 4284 13076
rect 4340 13020 4350 13076
rect 5740 12964 5796 13132
rect 7074 13020 7084 13076
rect 7140 13020 7644 13076
rect 7700 13020 7710 13076
rect 14578 13020 14588 13076
rect 14644 13020 15372 13076
rect 15428 13020 15438 13076
rect 2370 12908 2380 12964
rect 2436 12908 3836 12964
rect 3892 12908 3902 12964
rect 5058 12908 5068 12964
rect 5124 12908 5740 12964
rect 5796 12908 5806 12964
rect 5954 12908 5964 12964
rect 6020 12908 7252 12964
rect 7308 12908 7318 12964
rect 23426 12908 23436 12964
rect 23492 12908 23996 12964
rect 24052 12908 24062 12964
rect 7410 12796 7420 12852
rect 7476 12796 7532 12852
rect 7588 12796 7598 12852
rect 14820 12796 14830 12852
rect 14886 12796 15596 12852
rect 15652 12796 15662 12852
rect 21074 12796 21084 12852
rect 21140 12796 22559 12852
rect 22615 12796 22625 12852
rect 4274 12684 4284 12740
rect 4340 12684 5964 12740
rect 6020 12684 6030 12740
rect 7026 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7310 12572
rect 12850 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13134 12572
rect 18674 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18958 12572
rect 24498 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24782 12572
rect 5170 12348 5180 12404
rect 5236 12348 9996 12404
rect 10052 12348 10062 12404
rect 10658 12348 10668 12404
rect 10724 12348 11116 12404
rect 11172 12348 13356 12404
rect 13412 12348 13422 12404
rect 15922 12348 15932 12404
rect 15988 12348 17276 12404
rect 17332 12348 17342 12404
rect 3266 12236 3276 12292
rect 3332 12236 3836 12292
rect 3892 12236 4732 12292
rect 4788 12236 5068 12292
rect 5124 12236 5134 12292
rect 6178 12236 6188 12292
rect 6244 12236 6636 12292
rect 6692 12236 8204 12292
rect 8260 12236 8270 12292
rect 10490 12236 10500 12292
rect 10556 12236 11900 12292
rect 11956 12236 11966 12292
rect 23202 12236 23212 12292
rect 23268 12236 24052 12292
rect 24108 12236 24118 12292
rect 4162 12124 4172 12180
rect 4228 12124 4956 12180
rect 5012 12124 5404 12180
rect 5460 12124 6782 12180
rect 6838 12124 6848 12180
rect 7186 12124 7196 12180
rect 7252 12124 8316 12180
rect 8372 12124 8382 12180
rect 8548 12124 8558 12180
rect 8614 12124 9660 12180
rect 9716 12124 9726 12180
rect 10994 12124 11004 12180
rect 11060 12124 15036 12180
rect 15092 12124 15102 12180
rect 22978 12124 22988 12180
rect 23044 12124 23884 12180
rect 23940 12124 23950 12180
rect 7410 12012 7420 12068
rect 7476 12012 8092 12068
rect 8148 12012 8158 12068
rect 10322 12012 10332 12068
rect 10388 12012 12012 12068
rect 12068 12012 12078 12068
rect 20132 12012 22092 12068
rect 22148 12012 22158 12068
rect 13906 11900 13916 11956
rect 13972 11900 14700 11956
rect 14756 11900 14766 11956
rect 20132 11844 20188 12012
rect 25200 11956 26000 11984
rect 24266 11900 24276 11956
rect 24332 11900 26000 11956
rect 25200 11872 26000 11900
rect 6066 11788 6076 11844
rect 6132 11788 6860 11844
rect 6916 11788 6926 11844
rect 19842 11788 19852 11844
rect 19908 11788 20188 11844
rect 4114 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4398 11788
rect 9938 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10222 11788
rect 15762 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16046 11788
rect 21586 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21870 11788
rect 11236 11676 11246 11732
rect 11302 11676 12684 11732
rect 12740 11676 12750 11732
rect 22866 11564 22876 11620
rect 22932 11564 23660 11620
rect 23716 11564 23726 11620
rect 3938 11452 3948 11508
rect 4004 11452 5796 11508
rect 5852 11452 6412 11508
rect 6468 11452 6478 11508
rect 21746 11452 21756 11508
rect 21812 11452 22652 11508
rect 22708 11452 23324 11508
rect 23380 11452 23390 11508
rect 5058 11340 5068 11396
rect 5124 11340 5628 11396
rect 5684 11340 5694 11396
rect 9650 11340 9660 11396
rect 9716 11340 10892 11396
rect 10948 11340 10958 11396
rect 4610 11228 4620 11284
rect 4676 11228 6076 11284
rect 6132 11228 6142 11284
rect 7970 11228 7980 11284
rect 8036 11228 8428 11284
rect 8484 11228 8494 11284
rect 15250 11228 15260 11284
rect 15316 11228 16044 11284
rect 16100 11228 16110 11284
rect 12786 11116 12796 11172
rect 12852 11116 13636 11172
rect 13692 11116 13702 11172
rect 7410 11004 7420 11060
rect 7476 11004 7486 11060
rect 7026 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7310 11004
rect 7420 10836 7476 11004
rect 12850 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13134 11004
rect 18674 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18958 11004
rect 24498 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24782 11004
rect 7298 10780 7308 10836
rect 7364 10780 7476 10836
rect 7644 10780 7756 10836
rect 7812 10780 7822 10836
rect 16258 10780 16268 10836
rect 16324 10780 17948 10836
rect 18004 10780 18014 10836
rect 5282 10556 5292 10612
rect 5348 10556 6412 10612
rect 6468 10556 6478 10612
rect 6962 10444 6972 10500
rect 7028 10444 7420 10500
rect 7476 10444 7486 10500
rect 7644 10388 7700 10780
rect 14130 10556 14140 10612
rect 14196 10556 15260 10612
rect 15316 10556 15326 10612
rect 3602 10332 3612 10388
rect 3668 10332 7700 10388
rect 7644 10276 7700 10332
rect 7634 10220 7644 10276
rect 7700 10220 7710 10276
rect 4114 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4398 10220
rect 9938 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10222 10220
rect 15762 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16046 10220
rect 21586 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21870 10220
rect 22250 10108 22260 10164
rect 22316 10108 23772 10164
rect 23828 10108 23838 10164
rect 6682 9996 6692 10052
rect 6748 9996 7308 10052
rect 7364 9996 7532 10052
rect 7588 9996 7598 10052
rect 23772 9940 23828 10108
rect 25200 9940 26000 9968
rect 7410 9884 7420 9940
rect 7476 9884 9884 9940
rect 9940 9884 9950 9940
rect 12338 9884 12348 9940
rect 12404 9884 13636 9940
rect 13692 9884 13702 9940
rect 21410 9884 21420 9940
rect 21476 9884 21980 9940
rect 22036 9884 22046 9940
rect 23772 9884 26000 9940
rect 25200 9856 26000 9884
rect 8642 9772 8652 9828
rect 8708 9772 10220 9828
rect 10276 9772 10286 9828
rect 14130 9772 14140 9828
rect 14196 9772 15484 9828
rect 15540 9772 16492 9828
rect 16548 9772 16558 9828
rect 19170 9548 19180 9604
rect 19236 9548 21196 9604
rect 21252 9548 21262 9604
rect 23333 9548 23343 9604
rect 23399 9548 23548 9604
rect 23604 9548 23884 9604
rect 23940 9548 23950 9604
rect 7026 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7310 9436
rect 12850 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13134 9436
rect 18674 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18958 9436
rect 24498 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24782 9436
rect 16594 9212 16604 9268
rect 16660 9212 18396 9268
rect 18452 9212 18462 9268
rect 12898 9100 12908 9156
rect 12964 9100 13244 9156
rect 13300 9100 13804 9156
rect 13860 9100 13870 9156
rect 7634 8876 7644 8932
rect 7700 8876 13748 8932
rect 13804 8876 13814 8932
rect 7746 8764 7756 8820
rect 7812 8764 10556 8820
rect 10612 8764 10622 8820
rect 4114 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4398 8652
rect 9938 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10222 8652
rect 15762 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16046 8652
rect 21586 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21870 8652
rect 8082 8540 8092 8596
rect 8148 8540 8158 8596
rect 8092 8372 8148 8540
rect 5170 8316 5180 8372
rect 5236 8316 6860 8372
rect 6916 8316 7532 8372
rect 7588 8316 9772 8372
rect 9828 8316 9838 8372
rect 11116 8316 12348 8372
rect 12404 8316 13468 8372
rect 13524 8316 13534 8372
rect 14354 8316 14364 8372
rect 14420 8316 14924 8372
rect 14980 8316 15708 8372
rect 15764 8316 15774 8372
rect 23090 8316 23100 8372
rect 23156 8316 24892 8372
rect 24948 8316 24958 8372
rect 11116 8036 11172 8316
rect 19954 8204 19964 8260
rect 20020 8204 22092 8260
rect 22148 8204 22158 8260
rect 11106 7980 11116 8036
rect 11172 7980 11676 8036
rect 11732 7980 11742 8036
rect 25200 7924 26000 7952
rect 24892 7868 26000 7924
rect 7026 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7310 7868
rect 12850 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13134 7868
rect 18674 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18958 7868
rect 24498 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24782 7868
rect 24892 7700 24948 7868
rect 25200 7840 26000 7868
rect 16146 7644 16156 7700
rect 16212 7644 17612 7700
rect 17668 7644 17678 7700
rect 21634 7644 21644 7700
rect 21700 7644 23100 7700
rect 23156 7644 23343 7700
rect 23399 7644 23409 7700
rect 23762 7644 23772 7700
rect 23828 7644 24948 7700
rect 9538 7532 9548 7588
rect 9604 7532 13636 7588
rect 13692 7532 13702 7588
rect 21970 7532 21980 7588
rect 22036 7532 22428 7588
rect 22484 7532 22494 7588
rect 18722 7420 18732 7476
rect 18788 7420 19852 7476
rect 19908 7420 19918 7476
rect 7858 7308 7868 7364
rect 7924 7308 11284 7364
rect 11340 7308 11350 7364
rect 4114 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4398 7084
rect 9938 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10222 7084
rect 15762 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16046 7084
rect 21586 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21870 7084
rect 23202 6860 23212 6916
rect 23268 6860 23884 6916
rect 23940 6860 23950 6916
rect 14690 6748 14700 6804
rect 14756 6748 15820 6804
rect 15876 6748 15886 6804
rect 10210 6636 10220 6692
rect 10276 6636 11844 6692
rect 11900 6636 11910 6692
rect 12580 6524 12590 6580
rect 12646 6524 13356 6580
rect 13412 6524 13422 6580
rect 16706 6412 16716 6468
rect 16772 6412 18284 6468
rect 18340 6412 18956 6468
rect 19012 6412 19022 6468
rect 21970 6412 21980 6468
rect 22036 6412 22876 6468
rect 22932 6412 22942 6468
rect 7026 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7310 6300
rect 12850 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13134 6300
rect 18674 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18958 6300
rect 24498 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24782 6300
rect 22642 6188 22652 6244
rect 22708 6188 24332 6244
rect 24388 6188 24398 6244
rect 18741 6076 18751 6132
rect 18807 6076 20300 6132
rect 20356 6076 20804 6132
rect 20860 6076 20870 6132
rect 12674 5964 12684 6020
rect 12740 5964 13244 6020
rect 13300 5964 13310 6020
rect 19618 5964 19628 6020
rect 19684 5964 22092 6020
rect 22148 5964 22559 6020
rect 22615 5964 22625 6020
rect 25200 5908 26000 5936
rect 11218 5852 11228 5908
rect 11284 5852 11770 5908
rect 11826 5852 11836 5908
rect 20962 5852 20972 5908
rect 21028 5852 21420 5908
rect 21476 5852 22204 5908
rect 22260 5852 22270 5908
rect 23426 5852 23436 5908
rect 23492 5852 23996 5908
rect 24052 5852 24062 5908
rect 24210 5852 24220 5908
rect 24276 5852 26000 5908
rect 25200 5824 26000 5852
rect 20178 5740 20188 5796
rect 20244 5740 21196 5796
rect 21252 5740 21756 5796
rect 21812 5740 21822 5796
rect 20290 5628 20300 5684
rect 20356 5628 21084 5684
rect 21140 5628 21980 5684
rect 22036 5628 22046 5684
rect 4114 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4398 5516
rect 9938 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10222 5516
rect 15762 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16046 5516
rect 21586 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21870 5516
rect 22418 5292 22428 5348
rect 22484 5292 23996 5348
rect 24052 5292 24062 5348
rect 20962 5180 20972 5236
rect 21028 5180 21588 5236
rect 23314 5180 23324 5236
rect 23380 5180 25004 5236
rect 25060 5180 25070 5236
rect 21532 5124 21588 5180
rect 18274 5068 18284 5124
rect 18340 5068 21308 5124
rect 21364 5068 21374 5124
rect 21522 5068 21532 5124
rect 21588 5068 21598 5124
rect 22530 5068 22540 5124
rect 22596 5068 23660 5124
rect 23716 5068 23726 5124
rect 7026 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7310 4732
rect 12850 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13134 4732
rect 18674 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18958 4732
rect 24498 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24782 4732
rect 19394 4508 19404 4564
rect 19460 4508 20188 4564
rect 20132 4340 20188 4508
rect 20132 4284 22092 4340
rect 22148 4284 22158 4340
rect 23182 3948 23192 4004
rect 23248 3948 23996 4004
rect 24052 3948 24062 4004
rect 4114 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4398 3948
rect 9938 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10222 3948
rect 15762 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16046 3948
rect 21586 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21870 3948
rect 25200 3892 26000 3920
rect 24322 3836 24332 3892
rect 24388 3836 26000 3892
rect 25200 3808 26000 3836
rect 7026 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7310 3164
rect 12850 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13134 3164
rect 18674 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18958 3164
rect 24498 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24782 3164
rect 25200 1876 26000 1904
rect 21522 1820 21532 1876
rect 21588 1820 26000 1876
rect 25200 1792 26000 1820
<< via3 >>
rect 4124 22708 4180 22764
rect 4228 22708 4284 22764
rect 4332 22708 4388 22764
rect 9948 22708 10004 22764
rect 10052 22708 10108 22764
rect 10156 22708 10212 22764
rect 15772 22708 15828 22764
rect 15876 22708 15932 22764
rect 15980 22708 16036 22764
rect 21596 22708 21652 22764
rect 21700 22708 21756 22764
rect 21804 22708 21860 22764
rect 7036 21924 7092 21980
rect 7140 21924 7196 21980
rect 7244 21924 7300 21980
rect 12860 21924 12916 21980
rect 12964 21924 13020 21980
rect 13068 21924 13124 21980
rect 18684 21924 18740 21980
rect 18788 21924 18844 21980
rect 18892 21924 18948 21980
rect 24508 21924 24564 21980
rect 24612 21924 24668 21980
rect 24716 21924 24772 21980
rect 4124 21140 4180 21196
rect 4228 21140 4284 21196
rect 4332 21140 4388 21196
rect 9948 21140 10004 21196
rect 10052 21140 10108 21196
rect 10156 21140 10212 21196
rect 15772 21140 15828 21196
rect 15876 21140 15932 21196
rect 15980 21140 16036 21196
rect 21596 21140 21652 21196
rect 21700 21140 21756 21196
rect 21804 21140 21860 21196
rect 7036 20356 7092 20412
rect 7140 20356 7196 20412
rect 7244 20356 7300 20412
rect 12860 20356 12916 20412
rect 12964 20356 13020 20412
rect 13068 20356 13124 20412
rect 18684 20356 18740 20412
rect 18788 20356 18844 20412
rect 18892 20356 18948 20412
rect 24508 20356 24564 20412
rect 24612 20356 24668 20412
rect 24716 20356 24772 20412
rect 22652 20300 22708 20356
rect 22652 19852 22708 19908
rect 4124 19572 4180 19628
rect 4228 19572 4284 19628
rect 4332 19572 4388 19628
rect 9948 19572 10004 19628
rect 10052 19572 10108 19628
rect 10156 19572 10212 19628
rect 15772 19572 15828 19628
rect 15876 19572 15932 19628
rect 15980 19572 16036 19628
rect 21596 19572 21652 19628
rect 21700 19572 21756 19628
rect 21804 19572 21860 19628
rect 7036 18788 7092 18844
rect 7140 18788 7196 18844
rect 7244 18788 7300 18844
rect 12860 18788 12916 18844
rect 12964 18788 13020 18844
rect 13068 18788 13124 18844
rect 18684 18788 18740 18844
rect 18788 18788 18844 18844
rect 18892 18788 18948 18844
rect 24508 18788 24564 18844
rect 24612 18788 24668 18844
rect 24716 18788 24772 18844
rect 6748 18620 6804 18676
rect 4124 18004 4180 18060
rect 4228 18004 4284 18060
rect 4332 18004 4388 18060
rect 9948 18004 10004 18060
rect 10052 18004 10108 18060
rect 10156 18004 10212 18060
rect 15772 18004 15828 18060
rect 15876 18004 15932 18060
rect 15980 18004 16036 18060
rect 21596 18004 21652 18060
rect 21700 18004 21756 18060
rect 21804 18004 21860 18060
rect 7532 17836 7588 17892
rect 7420 17276 7476 17332
rect 7036 17220 7092 17276
rect 7140 17220 7196 17276
rect 7244 17220 7300 17276
rect 12860 17220 12916 17276
rect 12964 17220 13020 17276
rect 13068 17220 13124 17276
rect 18684 17220 18740 17276
rect 18788 17220 18844 17276
rect 18892 17220 18948 17276
rect 24508 17220 24564 17276
rect 24612 17220 24668 17276
rect 24716 17220 24772 17276
rect 6748 16716 6804 16772
rect 7532 16604 7588 16660
rect 4124 16436 4180 16492
rect 4228 16436 4284 16492
rect 4332 16436 4388 16492
rect 9948 16436 10004 16492
rect 10052 16436 10108 16492
rect 10156 16436 10212 16492
rect 15772 16436 15828 16492
rect 15876 16436 15932 16492
rect 15980 16436 16036 16492
rect 21596 16436 21652 16492
rect 21700 16436 21756 16492
rect 21804 16436 21860 16492
rect 7036 15652 7092 15708
rect 7140 15652 7196 15708
rect 7244 15652 7300 15708
rect 12860 15652 12916 15708
rect 12964 15652 13020 15708
rect 13068 15652 13124 15708
rect 18684 15652 18740 15708
rect 18788 15652 18844 15708
rect 18892 15652 18948 15708
rect 24508 15652 24564 15708
rect 24612 15652 24668 15708
rect 24716 15652 24772 15708
rect 7420 15036 7476 15092
rect 4124 14868 4180 14924
rect 4228 14868 4284 14924
rect 4332 14868 4388 14924
rect 9948 14868 10004 14924
rect 10052 14868 10108 14924
rect 10156 14868 10212 14924
rect 15772 14868 15828 14924
rect 15876 14868 15932 14924
rect 15980 14868 16036 14924
rect 21596 14868 21652 14924
rect 21700 14868 21756 14924
rect 21804 14868 21860 14924
rect 7036 14084 7092 14140
rect 7140 14084 7196 14140
rect 7244 14084 7300 14140
rect 12860 14084 12916 14140
rect 12964 14084 13020 14140
rect 13068 14084 13124 14140
rect 18684 14084 18740 14140
rect 18788 14084 18844 14140
rect 18892 14084 18948 14140
rect 24508 14084 24564 14140
rect 24612 14084 24668 14140
rect 24716 14084 24772 14140
rect 4124 13300 4180 13356
rect 4228 13300 4284 13356
rect 4332 13300 4388 13356
rect 9948 13300 10004 13356
rect 10052 13300 10108 13356
rect 10156 13300 10212 13356
rect 15772 13300 15828 13356
rect 15876 13300 15932 13356
rect 15980 13300 16036 13356
rect 21596 13300 21652 13356
rect 21700 13300 21756 13356
rect 21804 13300 21860 13356
rect 7420 12796 7476 12852
rect 7036 12516 7092 12572
rect 7140 12516 7196 12572
rect 7244 12516 7300 12572
rect 12860 12516 12916 12572
rect 12964 12516 13020 12572
rect 13068 12516 13124 12572
rect 18684 12516 18740 12572
rect 18788 12516 18844 12572
rect 18892 12516 18948 12572
rect 24508 12516 24564 12572
rect 24612 12516 24668 12572
rect 24716 12516 24772 12572
rect 4124 11732 4180 11788
rect 4228 11732 4284 11788
rect 4332 11732 4388 11788
rect 9948 11732 10004 11788
rect 10052 11732 10108 11788
rect 10156 11732 10212 11788
rect 15772 11732 15828 11788
rect 15876 11732 15932 11788
rect 15980 11732 16036 11788
rect 21596 11732 21652 11788
rect 21700 11732 21756 11788
rect 21804 11732 21860 11788
rect 7036 10948 7092 11004
rect 7140 10948 7196 11004
rect 7244 10948 7300 11004
rect 12860 10948 12916 11004
rect 12964 10948 13020 11004
rect 13068 10948 13124 11004
rect 18684 10948 18740 11004
rect 18788 10948 18844 11004
rect 18892 10948 18948 11004
rect 24508 10948 24564 11004
rect 24612 10948 24668 11004
rect 24716 10948 24772 11004
rect 7420 10444 7476 10500
rect 4124 10164 4180 10220
rect 4228 10164 4284 10220
rect 4332 10164 4388 10220
rect 9948 10164 10004 10220
rect 10052 10164 10108 10220
rect 10156 10164 10212 10220
rect 15772 10164 15828 10220
rect 15876 10164 15932 10220
rect 15980 10164 16036 10220
rect 21596 10164 21652 10220
rect 21700 10164 21756 10220
rect 21804 10164 21860 10220
rect 7036 9380 7092 9436
rect 7140 9380 7196 9436
rect 7244 9380 7300 9436
rect 12860 9380 12916 9436
rect 12964 9380 13020 9436
rect 13068 9380 13124 9436
rect 18684 9380 18740 9436
rect 18788 9380 18844 9436
rect 18892 9380 18948 9436
rect 24508 9380 24564 9436
rect 24612 9380 24668 9436
rect 24716 9380 24772 9436
rect 4124 8596 4180 8652
rect 4228 8596 4284 8652
rect 4332 8596 4388 8652
rect 9948 8596 10004 8652
rect 10052 8596 10108 8652
rect 10156 8596 10212 8652
rect 15772 8596 15828 8652
rect 15876 8596 15932 8652
rect 15980 8596 16036 8652
rect 21596 8596 21652 8652
rect 21700 8596 21756 8652
rect 21804 8596 21860 8652
rect 7036 7812 7092 7868
rect 7140 7812 7196 7868
rect 7244 7812 7300 7868
rect 12860 7812 12916 7868
rect 12964 7812 13020 7868
rect 13068 7812 13124 7868
rect 18684 7812 18740 7868
rect 18788 7812 18844 7868
rect 18892 7812 18948 7868
rect 24508 7812 24564 7868
rect 24612 7812 24668 7868
rect 24716 7812 24772 7868
rect 4124 7028 4180 7084
rect 4228 7028 4284 7084
rect 4332 7028 4388 7084
rect 9948 7028 10004 7084
rect 10052 7028 10108 7084
rect 10156 7028 10212 7084
rect 15772 7028 15828 7084
rect 15876 7028 15932 7084
rect 15980 7028 16036 7084
rect 21596 7028 21652 7084
rect 21700 7028 21756 7084
rect 21804 7028 21860 7084
rect 7036 6244 7092 6300
rect 7140 6244 7196 6300
rect 7244 6244 7300 6300
rect 12860 6244 12916 6300
rect 12964 6244 13020 6300
rect 13068 6244 13124 6300
rect 18684 6244 18740 6300
rect 18788 6244 18844 6300
rect 18892 6244 18948 6300
rect 24508 6244 24564 6300
rect 24612 6244 24668 6300
rect 24716 6244 24772 6300
rect 4124 5460 4180 5516
rect 4228 5460 4284 5516
rect 4332 5460 4388 5516
rect 9948 5460 10004 5516
rect 10052 5460 10108 5516
rect 10156 5460 10212 5516
rect 15772 5460 15828 5516
rect 15876 5460 15932 5516
rect 15980 5460 16036 5516
rect 21596 5460 21652 5516
rect 21700 5460 21756 5516
rect 21804 5460 21860 5516
rect 7036 4676 7092 4732
rect 7140 4676 7196 4732
rect 7244 4676 7300 4732
rect 12860 4676 12916 4732
rect 12964 4676 13020 4732
rect 13068 4676 13124 4732
rect 18684 4676 18740 4732
rect 18788 4676 18844 4732
rect 18892 4676 18948 4732
rect 24508 4676 24564 4732
rect 24612 4676 24668 4732
rect 24716 4676 24772 4732
rect 4124 3892 4180 3948
rect 4228 3892 4284 3948
rect 4332 3892 4388 3948
rect 9948 3892 10004 3948
rect 10052 3892 10108 3948
rect 10156 3892 10212 3948
rect 15772 3892 15828 3948
rect 15876 3892 15932 3948
rect 15980 3892 16036 3948
rect 21596 3892 21652 3948
rect 21700 3892 21756 3948
rect 21804 3892 21860 3948
rect 7036 3108 7092 3164
rect 7140 3108 7196 3164
rect 7244 3108 7300 3164
rect 12860 3108 12916 3164
rect 12964 3108 13020 3164
rect 13068 3108 13124 3164
rect 18684 3108 18740 3164
rect 18788 3108 18844 3164
rect 18892 3108 18948 3164
rect 24508 3108 24564 3164
rect 24612 3108 24668 3164
rect 24716 3108 24772 3164
<< metal4 >>
rect 4096 22764 4416 22796
rect 4096 22708 4124 22764
rect 4180 22708 4228 22764
rect 4284 22708 4332 22764
rect 4388 22708 4416 22764
rect 4096 21196 4416 22708
rect 4096 21140 4124 21196
rect 4180 21140 4228 21196
rect 4284 21140 4332 21196
rect 4388 21140 4416 21196
rect 4096 19628 4416 21140
rect 4096 19572 4124 19628
rect 4180 19572 4228 19628
rect 4284 19572 4332 19628
rect 4388 19572 4416 19628
rect 4096 18060 4416 19572
rect 7008 21980 7328 22796
rect 7008 21924 7036 21980
rect 7092 21924 7140 21980
rect 7196 21924 7244 21980
rect 7300 21924 7328 21980
rect 7008 20412 7328 21924
rect 7008 20356 7036 20412
rect 7092 20356 7140 20412
rect 7196 20356 7244 20412
rect 7300 20356 7328 20412
rect 7008 18844 7328 20356
rect 7008 18788 7036 18844
rect 7092 18788 7140 18844
rect 7196 18788 7244 18844
rect 7300 18788 7328 18844
rect 4096 18004 4124 18060
rect 4180 18004 4228 18060
rect 4284 18004 4332 18060
rect 4388 18004 4416 18060
rect 4096 16492 4416 18004
rect 6748 18676 6804 18686
rect 6748 16772 6804 18620
rect 6748 16706 6804 16716
rect 7008 17276 7328 18788
rect 9920 22764 10240 22796
rect 9920 22708 9948 22764
rect 10004 22708 10052 22764
rect 10108 22708 10156 22764
rect 10212 22708 10240 22764
rect 9920 21196 10240 22708
rect 9920 21140 9948 21196
rect 10004 21140 10052 21196
rect 10108 21140 10156 21196
rect 10212 21140 10240 21196
rect 9920 19628 10240 21140
rect 9920 19572 9948 19628
rect 10004 19572 10052 19628
rect 10108 19572 10156 19628
rect 10212 19572 10240 19628
rect 9920 18060 10240 19572
rect 9920 18004 9948 18060
rect 10004 18004 10052 18060
rect 10108 18004 10156 18060
rect 10212 18004 10240 18060
rect 7532 17892 7588 17902
rect 7008 17220 7036 17276
rect 7092 17220 7140 17276
rect 7196 17220 7244 17276
rect 7300 17220 7328 17276
rect 4096 16436 4124 16492
rect 4180 16436 4228 16492
rect 4284 16436 4332 16492
rect 4388 16436 4416 16492
rect 4096 14924 4416 16436
rect 4096 14868 4124 14924
rect 4180 14868 4228 14924
rect 4284 14868 4332 14924
rect 4388 14868 4416 14924
rect 4096 13356 4416 14868
rect 4096 13300 4124 13356
rect 4180 13300 4228 13356
rect 4284 13300 4332 13356
rect 4388 13300 4416 13356
rect 4096 11788 4416 13300
rect 4096 11732 4124 11788
rect 4180 11732 4228 11788
rect 4284 11732 4332 11788
rect 4388 11732 4416 11788
rect 4096 10220 4416 11732
rect 4096 10164 4124 10220
rect 4180 10164 4228 10220
rect 4284 10164 4332 10220
rect 4388 10164 4416 10220
rect 4096 8652 4416 10164
rect 4096 8596 4124 8652
rect 4180 8596 4228 8652
rect 4284 8596 4332 8652
rect 4388 8596 4416 8652
rect 4096 7084 4416 8596
rect 4096 7028 4124 7084
rect 4180 7028 4228 7084
rect 4284 7028 4332 7084
rect 4388 7028 4416 7084
rect 4096 5516 4416 7028
rect 4096 5460 4124 5516
rect 4180 5460 4228 5516
rect 4284 5460 4332 5516
rect 4388 5460 4416 5516
rect 4096 3948 4416 5460
rect 4096 3892 4124 3948
rect 4180 3892 4228 3948
rect 4284 3892 4332 3948
rect 4388 3892 4416 3948
rect 4096 3076 4416 3892
rect 7008 15708 7328 17220
rect 7008 15652 7036 15708
rect 7092 15652 7140 15708
rect 7196 15652 7244 15708
rect 7300 15652 7328 15708
rect 7008 14140 7328 15652
rect 7420 17332 7476 17342
rect 7420 15092 7476 17276
rect 7532 16660 7588 17836
rect 7532 16594 7588 16604
rect 7420 15026 7476 15036
rect 9920 16492 10240 18004
rect 9920 16436 9948 16492
rect 10004 16436 10052 16492
rect 10108 16436 10156 16492
rect 10212 16436 10240 16492
rect 7008 14084 7036 14140
rect 7092 14084 7140 14140
rect 7196 14084 7244 14140
rect 7300 14084 7328 14140
rect 7008 12572 7328 14084
rect 9920 14924 10240 16436
rect 9920 14868 9948 14924
rect 10004 14868 10052 14924
rect 10108 14868 10156 14924
rect 10212 14868 10240 14924
rect 9920 13356 10240 14868
rect 9920 13300 9948 13356
rect 10004 13300 10052 13356
rect 10108 13300 10156 13356
rect 10212 13300 10240 13356
rect 7008 12516 7036 12572
rect 7092 12516 7140 12572
rect 7196 12516 7244 12572
rect 7300 12516 7328 12572
rect 7008 11004 7328 12516
rect 7008 10948 7036 11004
rect 7092 10948 7140 11004
rect 7196 10948 7244 11004
rect 7300 10948 7328 11004
rect 7008 9436 7328 10948
rect 7420 12852 7476 12862
rect 7420 10500 7476 12796
rect 7420 10434 7476 10444
rect 9920 11788 10240 13300
rect 9920 11732 9948 11788
rect 10004 11732 10052 11788
rect 10108 11732 10156 11788
rect 10212 11732 10240 11788
rect 7008 9380 7036 9436
rect 7092 9380 7140 9436
rect 7196 9380 7244 9436
rect 7300 9380 7328 9436
rect 7008 7868 7328 9380
rect 7008 7812 7036 7868
rect 7092 7812 7140 7868
rect 7196 7812 7244 7868
rect 7300 7812 7328 7868
rect 7008 6300 7328 7812
rect 7008 6244 7036 6300
rect 7092 6244 7140 6300
rect 7196 6244 7244 6300
rect 7300 6244 7328 6300
rect 7008 4732 7328 6244
rect 7008 4676 7036 4732
rect 7092 4676 7140 4732
rect 7196 4676 7244 4732
rect 7300 4676 7328 4732
rect 7008 3164 7328 4676
rect 7008 3108 7036 3164
rect 7092 3108 7140 3164
rect 7196 3108 7244 3164
rect 7300 3108 7328 3164
rect 7008 3076 7328 3108
rect 9920 10220 10240 11732
rect 9920 10164 9948 10220
rect 10004 10164 10052 10220
rect 10108 10164 10156 10220
rect 10212 10164 10240 10220
rect 9920 8652 10240 10164
rect 9920 8596 9948 8652
rect 10004 8596 10052 8652
rect 10108 8596 10156 8652
rect 10212 8596 10240 8652
rect 9920 7084 10240 8596
rect 9920 7028 9948 7084
rect 10004 7028 10052 7084
rect 10108 7028 10156 7084
rect 10212 7028 10240 7084
rect 9920 5516 10240 7028
rect 9920 5460 9948 5516
rect 10004 5460 10052 5516
rect 10108 5460 10156 5516
rect 10212 5460 10240 5516
rect 9920 3948 10240 5460
rect 9920 3892 9948 3948
rect 10004 3892 10052 3948
rect 10108 3892 10156 3948
rect 10212 3892 10240 3948
rect 9920 3076 10240 3892
rect 12832 21980 13152 22796
rect 12832 21924 12860 21980
rect 12916 21924 12964 21980
rect 13020 21924 13068 21980
rect 13124 21924 13152 21980
rect 12832 20412 13152 21924
rect 12832 20356 12860 20412
rect 12916 20356 12964 20412
rect 13020 20356 13068 20412
rect 13124 20356 13152 20412
rect 12832 18844 13152 20356
rect 12832 18788 12860 18844
rect 12916 18788 12964 18844
rect 13020 18788 13068 18844
rect 13124 18788 13152 18844
rect 12832 17276 13152 18788
rect 12832 17220 12860 17276
rect 12916 17220 12964 17276
rect 13020 17220 13068 17276
rect 13124 17220 13152 17276
rect 12832 15708 13152 17220
rect 12832 15652 12860 15708
rect 12916 15652 12964 15708
rect 13020 15652 13068 15708
rect 13124 15652 13152 15708
rect 12832 14140 13152 15652
rect 12832 14084 12860 14140
rect 12916 14084 12964 14140
rect 13020 14084 13068 14140
rect 13124 14084 13152 14140
rect 12832 12572 13152 14084
rect 12832 12516 12860 12572
rect 12916 12516 12964 12572
rect 13020 12516 13068 12572
rect 13124 12516 13152 12572
rect 12832 11004 13152 12516
rect 12832 10948 12860 11004
rect 12916 10948 12964 11004
rect 13020 10948 13068 11004
rect 13124 10948 13152 11004
rect 12832 9436 13152 10948
rect 12832 9380 12860 9436
rect 12916 9380 12964 9436
rect 13020 9380 13068 9436
rect 13124 9380 13152 9436
rect 12832 7868 13152 9380
rect 12832 7812 12860 7868
rect 12916 7812 12964 7868
rect 13020 7812 13068 7868
rect 13124 7812 13152 7868
rect 12832 6300 13152 7812
rect 12832 6244 12860 6300
rect 12916 6244 12964 6300
rect 13020 6244 13068 6300
rect 13124 6244 13152 6300
rect 12832 4732 13152 6244
rect 12832 4676 12860 4732
rect 12916 4676 12964 4732
rect 13020 4676 13068 4732
rect 13124 4676 13152 4732
rect 12832 3164 13152 4676
rect 12832 3108 12860 3164
rect 12916 3108 12964 3164
rect 13020 3108 13068 3164
rect 13124 3108 13152 3164
rect 12832 3076 13152 3108
rect 15744 22764 16064 22796
rect 15744 22708 15772 22764
rect 15828 22708 15876 22764
rect 15932 22708 15980 22764
rect 16036 22708 16064 22764
rect 15744 21196 16064 22708
rect 15744 21140 15772 21196
rect 15828 21140 15876 21196
rect 15932 21140 15980 21196
rect 16036 21140 16064 21196
rect 15744 19628 16064 21140
rect 15744 19572 15772 19628
rect 15828 19572 15876 19628
rect 15932 19572 15980 19628
rect 16036 19572 16064 19628
rect 15744 18060 16064 19572
rect 15744 18004 15772 18060
rect 15828 18004 15876 18060
rect 15932 18004 15980 18060
rect 16036 18004 16064 18060
rect 15744 16492 16064 18004
rect 15744 16436 15772 16492
rect 15828 16436 15876 16492
rect 15932 16436 15980 16492
rect 16036 16436 16064 16492
rect 15744 14924 16064 16436
rect 15744 14868 15772 14924
rect 15828 14868 15876 14924
rect 15932 14868 15980 14924
rect 16036 14868 16064 14924
rect 15744 13356 16064 14868
rect 15744 13300 15772 13356
rect 15828 13300 15876 13356
rect 15932 13300 15980 13356
rect 16036 13300 16064 13356
rect 15744 11788 16064 13300
rect 15744 11732 15772 11788
rect 15828 11732 15876 11788
rect 15932 11732 15980 11788
rect 16036 11732 16064 11788
rect 15744 10220 16064 11732
rect 15744 10164 15772 10220
rect 15828 10164 15876 10220
rect 15932 10164 15980 10220
rect 16036 10164 16064 10220
rect 15744 8652 16064 10164
rect 15744 8596 15772 8652
rect 15828 8596 15876 8652
rect 15932 8596 15980 8652
rect 16036 8596 16064 8652
rect 15744 7084 16064 8596
rect 15744 7028 15772 7084
rect 15828 7028 15876 7084
rect 15932 7028 15980 7084
rect 16036 7028 16064 7084
rect 15744 5516 16064 7028
rect 15744 5460 15772 5516
rect 15828 5460 15876 5516
rect 15932 5460 15980 5516
rect 16036 5460 16064 5516
rect 15744 3948 16064 5460
rect 15744 3892 15772 3948
rect 15828 3892 15876 3948
rect 15932 3892 15980 3948
rect 16036 3892 16064 3948
rect 15744 3076 16064 3892
rect 18656 21980 18976 22796
rect 18656 21924 18684 21980
rect 18740 21924 18788 21980
rect 18844 21924 18892 21980
rect 18948 21924 18976 21980
rect 18656 20412 18976 21924
rect 18656 20356 18684 20412
rect 18740 20356 18788 20412
rect 18844 20356 18892 20412
rect 18948 20356 18976 20412
rect 18656 18844 18976 20356
rect 18656 18788 18684 18844
rect 18740 18788 18788 18844
rect 18844 18788 18892 18844
rect 18948 18788 18976 18844
rect 18656 17276 18976 18788
rect 18656 17220 18684 17276
rect 18740 17220 18788 17276
rect 18844 17220 18892 17276
rect 18948 17220 18976 17276
rect 18656 15708 18976 17220
rect 18656 15652 18684 15708
rect 18740 15652 18788 15708
rect 18844 15652 18892 15708
rect 18948 15652 18976 15708
rect 18656 14140 18976 15652
rect 18656 14084 18684 14140
rect 18740 14084 18788 14140
rect 18844 14084 18892 14140
rect 18948 14084 18976 14140
rect 18656 12572 18976 14084
rect 18656 12516 18684 12572
rect 18740 12516 18788 12572
rect 18844 12516 18892 12572
rect 18948 12516 18976 12572
rect 18656 11004 18976 12516
rect 18656 10948 18684 11004
rect 18740 10948 18788 11004
rect 18844 10948 18892 11004
rect 18948 10948 18976 11004
rect 18656 9436 18976 10948
rect 18656 9380 18684 9436
rect 18740 9380 18788 9436
rect 18844 9380 18892 9436
rect 18948 9380 18976 9436
rect 18656 7868 18976 9380
rect 18656 7812 18684 7868
rect 18740 7812 18788 7868
rect 18844 7812 18892 7868
rect 18948 7812 18976 7868
rect 18656 6300 18976 7812
rect 18656 6244 18684 6300
rect 18740 6244 18788 6300
rect 18844 6244 18892 6300
rect 18948 6244 18976 6300
rect 18656 4732 18976 6244
rect 18656 4676 18684 4732
rect 18740 4676 18788 4732
rect 18844 4676 18892 4732
rect 18948 4676 18976 4732
rect 18656 3164 18976 4676
rect 18656 3108 18684 3164
rect 18740 3108 18788 3164
rect 18844 3108 18892 3164
rect 18948 3108 18976 3164
rect 18656 3076 18976 3108
rect 21568 22764 21888 22796
rect 21568 22708 21596 22764
rect 21652 22708 21700 22764
rect 21756 22708 21804 22764
rect 21860 22708 21888 22764
rect 21568 21196 21888 22708
rect 21568 21140 21596 21196
rect 21652 21140 21700 21196
rect 21756 21140 21804 21196
rect 21860 21140 21888 21196
rect 21568 19628 21888 21140
rect 24480 21980 24800 22796
rect 24480 21924 24508 21980
rect 24564 21924 24612 21980
rect 24668 21924 24716 21980
rect 24772 21924 24800 21980
rect 24480 20412 24800 21924
rect 22652 20356 22708 20366
rect 22652 19908 22708 20300
rect 22652 19842 22708 19852
rect 24480 20356 24508 20412
rect 24564 20356 24612 20412
rect 24668 20356 24716 20412
rect 24772 20356 24800 20412
rect 21568 19572 21596 19628
rect 21652 19572 21700 19628
rect 21756 19572 21804 19628
rect 21860 19572 21888 19628
rect 21568 18060 21888 19572
rect 21568 18004 21596 18060
rect 21652 18004 21700 18060
rect 21756 18004 21804 18060
rect 21860 18004 21888 18060
rect 21568 16492 21888 18004
rect 21568 16436 21596 16492
rect 21652 16436 21700 16492
rect 21756 16436 21804 16492
rect 21860 16436 21888 16492
rect 21568 14924 21888 16436
rect 21568 14868 21596 14924
rect 21652 14868 21700 14924
rect 21756 14868 21804 14924
rect 21860 14868 21888 14924
rect 21568 13356 21888 14868
rect 21568 13300 21596 13356
rect 21652 13300 21700 13356
rect 21756 13300 21804 13356
rect 21860 13300 21888 13356
rect 21568 11788 21888 13300
rect 21568 11732 21596 11788
rect 21652 11732 21700 11788
rect 21756 11732 21804 11788
rect 21860 11732 21888 11788
rect 21568 10220 21888 11732
rect 21568 10164 21596 10220
rect 21652 10164 21700 10220
rect 21756 10164 21804 10220
rect 21860 10164 21888 10220
rect 21568 8652 21888 10164
rect 21568 8596 21596 8652
rect 21652 8596 21700 8652
rect 21756 8596 21804 8652
rect 21860 8596 21888 8652
rect 21568 7084 21888 8596
rect 21568 7028 21596 7084
rect 21652 7028 21700 7084
rect 21756 7028 21804 7084
rect 21860 7028 21888 7084
rect 21568 5516 21888 7028
rect 21568 5460 21596 5516
rect 21652 5460 21700 5516
rect 21756 5460 21804 5516
rect 21860 5460 21888 5516
rect 21568 3948 21888 5460
rect 21568 3892 21596 3948
rect 21652 3892 21700 3948
rect 21756 3892 21804 3948
rect 21860 3892 21888 3948
rect 21568 3076 21888 3892
rect 24480 18844 24800 20356
rect 24480 18788 24508 18844
rect 24564 18788 24612 18844
rect 24668 18788 24716 18844
rect 24772 18788 24800 18844
rect 24480 17276 24800 18788
rect 24480 17220 24508 17276
rect 24564 17220 24612 17276
rect 24668 17220 24716 17276
rect 24772 17220 24800 17276
rect 24480 15708 24800 17220
rect 24480 15652 24508 15708
rect 24564 15652 24612 15708
rect 24668 15652 24716 15708
rect 24772 15652 24800 15708
rect 24480 14140 24800 15652
rect 24480 14084 24508 14140
rect 24564 14084 24612 14140
rect 24668 14084 24716 14140
rect 24772 14084 24800 14140
rect 24480 12572 24800 14084
rect 24480 12516 24508 12572
rect 24564 12516 24612 12572
rect 24668 12516 24716 12572
rect 24772 12516 24800 12572
rect 24480 11004 24800 12516
rect 24480 10948 24508 11004
rect 24564 10948 24612 11004
rect 24668 10948 24716 11004
rect 24772 10948 24800 11004
rect 24480 9436 24800 10948
rect 24480 9380 24508 9436
rect 24564 9380 24612 9436
rect 24668 9380 24716 9436
rect 24772 9380 24800 9436
rect 24480 7868 24800 9380
rect 24480 7812 24508 7868
rect 24564 7812 24612 7868
rect 24668 7812 24716 7868
rect 24772 7812 24800 7868
rect 24480 6300 24800 7812
rect 24480 6244 24508 6300
rect 24564 6244 24612 6300
rect 24668 6244 24716 6300
rect 24772 6244 24800 6300
rect 24480 4732 24800 6244
rect 24480 4676 24508 4732
rect 24564 4676 24612 4732
rect 24668 4676 24716 4732
rect 24772 4676 24800 4732
rect 24480 3164 24800 4676
rect 24480 3108 24508 3164
rect 24564 3108 24612 3164
rect 24668 3108 24716 3164
rect 24772 3108 24800 3164
rect 24480 3076 24800 3108
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _197_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform 1 0 10192 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _198_
timestamp 1751914308
transform -1 0 13104 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform -1 0 11760 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _200_
timestamp 1751914308
transform 1 0 13328 0 1 14112
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _201_
timestamp 1751534193
transform -1 0 13104 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _202_
timestamp 1751534193
transform 1 0 21392 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _203_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform 1 0 11200 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _204_
timestamp 1751534193
transform -1 0 19936 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform -1 0 20608 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _206_
timestamp 1751534193
transform -1 0 23296 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform -1 0 21392 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _208_
timestamp 1751740063
transform 1 0 19824 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _209_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 19712 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _210_
timestamp 1751534193
transform -1 0 19824 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _211_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform -1 0 19824 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _212_
timestamp 1751740063
transform -1 0 18928 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _213_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform 1 0 21952 0 -1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform 1 0 21504 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _215_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform -1 0 22736 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _216_
timestamp 1751740063
transform 1 0 19488 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _217_
timestamp 1751534193
transform 1 0 19376 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _218_
timestamp 1751534193
transform -1 0 19712 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _219_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform -1 0 23632 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _220_
timestamp 1751740063
transform -1 0 23968 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _221_
timestamp 1751889408
transform -1 0 23184 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _222_
timestamp 1753182340
transform 1 0 21168 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _223_
timestamp 1751534193
transform -1 0 21840 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _224_
timestamp 1751532043
transform 1 0 23856 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _225_
timestamp 1753182340
transform 1 0 22624 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _226_
timestamp 1751740063
transform -1 0 23184 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _227_
timestamp 1753182340
transform 1 0 21392 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _228_
timestamp 1751534193
transform -1 0 19936 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _229_
timestamp 1751889408
transform -1 0 20944 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _230_
timestamp 1751740063
transform 1 0 21168 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _231_
timestamp 1753182340
transform 1 0 21168 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _232_
timestamp 1751534193
transform -1 0 19488 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _233_
timestamp 1751740063
transform -1 0 21056 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _234_
timestamp 1751889408
transform -1 0 21840 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _235_
timestamp 1753182340
transform -1 0 20944 0 1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _236_
timestamp 1751534193
transform -1 0 18592 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _237_
timestamp 1751740063
transform 1 0 19152 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _238_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform -1 0 23296 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _239_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform -1 0 22512 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _240_
timestamp 1753182340
transform 1 0 19936 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _241_
timestamp 1751534193
transform -1 0 18592 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _242_
timestamp 1751740063
transform -1 0 21952 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _243_
timestamp 1751889408
transform -1 0 20944 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _244_
timestamp 1753182340
transform 1 0 19824 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _245_
timestamp 1751534193
transform -1 0 18256 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _246_
timestamp 1751740063
transform 1 0 18704 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _247_
timestamp 1751889408
transform -1 0 21952 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _248_
timestamp 1753182340
transform 1 0 19488 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _249_
timestamp 1751534193
transform -1 0 18480 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _250_
timestamp 1751740063
transform 1 0 20608 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _251_
timestamp 1753960525
transform 1 0 20048 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _252_
timestamp 1751740063
transform 1 0 21168 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _253_
timestamp 1752061876
transform 1 0 11648 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _254_
timestamp 1751534193
transform 1 0 13328 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _255_
timestamp 1751534193
transform -1 0 8400 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _256_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform 1 0 14000 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _257_
timestamp 1751531619
transform 1 0 14784 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _258_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform 1 0 14896 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _259_
timestamp 1751534193
transform 1 0 15568 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _260_
timestamp 1751532043
transform -1 0 2912 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _261_
timestamp 1751889408
transform 1 0 12880 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _262_
timestamp 1751532043
transform 1 0 14336 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _263_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 14448 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _264_
timestamp 1751534193
transform 1 0 15120 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _265_
timestamp 1753868718
transform 1 0 14224 0 -1 15680
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _266_
timestamp 1751534193
transform 1 0 15456 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _267_
timestamp 1751534193
transform 1 0 8624 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _268_
timestamp 1751889808
transform 1 0 9632 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _269_
timestamp 1751534193
transform -1 0 11984 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _270_
timestamp 1751531619
transform 1 0 10864 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _271_
timestamp 1751889408
transform 1 0 10416 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _272_
timestamp 1751889408
transform 1 0 11200 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _273_
timestamp 1751534193
transform -1 0 6272 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _274_
timestamp 1751531619
transform -1 0 12768 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _275_
timestamp 1751532043
transform -1 0 9744 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _276_
timestamp 1753960525
transform 1 0 10528 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _277_
timestamp 1753960525
transform 1 0 11760 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _278_
timestamp 1751534193
transform 1 0 13328 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _279_
timestamp 1751740063
transform -1 0 10528 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _280_
timestamp 1751889808
transform -1 0 7504 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _281_
timestamp 1751531619
transform -1 0 8288 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _282_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform -1 0 8848 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _283_
timestamp 1752345181
transform 1 0 9072 0 1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _284_
timestamp 1753277515
transform -1 0 10976 0 -1 21952
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _285_
timestamp 1751905124
transform -1 0 13104 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _286_
timestamp 1751531619
transform 1 0 11200 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _287_
timestamp 1753441877
transform 1 0 11312 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _288_
timestamp 1751534193
transform -1 0 11760 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _289_
timestamp 1751905124
transform 1 0 4256 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _290_
timestamp 1751889408
transform 1 0 7280 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _291_
timestamp 1751534193
transform 1 0 8176 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _292_
timestamp 1751531619
transform -1 0 11088 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _293_
timestamp 1753182340
transform 1 0 7952 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _294_
timestamp 1751534193
transform 1 0 8848 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _295_
timestamp 1753277515
transform -1 0 23632 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _296_
timestamp 1753277515
transform 1 0 21952 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _297_
timestamp 1753277515
transform -1 0 23856 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _298_
timestamp 1753277515
transform -1 0 24416 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _299_
timestamp 1753172561
transform 1 0 22736 0 -1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _300_
timestamp 1753277515
transform 1 0 22064 0 1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _301_
timestamp 1753277515
transform 1 0 22736 0 -1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _302_
timestamp 1753277515
transform -1 0 24416 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _303_
timestamp 1753277515
transform -1 0 24304 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _304_
timestamp 1753172561
transform 1 0 22848 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _305_
timestamp 1753277515
transform -1 0 23632 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _306_
timestamp 1753277515
transform 1 0 22176 0 1 3136
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _307_
timestamp 1753277515
transform 1 0 21280 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _308_
timestamp 1753277515
transform -1 0 24416 0 -1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _309_
timestamp 1753172561
transform 1 0 22848 0 1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _310_
timestamp 1753182340
transform 1 0 22848 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _311_
timestamp 1751534193
transform -1 0 9072 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _312_
timestamp 1751532043
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _313_
timestamp 1753441877
transform -1 0 6608 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _314_
timestamp 1751534193
transform 1 0 9296 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _315_
timestamp 1751534193
transform -1 0 7952 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _316_
timestamp 1752061876
transform -1 0 3920 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _317_
timestamp 1751532043
transform -1 0 5264 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _318_
timestamp 1751889408
transform -1 0 5264 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _319_
timestamp 1751531619
transform 1 0 3696 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _320_
timestamp 1753277515
transform 1 0 5712 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _321_
timestamp 1753172561
transform 1 0 6048 0 1 15680
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _322_
timestamp 1751532043
transform -1 0 12096 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _323_
timestamp 1751534193
transform -1 0 11200 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _324_
timestamp 1753441877
transform -1 0 7728 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _325_
timestamp 1751532043
transform 1 0 4704 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _326_
timestamp 1753172561
transform 1 0 9408 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _327_
timestamp 1753441877
transform 1 0 8064 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _328_
timestamp 1751889408
transform -1 0 5376 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _329_
timestamp 1751889408
transform 1 0 3360 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _330_
timestamp 1753960525
transform 1 0 5712 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _331_
timestamp 1753868718
transform 1 0 3920 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _332_
timestamp 1753960525
transform -1 0 8848 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _333_
timestamp 1752061876
transform 1 0 6608 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _334_
timestamp 1751534193
transform -1 0 6944 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _335_
timestamp 1751740063
transform 1 0 2576 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_4  _336_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753952639
transform -1 0 6496 0 -1 15680
box -86 -86 2998 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _337_
timestamp 1753441877
transform 1 0 4144 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _338_
timestamp 1751531619
transform -1 0 6272 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _339_
timestamp 1751889408
transform 1 0 5376 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _340_
timestamp 1753172561
transform 1 0 8960 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _341_
timestamp 1753441877
transform -1 0 10528 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _342_
timestamp 1751534193
transform -1 0 8736 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _343_
timestamp 1753441877
transform 1 0 6384 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _344_
timestamp 1751889408
transform 1 0 7728 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _345_
timestamp 1751532043
transform -1 0 8960 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _346_
timestamp 1753441877
transform 1 0 7728 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _347_
timestamp 1751534193
transform -1 0 12992 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _348_
timestamp 1752345181
transform -1 0 7728 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _349_
timestamp 1751914308
transform 1 0 7504 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _350_
timestamp 1751889408
transform 1 0 9408 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _351_
timestamp 1751534193
transform -1 0 10080 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _352_
timestamp 1751534193
transform -1 0 4256 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _353_
timestamp 1751534193
transform -1 0 4928 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _354_
timestamp 1751740063
transform 1 0 3024 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _355_
timestamp 1751531619
transform 1 0 7280 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _356_
timestamp 1751531619
transform 1 0 9408 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _357_
timestamp 1751531619
transform 1 0 3808 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _358_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform 1 0 3696 0 1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _359_
timestamp 1751889408
transform -1 0 7280 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _360_
timestamp 1751905124
transform 1 0 5824 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _361_
timestamp 1753868718
transform 1 0 4592 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _362_
timestamp 1751534193
transform 1 0 5488 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _363_
timestamp 1753960525
transform 1 0 6944 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _364_
timestamp 1751531619
transform 1 0 7056 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _365_
timestamp 1752345181
transform -1 0 9072 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _366_
timestamp 1751534193
transform 1 0 10192 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _367_
timestamp 1753960525
transform 1 0 5488 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _368_
timestamp 1751534193
transform 1 0 6160 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _369_
timestamp 1751534193
transform 1 0 10528 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _370_
timestamp 1751534193
transform 1 0 11984 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _371_
timestamp 1751914308
transform 1 0 13328 0 -1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _372_
timestamp 1751534193
transform 1 0 7616 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _373_
timestamp 1751889408
transform 1 0 11984 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _374_
timestamp 1751534193
transform 1 0 14336 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _375_
timestamp 1751914308
transform 1 0 13776 0 1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _376_
timestamp 1751534193
transform 1 0 15568 0 -1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _377_
timestamp 1751914308
transform 1 0 13328 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _378_
timestamp 1751914308
transform 1 0 14448 0 1 10976
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _379_
timestamp 1751534193
transform 1 0 15904 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _380_
timestamp 1751534193
transform 1 0 11872 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _381_
timestamp 1751914308
transform 1 0 13440 0 -1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _382_
timestamp 1751914308
transform 1 0 14672 0 1 9408
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _383_
timestamp 1751534193
transform 1 0 16240 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _384_
timestamp 1751914308
transform 1 0 13328 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _385_
timestamp 1751914308
transform 1 0 14112 0 1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _386_
timestamp 1751534193
transform 1 0 15792 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _387_
timestamp 1751914308
transform 1 0 11536 0 1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _388_
timestamp 1751534193
transform 1 0 14560 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _389_
timestamp 1751914308
transform 1 0 13104 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _390_
timestamp 1751534193
transform 1 0 14448 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _391_
timestamp 1751914308
transform 1 0 10976 0 -1 7840
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _392_
timestamp 1751914308
transform -1 0 12880 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _393_
timestamp 1751534193
transform -1 0 11312 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _394_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform -1 0 18144 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _395_
timestamp 1751632746
transform -1 0 18816 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _396_
timestamp 1751632746
transform -1 0 19264 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _397_
timestamp 1751632746
transform -1 0 18480 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _398_
timestamp 1751632746
transform -1 0 16688 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _399_
timestamp 1751632746
transform 1 0 9744 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _400_
timestamp 1751632746
transform 1 0 9856 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _401_
timestamp 1751632746
transform 1 0 11536 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _402_
timestamp 1751632746
transform 1 0 18256 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _403_
timestamp 1751632746
transform 1 0 21280 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _404_
timestamp 1751632746
transform 1 0 16688 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _405_
timestamp 1751632746
transform 1 0 18928 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _406_
timestamp 1751632746
transform 1 0 21168 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _407_
timestamp 1751632746
transform 1 0 18368 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _408_
timestamp 1751632746
transform 1 0 18144 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _409_
timestamp 1751632746
transform 1 0 17248 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _410_
timestamp 1751632746
transform 1 0 17360 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _411_
timestamp 1751632746
transform 1 0 16800 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _412_
timestamp 1751632746
transform 1 0 17248 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _413_
timestamp 1751632746
transform 1 0 20832 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _414_
timestamp 1751632746
transform 1 0 15120 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _415_
timestamp 1751632746
transform 1 0 2016 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _416_
timestamp 1751632746
transform 1 0 1568 0 -1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _417_
timestamp 1751632746
transform 1 0 1568 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _418_
timestamp 1751632746
transform 1 0 1568 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _419_
timestamp 1751632746
transform -1 0 17360 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _420_
timestamp 1751632746
transform -1 0 17920 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _421_
timestamp 1751632746
transform 1 0 5488 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _422_
timestamp 1751632746
transform -1 0 16352 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _423_
timestamp 1751632746
transform 1 0 4704 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _424_
timestamp 1751632746
transform -1 0 14784 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _425_
timestamp 1751632746
transform 1 0 10080 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _426_
timestamp 1751632746
transform 1 0 9632 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _427_
timestamp 1751632746
transform 1 0 4928 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _428_
timestamp 1751632746
transform 1 0 6832 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _429_
timestamp 1751632746
transform 1 0 5152 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _430_
timestamp 1751632746
transform 1 0 9184 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _431_
timestamp 1751632746
transform 1 0 7504 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__204__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform -1 0 19264 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__217__A
timestamp 1751532392
transform -1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__251__D
timestamp 1751532392
transform -1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__401__CLK
timestamp 1751532392
transform 1 0 11312 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__415__CLK
timestamp 1751532392
transform 1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__416__CLK
timestamp 1751532392
transform 1 0 4592 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__417__CLK
timestamp 1751532392
transform 1 0 5712 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__418__CLK
timestamp 1751532392
transform -1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__421__CLK
timestamp 1751532392
transform 1 0 8736 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__423__CLK
timestamp 1751532392
transform -1 0 8736 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__430__CLK
timestamp 1751532392
transform -1 0 9184 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 10864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload1_A
timestamp 1751532392
transform 1 0 7840 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 21504 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input2_A
timestamp 1751532392
transform -1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input3_A
timestamp 1751532392
transform -1 0 22736 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input4_A
timestamp 1751532392
transform -1 0 22848 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input5_A
timestamp 1751532392
transform -1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input6_A
timestamp 1751532392
transform -1 0 23744 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input7_A
timestamp 1751532392
transform -1 0 22400 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input8_A
timestamp 1751532392
transform -1 0 24416 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input9_A
timestamp 1751532392
transform -1 0 23744 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input10_A
timestamp 1751532392
transform 1 0 24192 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input11_A
timestamp 1751532392
transform -1 0 22176 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input12_A
timestamp 1751532392
transform -1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input13_A
timestamp 1751532392
transform 1 0 13888 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 11536 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_0__f_wb_clk_i
timestamp 1751661108
transform -1 0 10864 0 1 9408
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_1__f_wb_clk_i
timestamp 1751661108
transform -1 0 8960 0 1 14112
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_2__f_wb_clk_i
timestamp 1751661108
transform 1 0 17248 0 -1 10976
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_2_3__f_wb_clk_i
timestamp 1751661108
transform 1 0 16240 0 1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 8064 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload1
timestamp 1751633659
transform 1 0 6832 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_18
timestamp 1751532351
transform 1 0 3360 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_36
timestamp 1751532351
transform 1 0 5376 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_52
timestamp 1751532351
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_70
timestamp 1751532351
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_86
timestamp 1751532351
transform 1 0 10976 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_104
timestamp 1751532351
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_120
timestamp 1751532351
transform 1 0 14784 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_138
timestamp 1751532351
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_154
timestamp 1751532351
transform 1 0 18592 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_172 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_176 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_200
timestamp 1751532440
transform 1 0 23744 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_2
timestamp 1751532351
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_18
timestamp 1751532351
transform 1 0 3360 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_34
timestamp 1751532351
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_50
timestamp 1751532351
transform 1 0 6944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_66
timestamp 1751532246
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_72
timestamp 1751532351
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_88
timestamp 1751532351
transform 1 0 11200 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_104
timestamp 1751532351
transform 1 0 12992 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_1_120
timestamp 1751532351
transform 1 0 14784 0 -1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_136
timestamp 1751532246
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_150 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 18144 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_205
timestamp 1751532423
transform 1 0 24304 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_2
timestamp 1751532351
transform 1 0 1568 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_18
timestamp 1751532351
transform 1 0 3360 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_34
timestamp 1751532423
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_37
timestamp 1751532351
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_53
timestamp 1751532351
transform 1 0 7280 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_69
timestamp 1751532246
transform 1 0 9072 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_73
timestamp 1751532440
transform 1 0 9520 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_102
timestamp 1751532440
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_104
timestamp 1751532423
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_107
timestamp 1751532351
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_123
timestamp 1751532351
transform 1 0 15120 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_2_139
timestamp 1751532351
transform 1 0 16912 0 1 4704
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_155
timestamp 1751532246
transform 1 0 18704 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_172
timestamp 1751532440
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_174
timestamp 1751532423
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_177
timestamp 1751532423
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_2
timestamp 1751532351
transform 1 0 1568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_18
timestamp 1751532351
transform 1 0 3360 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_34
timestamp 1751532351
transform 1 0 5152 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_50
timestamp 1751532351
transform 1 0 6944 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_66
timestamp 1751532246
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_72
timestamp 1751532312
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_80
timestamp 1751532440
transform 1 0 10304 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_82
timestamp 1751532423
transform 1 0 10528 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_89
timestamp 1751532440
transform 1 0 11312 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_103
timestamp 1751532440
transform 1 0 12880 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_123
timestamp 1751532351
transform 1 0 15120 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_139
timestamp 1751532423
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_142
timestamp 1751532312
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_150
timestamp 1751532423
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_199
timestamp 1751532423
transform 1 0 23632 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_2
timestamp 1751532351
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_18
timestamp 1751532351
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_34
timestamp 1751532423
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_37
timestamp 1751532351
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_53
timestamp 1751532440
transform 1 0 7280 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_82
timestamp 1751532312
transform 1 0 10528 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_90
timestamp 1751532423
transform 1 0 11424 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_103
timestamp 1751532440
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_107
timestamp 1751532440
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_109
timestamp 1751532423
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_177
timestamp 1751532440
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_179
timestamp 1751532423
transform 1 0 21392 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_196
timestamp 1751532440
transform 1 0 23296 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_2
timestamp 1751532351
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_18
timestamp 1751532351
transform 1 0 3360 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_67
timestamp 1751532440
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_69
timestamp 1751532423
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_72
timestamp 1751532312
transform 1 0 9408 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_80
timestamp 1751532246
transform 1 0 10304 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_84
timestamp 1751532440
transform 1 0 10752 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_98
timestamp 1751532312
transform 1 0 12320 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_106
timestamp 1751532423
transform 1 0 13216 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_119
timestamp 1751532312
transform 1 0 14672 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_127
timestamp 1751532440
transform 1 0 15568 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_135
timestamp 1751532246
transform 1 0 16464 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_139
timestamp 1751532423
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_142
timestamp 1751532312
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_198
timestamp 1751532440
transform 1 0 23520 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_2
timestamp 1751532351
transform 1 0 1568 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_18
timestamp 1751532351
transform 1 0 3360 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_34
timestamp 1751532423
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_103
timestamp 1751532440
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_107
timestamp 1751532246
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_111
timestamp 1751532440
transform 1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_113
timestamp 1751532423
transform 1 0 14000 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_153
timestamp 1751532312
transform 1 0 18480 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_161
timestamp 1751532423
transform 1 0 19376 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_169
timestamp 1751532246
transform 1 0 20272 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_173
timestamp 1751532440
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_177
timestamp 1751532246
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_181
timestamp 1751532440
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_183
timestamp 1751532423
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_191
timestamp 1751532423
transform 1 0 22736 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_2
timestamp 1751532351
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_18
timestamp 1751532312
transform 1 0 3360 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_26
timestamp 1751532246
transform 1 0 4256 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_30
timestamp 1751532440
transform 1 0 4704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_59
timestamp 1751532423
transform 1 0 7952 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_67
timestamp 1751532440
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_69
timestamp 1751532423
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_85
timestamp 1751532440
transform 1 0 10864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_105
timestamp 1751532440
transform 1 0 13104 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_107
timestamp 1751532423
transform 1 0 13328 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_120
timestamp 1751532312
transform 1 0 14784 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_128
timestamp 1751532246
transform 1 0 15680 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_132
timestamp 1751532423
transform 1 0 16128 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_139
timestamp 1751532423
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_142
timestamp 1751532351
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_160
timestamp 1751532351
transform 1 0 19264 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_176
timestamp 1751532312
transform 1 0 21056 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_184
timestamp 1751532246
transform 1 0 21952 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_188
timestamp 1751532440
transform 1 0 22400 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_2
timestamp 1751532351
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_18
timestamp 1751532351
transform 1 0 3360 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_34
timestamp 1751532423
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_37
timestamp 1751532312
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_45
timestamp 1751532423
transform 1 0 6384 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_85
timestamp 1751532312
transform 1 0 10864 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_93
timestamp 1751532423
transform 1 0 11760 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_100
timestamp 1751532246
transform 1 0 12544 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_104
timestamp 1751532423
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_131
timestamp 1751532440
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_166
timestamp 1751532312
transform 1 0 19936 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_174
timestamp 1751532423
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_204
timestamp 1751532440
transform 1 0 24192 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_2
timestamp 1751532312
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_10
timestamp 1751532246
transform 1 0 2464 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_14
timestamp 1751532423
transform 1 0 2912 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_50
timestamp 1751532423
transform 1 0 6944 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_69
timestamp 1751532423
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_72
timestamp 1751532440
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_101
timestamp 1751532246
transform 1 0 12656 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_105
timestamp 1751532440
transform 1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_119
timestamp 1751532312
transform 1 0 14672 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_127
timestamp 1751532440
transform 1 0 15568 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_129
timestamp 1751532423
transform 1 0 15792 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_136
timestamp 1751532246
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_167
timestamp 1751532312
transform 1 0 20048 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_175
timestamp 1751532440
transform 1 0 20944 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_183
timestamp 1751532440
transform 1 0 21840 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_185
timestamp 1751532423
transform 1 0 22064 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_199
timestamp 1751532423
transform 1 0 23632 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_2
timestamp 1751532351
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_18
timestamp 1751532440
transform 1 0 3360 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_20
timestamp 1751532423
transform 1 0 3584 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_47
timestamp 1751532246
transform 1 0 6608 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_51
timestamp 1751532440
transform 1 0 7056 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_60
timestamp 1751532312
transform 1 0 8064 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_68
timestamp 1751532246
transform 1 0 8960 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_107
timestamp 1751532312
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_115
timestamp 1751532440
transform 1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_156
timestamp 1751532246
transform 1 0 18816 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_166
timestamp 1751532312
transform 1 0 19936 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_174
timestamp 1751532423
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_202
timestamp 1751532440
transform 1 0 23968 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_11_2
timestamp 1751532351
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_18
timestamp 1751532440
transform 1 0 3360 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_43
timestamp 1751532440
transform 1 0 6160 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_67
timestamp 1751532440
transform 1 0 8848 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_69
timestamp 1751532423
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_122
timestamp 1751532246
transform 1 0 15008 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_126
timestamp 1751532423
transform 1 0 15456 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_133
timestamp 1751532246
transform 1 0 16240 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_137
timestamp 1751532440
transform 1 0 16688 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_139
timestamp 1751532423
transform 1 0 16912 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_142
timestamp 1751532312
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_150
timestamp 1751532440
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_205
timestamp 1751532423
transform 1 0 24304 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_29
timestamp 1751532440
transform 1 0 4592 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_33
timestamp 1751532440
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_66
timestamp 1751532440
transform 1 0 8736 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_97
timestamp 1751532312
transform 1 0 12208 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_107
timestamp 1751532246
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_150
timestamp 1751532246
transform 1 0 18144 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_154
timestamp 1751532440
transform 1 0 18592 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_162
timestamp 1751532312
transform 1 0 19488 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_170
timestamp 1751532246
transform 1 0 20384 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_174
timestamp 1751532423
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_177
timestamp 1751532312
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_199
timestamp 1751532423
transform 1 0 23632 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_2
timestamp 1751532312
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_14
timestamp 1751532312
transform 1 0 2912 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_22
timestamp 1751532246
transform 1 0 3808 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_32
timestamp 1751532312
transform 1 0 4928 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_40
timestamp 1751532246
transform 1 0 5824 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_44
timestamp 1751532440
transform 1 0 6272 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_67
timestamp 1751532440
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_69
timestamp 1751532423
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_72
timestamp 1751532312
transform 1 0 9408 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_80
timestamp 1751532246
transform 1 0 10304 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_84
timestamp 1751532423
transform 1 0 10752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_87
timestamp 1751532440
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_124
timestamp 1751532351
transform 1 0 15232 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_142
timestamp 1751532312
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_184
timestamp 1751532423
transform 1 0 21952 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_196
timestamp 1751532440
transform 1 0 23296 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_29
timestamp 1751532423
transform 1 0 4592 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_34
timestamp 1751532423
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_37
timestamp 1751532440
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_41
timestamp 1751532440
transform 1 0 5936 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_82
timestamp 1751532351
transform 1 0 10528 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_98
timestamp 1751532423
transform 1 0 12320 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_119
timestamp 1751532440
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_154
timestamp 1751532312
transform 1 0 18592 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_162
timestamp 1751532246
transform 1 0 19488 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_166
timestamp 1751532440
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_188
timestamp 1751532246
transform 1 0 22400 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_2
timestamp 1751532351
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_18
timestamp 1751532440
transform 1 0 3360 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_46
timestamp 1751532423
transform 1 0 6496 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_68
timestamp 1751532440
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_88
timestamp 1751532246
transform 1 0 11200 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_92
timestamp 1751532440
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_94
timestamp 1751532423
transform 1 0 11872 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_101
timestamp 1751532312
transform 1 0 12656 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_109
timestamp 1751532246
transform 1 0 13552 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_113
timestamp 1751532440
transform 1 0 14000 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_132
timestamp 1751532312
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_183
timestamp 1751532312
transform 1 0 21840 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_205
timestamp 1751532423
transform 1 0 24304 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_2
timestamp 1751532312
transform 1 0 1568 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_10
timestamp 1751532423
transform 1 0 2464 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_37
timestamp 1751532246
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_41
timestamp 1751532423
transform 1 0 5936 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_62
timestamp 1751532423
transform 1 0 8288 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_69
timestamp 1751532440
transform 1 0 9072 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_77
timestamp 1751532312
transform 1 0 9968 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_85
timestamp 1751532440
transform 1 0 10864 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_87
timestamp 1751532423
transform 1 0 11088 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_102
timestamp 1751532440
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_104
timestamp 1751532423
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_107
timestamp 1751532312
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_115
timestamp 1751532423
transform 1 0 14224 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_120
timestamp 1751532312
transform 1 0 14784 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_128
timestamp 1751532246
transform 1 0 15680 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_132
timestamp 1751532423
transform 1 0 16128 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_177
timestamp 1751532312
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_185
timestamp 1751532440
transform 1 0 22064 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_201
timestamp 1751532440
transform 1 0 23856 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_203
timestamp 1751532423
transform 1 0 24080 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_2
timestamp 1751532312
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_10
timestamp 1751532440
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_12
timestamp 1751532423
transform 1 0 2688 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_34
timestamp 1751532246
transform 1 0 5152 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_38
timestamp 1751532423
transform 1 0 5600 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_56
timestamp 1751532440
transform 1 0 7616 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_86
timestamp 1751532246
transform 1 0 10976 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_90
timestamp 1751532440
transform 1 0 11424 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_102
timestamp 1751532423
transform 1 0 12768 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_110
timestamp 1751532246
transform 1 0 13664 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_114
timestamp 1751532440
transform 1 0 14112 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_116
timestamp 1751532423
transform 1 0 14336 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_128
timestamp 1751532312
transform 1 0 15680 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_136
timestamp 1751532246
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_142
timestamp 1751532246
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_146
timestamp 1751532440
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_154
timestamp 1751532246
transform 1 0 18592 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_158
timestamp 1751532423
transform 1 0 19040 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_177
timestamp 1751532440
transform 1 0 21168 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_189
timestamp 1751532440
transform 1 0 22512 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_191
timestamp 1751532423
transform 1 0 22736 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_203
timestamp 1751532440
transform 1 0 24080 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_205
timestamp 1751532423
transform 1 0 24304 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_2
timestamp 1751532351
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_18
timestamp 1751532440
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_20
timestamp 1751532423
transform 1 0 3584 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_73
timestamp 1751532312
transform 1 0 9520 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_81
timestamp 1751532423
transform 1 0 10416 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_88
timestamp 1751532423
transform 1 0 11200 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_102
timestamp 1751532440
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_104
timestamp 1751532423
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_113
timestamp 1751532440
transform 1 0 14000 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_115
timestamp 1751532423
transform 1 0 14224 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_170
timestamp 1751532246
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_174
timestamp 1751532423
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_177
timestamp 1751532246
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_181
timestamp 1751532440
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_183
timestamp 1751532423
transform 1 0 21840 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_198
timestamp 1751532440
transform 1 0 23520 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_36
timestamp 1751532440
transform 1 0 5376 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_38
timestamp 1751532423
transform 1 0 5600 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_59
timestamp 1751532312
transform 1 0 7952 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_67
timestamp 1751532440
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_69
timestamp 1751532423
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_72
timestamp 1751532312
transform 1 0 9408 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_80
timestamp 1751532246
transform 1 0 10304 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_84
timestamp 1751532423
transform 1 0 10752 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_96
timestamp 1751532440
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_104
timestamp 1751532440
transform 1 0 12992 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_106
timestamp 1751532423
transform 1 0 13216 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_113
timestamp 1751532312
transform 1 0 14000 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_121
timestamp 1751532440
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_129
timestamp 1751532312
transform 1 0 15792 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_137
timestamp 1751532440
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_139
timestamp 1751532423
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_142
timestamp 1751532440
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_144
timestamp 1751532423
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_151
timestamp 1751532312
transform 1 0 18256 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_159
timestamp 1751532246
transform 1 0 19152 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_163
timestamp 1751532440
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_176
timestamp 1751532312
transform 1 0 21056 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_2
timestamp 1751532246
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_33
timestamp 1751532440
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_41
timestamp 1751532440
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_45
timestamp 1751532312
transform 1 0 6384 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_53
timestamp 1751532246
transform 1 0 7280 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_63
timestamp 1751532440
transform 1 0 8400 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_92
timestamp 1751532423
transform 1 0 11648 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_103
timestamp 1751532440
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_134
timestamp 1751532246
transform 1 0 16352 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_165
timestamp 1751532440
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_167
timestamp 1751532423
transform 1 0 20048 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_184
timestamp 1751532246
transform 1 0 21952 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_188
timestamp 1751532423
transform 1 0 22400 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_205
timestamp 1751532423
transform 1 0 24304 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_2
timestamp 1751532351
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_18
timestamp 1751532312
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_26
timestamp 1751532440
transform 1 0 4256 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_28
timestamp 1751532423
transform 1 0 4480 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_35
timestamp 1751532440
transform 1 0 5264 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_37
timestamp 1751532423
transform 1 0 5488 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_44
timestamp 1751532312
transform 1 0 6272 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_52
timestamp 1751532246
transform 1 0 7168 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_56
timestamp 1751532440
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_58
timestamp 1751532423
transform 1 0 7840 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_72
timestamp 1751532440
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_21_95
timestamp 1751532351
transform 1 0 11984 0 -1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_111
timestamp 1751532312
transform 1 0 13776 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_119
timestamp 1751532440
transform 1 0 14672 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_131
timestamp 1751532312
transform 1 0 16016 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_139
timestamp 1751532423
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_142
timestamp 1751532246
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_146
timestamp 1751532423
transform 1 0 17696 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_153
timestamp 1751532440
transform 1 0 18480 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_157
timestamp 1751532440
transform 1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_184
timestamp 1751532423
transform 1 0 21952 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_205
timestamp 1751532423
transform 1 0 24304 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_2
timestamp 1751532351
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_18
timestamp 1751532351
transform 1 0 3360 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_34
timestamp 1751532423
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_64
timestamp 1751532440
transform 1 0 8512 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_68
timestamp 1751532423
transform 1 0 8960 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_87
timestamp 1751532423
transform 1 0 11088 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_107
timestamp 1751532246
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_111
timestamp 1751532440
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_150
timestamp 1751532246
transform 1 0 18144 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_154
timestamp 1751532423
transform 1 0 18592 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_173
timestamp 1751532440
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_184
timestamp 1751532423
transform 1 0 21952 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_199
timestamp 1751532423
transform 1 0 23632 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_2
timestamp 1751532351
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_18
timestamp 1751532312
transform 1 0 3360 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_26
timestamp 1751532246
transform 1 0 4256 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_67
timestamp 1751532440
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_69
timestamp 1751532423
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_86
timestamp 1751532423
transform 1 0 10976 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_133
timestamp 1751532246
transform 1 0 16240 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_137
timestamp 1751532440
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_139
timestamp 1751532423
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_169
timestamp 1751532246
transform 1 0 20272 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_173
timestamp 1751532423
transform 1 0 20720 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_201
timestamp 1751532440
transform 1 0 23856 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_203
timestamp 1751532423
transform 1 0 24080 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_2
timestamp 1751532351
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_18
timestamp 1751532351
transform 1 0 3360 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_36
timestamp 1751532312
transform 1 0 5376 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_44
timestamp 1751532246
transform 1 0 6272 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_62
timestamp 1751532440
transform 1 0 8288 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_66
timestamp 1751532440
transform 1 0 8736 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_70
timestamp 1751532351
transform 1 0 9184 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_86
timestamp 1751532440
transform 1 0 10976 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_88
timestamp 1751532423
transform 1 0 11200 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_99
timestamp 1751532440
transform 1 0 12432 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_101
timestamp 1751532423
transform 1 0 12656 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_110
timestamp 1751532440
transform 1 0 13664 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_114
timestamp 1751532351
transform 1 0 14112 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_130
timestamp 1751532246
transform 1 0 15904 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_134
timestamp 1751532440
transform 1 0 16352 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_138
timestamp 1751532351
transform 1 0 16800 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_154
timestamp 1751532312
transform 1 0 18592 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform 1 0 21504 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input2
timestamp 1751534193
transform 1 0 19712 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input3
timestamp 1751534193
transform -1 0 22736 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input4
timestamp 1751534193
transform -1 0 24416 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input5
timestamp 1751534193
transform -1 0 24416 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input6
timestamp 1751534193
transform 1 0 23744 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input7
timestamp 1751534193
transform 1 0 23744 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input8
timestamp 1751534193
transform -1 0 24416 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input9
timestamp 1751534193
transform 1 0 23744 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input10
timestamp 1751534193
transform -1 0 24416 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input11
timestamp 1751534193
transform -1 0 22848 0 -1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input12
timestamp 1751534193
transform -1 0 24416 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input13
timestamp 1751534193
transform -1 0 13664 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output14
timestamp 1751661108
transform 1 0 21392 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 24640 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_26
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_27
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_28
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_29
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_30
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_31
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 24640 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_32
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_33
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 24640 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_34
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_35
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 24640 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_36
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_37
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_38
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_39
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_40
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_41
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 24640 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_42
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_43
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 24640 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_44
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_45
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_46
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_47
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_48
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_49
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 24640 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_50
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_51
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_52
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_53
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_54
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_55
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_56
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_57
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_58
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_59
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_60
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_61
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_62
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_63
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_64
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_65
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_66
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_67
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_68
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_69
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_70
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_71
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_72
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_73
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_74
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_75
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_76
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_77
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_78
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_79
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_80
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_81
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_82
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_83
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_84
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_85
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_86
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_87
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_88
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_89
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_90
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_91
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_92
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_93
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_94
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_95
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_96
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_97
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_98
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_99
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_100
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_101
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_102
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_103
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_104
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_105
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_106
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_107
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_108
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_109
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_110
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_111
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_112
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_113
timestamp 1751532504
transform 1 0 5152 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_114
timestamp 1751532504
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_115
timestamp 1751532504
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_116
timestamp 1751532504
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_117
timestamp 1751532504
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_118
timestamp 1751532504
transform 1 0 24192 0 1 21952
box -86 -86 310 870
<< labels >>
flabel metal3 s 25200 1792 26000 1904 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 25200 21952 26000 22064 0 FreeSans 448 0 0 0 custom_settings[10]
port 1 nsew signal input
flabel metal3 s 25200 23968 26000 24080 0 FreeSans 448 0 0 0 custom_settings[11]
port 2 nsew signal input
flabel metal3 s 25200 3808 26000 3920 0 FreeSans 448 0 0 0 custom_settings[1]
port 3 nsew signal input
flabel metal3 s 25200 5824 26000 5936 0 FreeSans 448 0 0 0 custom_settings[2]
port 4 nsew signal input
flabel metal3 s 25200 7840 26000 7952 0 FreeSans 448 0 0 0 custom_settings[3]
port 5 nsew signal input
flabel metal3 s 25200 9856 26000 9968 0 FreeSans 448 0 0 0 custom_settings[4]
port 6 nsew signal input
flabel metal3 s 25200 11872 26000 11984 0 FreeSans 448 0 0 0 custom_settings[5]
port 7 nsew signal input
flabel metal3 s 25200 13888 26000 14000 0 FreeSans 448 0 0 0 custom_settings[6]
port 8 nsew signal input
flabel metal3 s 25200 15904 26000 16016 0 FreeSans 448 0 0 0 custom_settings[7]
port 9 nsew signal input
flabel metal3 s 25200 17920 26000 18032 0 FreeSans 448 0 0 0 custom_settings[8]
port 10 nsew signal input
flabel metal3 s 25200 19936 26000 20048 0 FreeSans 448 0 0 0 custom_settings[9]
port 11 nsew signal input
flabel metal2 s 21280 25200 21392 26000 0 FreeSans 448 90 0 0 io_out
port 12 nsew signal output
flabel metal2 s 12768 25200 12880 26000 0 FreeSans 448 90 0 0 rst_n
port 13 nsew signal input
flabel metal4 s 4096 3076 4416 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 9920 3076 10240 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 15744 3076 16064 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 21568 3076 21888 22796 0 FreeSans 1280 90 0 0 vdd
port 14 nsew power bidirectional
flabel metal4 s 7008 3076 7328 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 12832 3076 13152 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 18656 3076 18976 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal4 s 24480 3076 24800 22796 0 FreeSans 1280 90 0 0 vss
port 15 nsew ground bidirectional
flabel metal2 s 4256 25200 4368 26000 0 FreeSans 448 90 0 0 wb_clk_i
port 16 nsew signal input
rlabel metal1 12992 22736 12992 22736 0 vdd
rlabel via1 13072 21952 13072 21952 0 vss
rlabel metal3 10304 11368 10304 11368 0 _000_
rlabel metal2 10024 9436 10024 9436 0 _001_
rlabel metal2 5824 8456 5824 8456 0 _002_
rlabel metal2 7672 8372 7672 8372 0 _003_
rlabel metal2 5992 7728 5992 7728 0 _004_
rlabel metal3 16632 12376 16632 12376 0 _005_
rlabel metal3 17136 10808 17136 10808 0 _006_
rlabel metal3 17528 9240 17528 9240 0 _007_
rlabel metal3 16912 7672 16912 7672 0 _008_
rlabel metal2 14784 6104 14784 6104 0 _009_
rlabel metal2 10584 5432 10584 5432 0 _010_
rlabel metal2 11032 8792 11032 8792 0 _011_
rlabel metal2 12376 14000 12376 14000 0 _012_
rlabel metal2 19096 4696 19096 4696 0 _013_
rlabel metal3 21140 4312 21140 4312 0 _014_
rlabel metal2 17528 7056 17528 7056 0 _015_
rlabel metal2 19768 7756 19768 7756 0 _016_
rlabel metal3 21728 9912 21728 9912 0 _017_
rlabel metal2 19488 11592 19488 11592 0 _018_
rlabel metal2 19040 13160 19040 13160 0 _019_
rlabel metal2 18144 14728 18144 14728 0 _020_
rlabel metal2 18200 17360 18200 17360 0 _021_
rlabel metal2 17864 18928 17864 18928 0 _022_
rlabel metal2 18088 20832 18088 20832 0 _023_
rlabel metal2 21560 20580 21560 20580 0 _024_
rlabel metal2 16072 20888 16072 20888 0 _025_
rlabel metal4 6776 17696 6776 17696 0 _026_
rlabel metal3 4228 14280 4228 14280 0 _027_
rlabel metal2 2688 14224 2688 14224 0 _028_
rlabel metal2 3864 12656 3864 12656 0 _029_
rlabel metal2 16520 17976 16520 17976 0 _030_
rlabel metal2 17080 14840 17080 14840 0 _031_
rlabel metal2 5880 20496 5880 20496 0 _032_
rlabel metal2 13720 18816 13720 18816 0 _033_
rlabel metal3 6776 21448 6776 21448 0 _034_
rlabel metal3 12656 21448 12656 21448 0 _035_
rlabel metal2 5208 12180 5208 12180 0 _036_
rlabel metal2 8344 7000 8344 7000 0 _037_
rlabel metal2 23184 14728 23184 14728 0 _038_
rlabel metal3 23576 18424 23576 18424 0 _039_
rlabel metal2 23352 17612 23352 17612 0 _040_
rlabel metal2 23016 5208 23016 5208 0 _041_
rlabel metal2 23464 4396 23464 4396 0 _042_
rlabel metal3 23128 5096 23128 5096 0 _043_
rlabel metal3 23576 6888 23576 6888 0 _044_
rlabel metal3 24192 5208 24192 5208 0 _045_
rlabel metal2 8344 16912 8344 16912 0 _046_
rlabel metal2 6328 17528 6328 17528 0 _047_
rlabel metal2 5880 18704 5880 18704 0 _048_
rlabel metal2 7560 15344 7560 15344 0 _049_
rlabel metal2 6328 15960 6328 15960 0 _050_
rlabel metal2 7672 16352 7672 16352 0 _051_
rlabel metal2 4088 16940 4088 16940 0 _052_
rlabel metal2 4984 17584 4984 17584 0 _053_
rlabel metal3 4452 17640 4452 17640 0 _054_
rlabel metal2 6888 16352 6888 16352 0 _055_
rlabel metal2 7224 16576 7224 16576 0 _056_
rlabel metal2 7448 15400 7448 15400 0 _057_
rlabel metal2 11144 17752 11144 17752 0 _058_
rlabel metal2 7282 15232 7282 15232 0 _059_
rlabel metal2 4760 14784 4760 14784 0 _060_
rlabel metal3 10080 15288 10080 15288 0 _061_
rlabel metal2 10248 15400 10248 15400 0 _062_
rlabel metal2 3640 16408 3640 16408 0 _063_
rlabel metal2 4424 16940 4424 16940 0 _064_
rlabel metal2 6692 16968 6692 16968 0 _065_
rlabel metal2 5012 16632 5012 16632 0 _066_
rlabel metal2 7700 17640 7700 17640 0 _067_
rlabel metal2 8154 14019 8154 14019 0 _068_
rlabel metal2 6810 12451 6810 12451 0 _069_
rlabel metal2 3192 15960 3192 15960 0 _070_
rlabel metal2 4356 12451 4356 12451 0 _071_
rlabel metal3 5432 12936 5432 12936 0 _072_
rlabel metal2 5600 12152 5600 12152 0 _073_
rlabel metal2 5992 11480 5992 11480 0 _074_
rlabel metal2 9464 13384 9464 13384 0 _075_
rlabel metal2 8904 14112 8904 14112 0 _076_
rlabel metal2 6664 12208 6664 12208 0 _077_
rlabel metal3 7784 12152 7784 12152 0 _078_
rlabel metal2 7896 14112 7896 14112 0 _079_
rlabel metal2 7112 12992 7112 12992 0 _080_
rlabel metal2 8232 19208 8232 19208 0 _081_
rlabel metal2 7224 13552 7224 13552 0 _082_
rlabel metal3 9137 12152 9137 12152 0 _083_
rlabel metal2 9912 11368 9912 11368 0 _084_
rlabel metal3 3696 13720 3696 13720 0 _085_
rlabel metal2 7616 9800 7616 9800 0 _086_
rlabel metal2 7560 11172 7560 11172 0 _087_
rlabel metal2 4424 10444 4424 10444 0 _088_
rlabel metal2 5096 11312 5096 11312 0 _089_
rlabel metal3 7140 10024 7140 10024 0 _090_
rlabel via2 5320 10598 5320 10598 0 _091_
rlabel metal2 5572 10360 5572 10360 0 _092_
rlabel metal2 8008 12040 8008 12040 0 _093_
rlabel metal2 7672 10500 7672 10500 0 _094_
rlabel metal2 8680 10136 8680 10136 0 _095_
rlabel metal2 6216 8316 6216 8316 0 _096_
rlabel metal2 10360 12096 10360 12096 0 _097_
rlabel metal2 12376 15904 12376 15904 0 _098_
rlabel metal2 14345 10696 14345 10696 0 _099_
rlabel metal3 11872 16072 11872 16072 0 _100_
rlabel metal3 13468 16072 13468 16072 0 _101_
rlabel metal2 14224 8232 14224 8232 0 _102_
rlabel metal2 15624 12488 15624 12488 0 _103_
rlabel metal2 14410 10080 14410 10080 0 _104_
rlabel metal2 15960 10920 15960 10920 0 _105_
rlabel metal3 12936 8344 12936 8344 0 _106_
rlabel metal2 14522 9184 14522 9184 0 _107_
rlabel metal2 16016 9016 16016 9016 0 _108_
rlabel via1 14429 7560 14429 7560 0 _109_
rlabel metal2 15848 7616 15848 7616 0 _110_
rlabel metal2 13440 6244 13440 6244 0 _111_
rlabel metal3 12992 5992 12992 5992 0 _112_
rlabel metal2 14345 5880 14345 5880 0 _113_
rlabel metal2 12544 6132 12544 6132 0 _114_
rlabel metal3 11527 5880 11527 5880 0 _115_
rlabel metal2 12768 9324 12768 9324 0 _116_
rlabel metal2 11863 9016 11863 9016 0 _117_
rlabel metal3 13729 14504 13729 14504 0 _118_
rlabel metal2 20272 5880 20272 5880 0 _119_
rlabel metal2 19656 9800 19656 9800 0 _120_
rlabel metal2 20048 6664 20048 6664 0 _121_
rlabel metal2 21112 5768 21112 5768 0 _122_
rlabel metal2 20832 6048 20832 6048 0 _123_
rlabel metal2 20496 6664 20496 6664 0 _124_
rlabel metal2 19824 5096 19824 5096 0 _125_
rlabel metal2 18536 6216 18536 6216 0 _126_
rlabel metal2 22568 7784 22568 7784 0 _127_
rlabel metal2 22372 6888 22372 6888 0 _128_
rlabel metal2 22120 8316 22120 8316 0 _129_
rlabel metal2 19712 19992 19712 19992 0 _130_
rlabel metal2 21336 14560 21336 14560 0 _131_
rlabel metal2 23688 11480 23688 11480 0 _132_
rlabel metal2 22680 11416 22680 11416 0 _133_
rlabel metal2 22540 10696 22540 10696 0 _134_
rlabel metal2 21784 10752 21784 10752 0 _135_
rlabel metal2 23240 12236 23240 12236 0 _136_
rlabel metal2 22008 12348 22008 12348 0 _137_
rlabel metal2 22232 11816 22232 11816 0 _138_
rlabel metal2 22120 12180 22120 12180 0 _139_
rlabel metal2 21532 14504 21532 14504 0 _140_
rlabel metal2 21784 14056 21784 14056 0 _141_
rlabel metal2 21448 13916 21448 13916 0 _142_
rlabel metal2 20440 15596 20440 15596 0 _143_
rlabel metal2 20160 16072 20160 16072 0 _144_
rlabel metal2 18536 14728 18536 14728 0 _145_
rlabel via2 20440 16869 20440 16869 0 _146_
rlabel metal3 22400 15848 22400 15848 0 _147_
rlabel metal2 20776 16940 20776 16940 0 _148_
rlabel metal2 18536 16968 18536 16968 0 _149_
rlabel metal2 21336 19096 21336 19096 0 _150_
rlabel metal2 20664 20160 20664 20160 0 _151_
rlabel metal3 19208 18424 19208 18424 0 _152_
rlabel metal2 19936 20748 19936 20748 0 _153_
rlabel metal3 21252 21000 21252 21000 0 _154_
rlabel metal2 18424 20104 18424 20104 0 _155_
rlabel metal2 21224 21224 21224 21224 0 _156_
rlabel via1 21616 20006 21616 20006 0 _157_
rlabel metal2 13216 16856 13216 16856 0 _158_
rlabel metal3 11536 20216 11536 20216 0 _159_
rlabel metal2 8064 21112 8064 21112 0 _160_
rlabel metal2 14952 21084 14952 21084 0 _161_
rlabel metal2 15322 20291 15322 20291 0 _162_
rlabel metal2 15680 19880 15680 19880 0 _163_
rlabel via2 14728 16870 14728 16870 0 _164_
rlabel metal2 14532 16296 14532 16296 0 _165_
rlabel metal2 15428 16968 15428 16968 0 _166_
rlabel metal2 15372 15288 15372 15288 0 _167_
rlabel metal2 9856 20776 9856 20776 0 _168_
rlabel metal2 10500 19768 10500 19768 0 _169_
rlabel metal1 12488 20216 12488 20216 0 _170_
rlabel metal2 11144 18396 11144 18396 0 _171_
rlabel metal2 11480 19880 11480 19880 0 _172_
rlabel metal2 6216 19936 6216 19936 0 _173_
rlabel metal2 12264 18452 12264 18452 0 _174_
rlabel metal3 9884 19208 9884 19208 0 _175_
rlabel metal3 11676 19208 11676 19208 0 _176_
rlabel metal2 13384 18760 13384 18760 0 _177_
rlabel metal2 7224 22232 7224 22232 0 _178_
rlabel metal2 7784 22624 7784 22624 0 _179_
rlabel metal2 7868 21616 7868 21616 0 _180_
rlabel metal2 9576 21224 9576 21224 0 _181_
rlabel metal2 9856 21336 9856 21336 0 _182_
rlabel metal3 11928 20776 11928 20776 0 _183_
rlabel metal2 11758 22456 11758 22456 0 _184_
rlabel metal2 11704 21784 11704 21784 0 _185_
rlabel metal2 7952 7896 7952 7896 0 _186_
rlabel metal3 9744 20552 9744 20552 0 _187_
rlabel metal2 8232 20020 8232 20020 0 _188_
rlabel metal2 6440 17528 6440 17528 0 _189_
rlabel metal2 22344 13272 22344 13272 0 _190_
rlabel metal2 23184 15372 23184 15372 0 _191_
rlabel metal3 23072 15288 23072 15288 0 _192_
rlabel metal3 24024 8344 24024 8344 0 _193_
rlabel metal2 23016 16744 23016 16744 0 _194_
rlabel metal2 22960 18424 22960 18424 0 _195_
rlabel metal2 23464 19012 23464 19012 0 _196_
rlabel metal3 21840 5880 21840 5880 0 baud_delay\[0\]
rlabel metal3 22502 20776 22502 20776 0 baud_delay\[10\]
rlabel metal2 20552 21224 20552 21224 0 baud_delay\[11\]
rlabel metal2 24024 4592 24024 4592 0 baud_delay\[1\]
rlabel metal2 22587 5964 22587 5964 0 baud_delay\[2\]
rlabel metal2 23128 7560 23128 7560 0 baud_delay\[3\]
rlabel metal2 23912 9632 23912 9632 0 baud_delay\[4\]
rlabel metal2 22587 12852 22587 12852 0 baud_delay\[5\]
rlabel metal2 23128 13888 23128 13888 0 baud_delay\[6\]
rlabel metal2 22568 14952 22568 14952 0 baud_delay\[7\]
rlabel metal3 19768 17528 19768 17528 0 baud_delay\[8\]
rlabel metal3 22521 19208 22521 19208 0 baud_delay\[9\]
rlabel metal2 13664 10892 13664 10892 0 char_at\[0\]
rlabel metal2 13664 9884 13664 9884 0 char_at\[1\]
rlabel metal2 13776 8932 13776 8932 0 char_at\[2\]
rlabel metal2 13664 7532 13664 7532 0 char_at\[3\]
rlabel metal3 11060 6664 11060 6664 0 char_at\[4\]
rlabel metal2 11312 7364 11312 7364 0 char_at\[5\]
rlabel metal2 10528 12236 10528 12236 0 char_at\[6\]
rlabel metal2 5096 18368 5096 18368 0 char_pointer\[0\]
rlabel metal2 5320 18816 5320 18816 0 char_pointer\[1\]
rlabel metal2 4590 15988 4590 15988 0 char_pointer\[2\]
rlabel metal2 3752 14952 3752 14952 0 char_pointer\[3\]
rlabel metal2 17752 11941 17752 11941 0 clknet_0_wb_clk_i
rlabel metal2 6888 8288 6888 8288 0 clknet_2_0__leaf_wb_clk_i
rlabel metal2 5544 20496 5544 20496 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 21336 4704 21336 4704 0 clknet_2_2__leaf_wb_clk_i
rlabel metal2 14728 21168 14728 21168 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 21560 2688 21560 2688 0 custom_settings[0]
rlabel metal3 22260 22232 22260 22232 0 custom_settings[10]
rlabel metal3 24066 24024 24066 24024 0 custom_settings[11]
rlabel metal2 24360 4872 24360 4872 0 custom_settings[1]
rlabel metal2 24304 6664 24304 6664 0 custom_settings[2]
rlabel metal2 23800 7560 23800 7560 0 custom_settings[3]
rlabel metal2 23800 10360 23800 10360 0 custom_settings[4]
rlabel metal2 24304 11704 24304 11704 0 custom_settings[5]
rlabel metal3 24430 13944 24430 13944 0 custom_settings[6]
rlabel metal3 24766 15960 24766 15960 0 custom_settings[7]
rlabel metal2 22792 18200 22792 18200 0 custom_settings[8]
rlabel metal2 24360 20720 24360 20720 0 custom_settings[9]
rlabel metal2 8288 20664 8288 20664 0 frame_counter\[0\]
rlabel via2 9688 20756 9688 20756 0 frame_counter\[1\]
rlabel metal2 7448 22008 7448 22008 0 frame_counter\[2\]
rlabel metal2 12152 21448 12152 21448 0 frame_counter\[3\]
rlabel metal3 21952 22568 21952 22568 0 io_out
rlabel metal2 22324 4844 22324 4844 0 net1
rlabel metal2 23800 16072 23800 16072 0 net10
rlabel metal3 22120 17752 22120 17752 0 net11
rlabel metal2 24248 19208 24248 19208 0 net12
rlabel metal2 12880 22120 12880 22120 0 net13
rlabel metal2 14840 20832 14840 20832 0 net14
rlabel metal2 22120 20776 22120 20776 0 net2
rlabel metal2 22848 19992 22848 19992 0 net3
rlabel metal2 22232 3528 22232 3528 0 net4
rlabel metal3 23744 5880 23744 5880 0 net5
rlabel metal2 24192 7672 24192 7672 0 net6
rlabel metal2 24248 9688 24248 9688 0 net7
rlabel metal3 23744 12936 23744 12936 0 net8
rlabel metal2 24192 13944 24192 13944 0 net9
rlabel metal3 13216 22344 13216 22344 0 rst_n
rlabel metal2 14616 17976 14616 17976 0 uart_frame\[0\]
rlabel metal2 14616 13216 14616 13216 0 uart_frame\[1\]
rlabel metal2 15288 10976 15288 10976 0 uart_frame\[2\]
rlabel metal3 14840 9800 14840 9800 0 uart_frame\[3\]
rlabel metal2 14952 8288 14952 8288 0 uart_frame\[4\]
rlabel metal2 13944 7112 13944 7112 0 uart_frame\[5\]
rlabel metal2 12040 5544 12040 5544 0 uart_frame\[6\]
rlabel metal2 12040 7448 12040 7448 0 uart_frame\[7\]
rlabel metal2 15120 14392 15120 14392 0 uart_frame\[8\]
rlabel metal2 14168 14896 14168 14896 0 uart_frame\[9\]
rlabel metal2 4424 22904 4424 22904 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 26000 26000
<< end >>
