magic
tech gf180mcuD
magscale 1 5
timestamp 1754400677
<< nwell >>
rect 629 1525 169331 78443
<< obsm1 >>
rect 672 1538 169288 78430
<< metal2 >>
rect 1232 0 1288 400
rect 3808 0 3864 400
rect 6384 0 6440 400
rect 8960 0 9016 400
rect 11536 0 11592 400
rect 14112 0 14168 400
rect 16688 0 16744 400
rect 19264 0 19320 400
rect 21840 0 21896 400
rect 24416 0 24472 400
rect 26992 0 27048 400
rect 29568 0 29624 400
rect 32144 0 32200 400
rect 34720 0 34776 400
rect 37296 0 37352 400
rect 39872 0 39928 400
rect 42448 0 42504 400
rect 45024 0 45080 400
rect 47600 0 47656 400
rect 50176 0 50232 400
rect 52752 0 52808 400
rect 55328 0 55384 400
rect 57904 0 57960 400
rect 60480 0 60536 400
rect 63056 0 63112 400
rect 65632 0 65688 400
rect 68208 0 68264 400
rect 70784 0 70840 400
rect 73360 0 73416 400
rect 75936 0 75992 400
rect 78512 0 78568 400
rect 81088 0 81144 400
rect 83664 0 83720 400
rect 86240 0 86296 400
rect 88816 0 88872 400
rect 91392 0 91448 400
rect 93968 0 94024 400
rect 96544 0 96600 400
rect 99120 0 99176 400
rect 101696 0 101752 400
rect 104272 0 104328 400
rect 106848 0 106904 400
rect 109424 0 109480 400
rect 112000 0 112056 400
rect 114576 0 114632 400
rect 117152 0 117208 400
rect 119728 0 119784 400
rect 122304 0 122360 400
rect 124880 0 124936 400
rect 127456 0 127512 400
rect 130032 0 130088 400
rect 132608 0 132664 400
rect 135184 0 135240 400
rect 137760 0 137816 400
rect 140336 0 140392 400
rect 142912 0 142968 400
rect 145488 0 145544 400
rect 148064 0 148120 400
rect 150640 0 150696 400
rect 153216 0 153272 400
rect 155792 0 155848 400
rect 158368 0 158424 400
rect 160944 0 161000 400
rect 163520 0 163576 400
rect 166096 0 166152 400
rect 168672 0 168728 400
<< obsm2 >>
rect 14 430 169134 78419
rect 14 345 1202 430
rect 1318 345 3778 430
rect 3894 345 6354 430
rect 6470 345 8930 430
rect 9046 345 11506 430
rect 11622 345 14082 430
rect 14198 345 16658 430
rect 16774 345 19234 430
rect 19350 345 21810 430
rect 21926 345 24386 430
rect 24502 345 26962 430
rect 27078 345 29538 430
rect 29654 345 32114 430
rect 32230 345 34690 430
rect 34806 345 37266 430
rect 37382 345 39842 430
rect 39958 345 42418 430
rect 42534 345 44994 430
rect 45110 345 47570 430
rect 47686 345 50146 430
rect 50262 345 52722 430
rect 52838 345 55298 430
rect 55414 345 57874 430
rect 57990 345 60450 430
rect 60566 345 63026 430
rect 63142 345 65602 430
rect 65718 345 68178 430
rect 68294 345 70754 430
rect 70870 345 73330 430
rect 73446 345 75906 430
rect 76022 345 78482 430
rect 78598 345 81058 430
rect 81174 345 83634 430
rect 83750 345 86210 430
rect 86326 345 88786 430
rect 88902 345 91362 430
rect 91478 345 93938 430
rect 94054 345 96514 430
rect 96630 345 99090 430
rect 99206 345 101666 430
rect 101782 345 104242 430
rect 104358 345 106818 430
rect 106934 345 109394 430
rect 109510 345 111970 430
rect 112086 345 114546 430
rect 114662 345 117122 430
rect 117238 345 119698 430
rect 119814 345 122274 430
rect 122390 345 124850 430
rect 124966 345 127426 430
rect 127542 345 130002 430
rect 130118 345 132578 430
rect 132694 345 135154 430
rect 135270 345 137730 430
rect 137846 345 140306 430
rect 140422 345 142882 430
rect 142998 345 145458 430
rect 145574 345 148034 430
rect 148150 345 150610 430
rect 150726 345 153186 430
rect 153302 345 155762 430
rect 155878 345 158338 430
rect 158454 345 160914 430
rect 161030 345 163490 430
rect 163606 345 166066 430
rect 166182 345 168642 430
rect 168758 345 169134 430
<< metal3 >>
rect 0 77504 400 77560
rect 169600 77504 170000 77560
rect 169600 75152 170000 75208
rect 0 73920 400 73976
rect 169600 72800 170000 72856
rect 169600 70448 170000 70504
rect 0 70336 400 70392
rect 169600 68096 170000 68152
rect 0 66752 400 66808
rect 169600 65744 170000 65800
rect 169600 63392 170000 63448
rect 0 63168 400 63224
rect 169600 61040 170000 61096
rect 0 59584 400 59640
rect 169600 58688 170000 58744
rect 169600 56336 170000 56392
rect 0 56000 400 56056
rect 169600 53984 170000 54040
rect 0 52416 400 52472
rect 169600 51632 170000 51688
rect 169600 49280 170000 49336
rect 0 48832 400 48888
rect 169600 46928 170000 46984
rect 0 45248 400 45304
rect 169600 44576 170000 44632
rect 169600 42224 170000 42280
rect 0 41664 400 41720
rect 169600 39872 170000 39928
rect 0 38080 400 38136
rect 169600 37520 170000 37576
rect 169600 35168 170000 35224
rect 0 34496 400 34552
rect 169600 32816 170000 32872
rect 0 30912 400 30968
rect 169600 30464 170000 30520
rect 169600 28112 170000 28168
rect 0 27328 400 27384
rect 169600 25760 170000 25816
rect 0 23744 400 23800
rect 169600 23408 170000 23464
rect 169600 21056 170000 21112
rect 0 20160 400 20216
rect 169600 18704 170000 18760
rect 0 16576 400 16632
rect 169600 16352 170000 16408
rect 169600 14000 170000 14056
rect 0 12992 400 13048
rect 169600 11648 170000 11704
rect 0 9408 400 9464
rect 169600 9296 170000 9352
rect 169600 6944 170000 7000
rect 0 5824 400 5880
rect 169600 4592 170000 4648
rect 0 2240 400 2296
rect 169600 2240 170000 2296
<< obsm3 >>
rect 9 77590 169600 78414
rect 430 77474 169570 77590
rect 9 75238 169600 77474
rect 9 75122 169570 75238
rect 9 74006 169600 75122
rect 430 73890 169600 74006
rect 9 72886 169600 73890
rect 9 72770 169570 72886
rect 9 70534 169600 72770
rect 9 70422 169570 70534
rect 430 70418 169570 70422
rect 430 70306 169600 70418
rect 9 68182 169600 70306
rect 9 68066 169570 68182
rect 9 66838 169600 68066
rect 430 66722 169600 66838
rect 9 65830 169600 66722
rect 9 65714 169570 65830
rect 9 63478 169600 65714
rect 9 63362 169570 63478
rect 9 63254 169600 63362
rect 430 63138 169600 63254
rect 9 61126 169600 63138
rect 9 61010 169570 61126
rect 9 59670 169600 61010
rect 430 59554 169600 59670
rect 9 58774 169600 59554
rect 9 58658 169570 58774
rect 9 56422 169600 58658
rect 9 56306 169570 56422
rect 9 56086 169600 56306
rect 430 55970 169600 56086
rect 9 54070 169600 55970
rect 9 53954 169570 54070
rect 9 52502 169600 53954
rect 430 52386 169600 52502
rect 9 51718 169600 52386
rect 9 51602 169570 51718
rect 9 49366 169600 51602
rect 9 49250 169570 49366
rect 9 48918 169600 49250
rect 430 48802 169600 48918
rect 9 47014 169600 48802
rect 9 46898 169570 47014
rect 9 45334 169600 46898
rect 430 45218 169600 45334
rect 9 44662 169600 45218
rect 9 44546 169570 44662
rect 9 42310 169600 44546
rect 9 42194 169570 42310
rect 9 41750 169600 42194
rect 430 41634 169600 41750
rect 9 39958 169600 41634
rect 9 39842 169570 39958
rect 9 38166 169600 39842
rect 430 38050 169600 38166
rect 9 37606 169600 38050
rect 9 37490 169570 37606
rect 9 35254 169600 37490
rect 9 35138 169570 35254
rect 9 34582 169600 35138
rect 430 34466 169600 34582
rect 9 32902 169600 34466
rect 9 32786 169570 32902
rect 9 30998 169600 32786
rect 430 30882 169600 30998
rect 9 30550 169600 30882
rect 9 30434 169570 30550
rect 9 28198 169600 30434
rect 9 28082 169570 28198
rect 9 27414 169600 28082
rect 430 27298 169600 27414
rect 9 25846 169600 27298
rect 9 25730 169570 25846
rect 9 23830 169600 25730
rect 430 23714 169600 23830
rect 9 23494 169600 23714
rect 9 23378 169570 23494
rect 9 21142 169600 23378
rect 9 21026 169570 21142
rect 9 20246 169600 21026
rect 430 20130 169600 20246
rect 9 18790 169600 20130
rect 9 18674 169570 18790
rect 9 16662 169600 18674
rect 430 16546 169600 16662
rect 9 16438 169600 16546
rect 9 16322 169570 16438
rect 9 14086 169600 16322
rect 9 13970 169570 14086
rect 9 13078 169600 13970
rect 430 12962 169600 13078
rect 9 11734 169600 12962
rect 9 11618 169570 11734
rect 9 9494 169600 11618
rect 430 9382 169600 9494
rect 430 9378 169570 9382
rect 9 9266 169570 9378
rect 9 7030 169600 9266
rect 9 6914 169570 7030
rect 9 5910 169600 6914
rect 430 5794 169600 5910
rect 9 4678 169600 5794
rect 9 4562 169570 4678
rect 9 2326 169600 4562
rect 430 2210 169570 2326
rect 9 350 169600 2210
<< metal4 >>
rect 2224 1538 2384 78430
rect 9904 1538 10064 78430
rect 17584 1538 17744 78430
rect 25264 1538 25424 78430
rect 32944 1538 33104 78430
rect 40624 1538 40784 78430
rect 48304 1538 48464 78430
rect 55984 1538 56144 78430
rect 63664 1538 63824 78430
rect 71344 1538 71504 78430
rect 79024 1538 79184 78430
rect 86704 1538 86864 78430
rect 94384 1538 94544 78430
rect 102064 1538 102224 78430
rect 109744 1538 109904 78430
rect 117424 1538 117584 78430
rect 125104 1538 125264 78430
rect 132784 1538 132944 78430
rect 140464 1538 140624 78430
rect 148144 1538 148304 78430
rect 155824 1538 155984 78430
rect 163504 1538 163664 78430
<< obsm4 >>
rect 6846 1508 9874 78223
rect 10094 1508 17554 78223
rect 17774 1508 25234 78223
rect 25454 1508 32914 78223
rect 33134 1508 40594 78223
rect 40814 1508 48274 78223
rect 48494 1508 55954 78223
rect 56174 1508 63634 78223
rect 63854 1508 71314 78223
rect 71534 1508 78994 78223
rect 79214 1508 86674 78223
rect 86894 1508 94354 78223
rect 94574 1508 102034 78223
rect 102254 1508 109714 78223
rect 109934 1508 117394 78223
rect 117614 1508 125074 78223
rect 125294 1508 132754 78223
rect 132974 1508 140434 78223
rect 140654 1508 144186 78223
rect 6846 625 144186 1508
<< labels >>
rlabel metal3 s 0 9408 400 9464 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 45248 400 45304 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 0 48832 400 48888 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 0 52416 400 52472 6 custom_settings[12]
port 4 nsew signal input
rlabel metal3 s 0 56000 400 56056 6 custom_settings[13]
port 5 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 custom_settings[14]
port 6 nsew signal input
rlabel metal3 s 0 63168 400 63224 6 custom_settings[15]
port 7 nsew signal input
rlabel metal3 s 0 66752 400 66808 6 custom_settings[16]
port 8 nsew signal input
rlabel metal3 s 0 70336 400 70392 6 custom_settings[17]
port 9 nsew signal input
rlabel metal3 s 0 73920 400 73976 6 custom_settings[18]
port 10 nsew signal input
rlabel metal3 s 0 77504 400 77560 6 custom_settings[19]
port 11 nsew signal input
rlabel metal3 s 0 12992 400 13048 6 custom_settings[1]
port 12 nsew signal input
rlabel metal3 s 0 16576 400 16632 6 custom_settings[2]
port 13 nsew signal input
rlabel metal3 s 0 20160 400 20216 6 custom_settings[3]
port 14 nsew signal input
rlabel metal3 s 0 23744 400 23800 6 custom_settings[4]
port 15 nsew signal input
rlabel metal3 s 0 27328 400 27384 6 custom_settings[5]
port 16 nsew signal input
rlabel metal3 s 0 30912 400 30968 6 custom_settings[6]
port 17 nsew signal input
rlabel metal3 s 0 34496 400 34552 6 custom_settings[7]
port 18 nsew signal input
rlabel metal3 s 0 38080 400 38136 6 custom_settings[8]
port 19 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 custom_settings[9]
port 20 nsew signal input
rlabel metal2 s 1232 0 1288 400 6 io_in[0]
port 21 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 io_in[10]
port 22 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 io_in[11]
port 23 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 io_in[12]
port 24 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 io_in[13]
port 25 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 io_in[14]
port 26 nsew signal input
rlabel metal2 s 39872 0 39928 400 6 io_in[15]
port 27 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 io_in[16]
port 28 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 io_in[17]
port 29 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 io_in[18]
port 30 nsew signal input
rlabel metal2 s 50176 0 50232 400 6 io_in[19]
port 31 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 io_in[1]
port 32 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 io_in[20]
port 33 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 io_in[21]
port 34 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 io_in[22]
port 35 nsew signal input
rlabel metal2 s 60480 0 60536 400 6 io_in[23]
port 36 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 io_in[24]
port 37 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 io_in[25]
port 38 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 io_in[26]
port 39 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 io_in[27]
port 40 nsew signal input
rlabel metal2 s 73360 0 73416 400 6 io_in[28]
port 41 nsew signal input
rlabel metal2 s 75936 0 75992 400 6 io_in[29]
port 42 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 io_in[2]
port 43 nsew signal input
rlabel metal2 s 78512 0 78568 400 6 io_in[30]
port 44 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 io_in[31]
port 45 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 io_in[32]
port 46 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 io_in[3]
port 47 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 io_in[4]
port 48 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 io_in[5]
port 49 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 io_in[6]
port 50 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 io_in[7]
port 51 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 io_in[8]
port 52 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 io_in[9]
port 53 nsew signal input
rlabel metal3 s 169600 2240 170000 2296 6 io_oeb[0]
port 54 nsew signal output
rlabel metal3 s 169600 25760 170000 25816 6 io_oeb[10]
port 55 nsew signal output
rlabel metal3 s 169600 28112 170000 28168 6 io_oeb[11]
port 56 nsew signal output
rlabel metal3 s 169600 30464 170000 30520 6 io_oeb[12]
port 57 nsew signal output
rlabel metal3 s 169600 32816 170000 32872 6 io_oeb[13]
port 58 nsew signal output
rlabel metal3 s 169600 35168 170000 35224 6 io_oeb[14]
port 59 nsew signal output
rlabel metal3 s 169600 37520 170000 37576 6 io_oeb[15]
port 60 nsew signal output
rlabel metal3 s 169600 39872 170000 39928 6 io_oeb[16]
port 61 nsew signal output
rlabel metal3 s 169600 42224 170000 42280 6 io_oeb[17]
port 62 nsew signal output
rlabel metal3 s 169600 44576 170000 44632 6 io_oeb[18]
port 63 nsew signal output
rlabel metal3 s 169600 46928 170000 46984 6 io_oeb[19]
port 64 nsew signal output
rlabel metal3 s 169600 4592 170000 4648 6 io_oeb[1]
port 65 nsew signal output
rlabel metal3 s 169600 49280 170000 49336 6 io_oeb[20]
port 66 nsew signal output
rlabel metal3 s 169600 51632 170000 51688 6 io_oeb[21]
port 67 nsew signal output
rlabel metal3 s 169600 53984 170000 54040 6 io_oeb[22]
port 68 nsew signal output
rlabel metal3 s 169600 56336 170000 56392 6 io_oeb[23]
port 69 nsew signal output
rlabel metal3 s 169600 58688 170000 58744 6 io_oeb[24]
port 70 nsew signal output
rlabel metal3 s 169600 61040 170000 61096 6 io_oeb[25]
port 71 nsew signal output
rlabel metal3 s 169600 63392 170000 63448 6 io_oeb[26]
port 72 nsew signal output
rlabel metal3 s 169600 65744 170000 65800 6 io_oeb[27]
port 73 nsew signal output
rlabel metal3 s 169600 68096 170000 68152 6 io_oeb[28]
port 74 nsew signal output
rlabel metal3 s 169600 70448 170000 70504 6 io_oeb[29]
port 75 nsew signal output
rlabel metal3 s 169600 6944 170000 7000 6 io_oeb[2]
port 76 nsew signal output
rlabel metal3 s 169600 72800 170000 72856 6 io_oeb[30]
port 77 nsew signal output
rlabel metal3 s 169600 75152 170000 75208 6 io_oeb[31]
port 78 nsew signal output
rlabel metal3 s 169600 77504 170000 77560 6 io_oeb[32]
port 79 nsew signal output
rlabel metal3 s 169600 9296 170000 9352 6 io_oeb[3]
port 80 nsew signal output
rlabel metal3 s 169600 11648 170000 11704 6 io_oeb[4]
port 81 nsew signal output
rlabel metal3 s 169600 14000 170000 14056 6 io_oeb[5]
port 82 nsew signal output
rlabel metal3 s 169600 16352 170000 16408 6 io_oeb[6]
port 83 nsew signal output
rlabel metal3 s 169600 18704 170000 18760 6 io_oeb[7]
port 84 nsew signal output
rlabel metal3 s 169600 21056 170000 21112 6 io_oeb[8]
port 85 nsew signal output
rlabel metal3 s 169600 23408 170000 23464 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 86240 0 86296 400 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 112000 0 112056 400 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 114576 0 114632 400 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 117152 0 117208 400 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 119728 0 119784 400 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 122304 0 122360 400 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 124880 0 124936 400 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 127456 0 127512 400 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 130032 0 130088 400 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 132608 0 132664 400 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 135184 0 135240 400 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 88816 0 88872 400 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 137760 0 137816 400 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 140336 0 140392 400 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 142912 0 142968 400 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 145488 0 145544 400 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 148064 0 148120 400 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 150640 0 150696 400 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 153216 0 153272 400 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 155792 0 155848 400 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 158368 0 158424 400 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 160944 0 161000 400 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 91392 0 91448 400 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 163520 0 163576 400 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 166096 0 166152 400 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 168672 0 168728 400 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 93968 0 94024 400 6 io_out[3]
port 113 nsew signal output
rlabel metal2 s 96544 0 96600 400 6 io_out[4]
port 114 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 io_out[5]
port 115 nsew signal output
rlabel metal2 s 101696 0 101752 400 6 io_out[6]
port 116 nsew signal output
rlabel metal2 s 104272 0 104328 400 6 io_out[7]
port 117 nsew signal output
rlabel metal2 s 106848 0 106904 400 6 io_out[8]
port 118 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 io_out[9]
port 119 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 rst_n
port 120 nsew signal input
rlabel metal4 s 2224 1538 2384 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 78430 6 vdd
port 121 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 78430 6 vss
port 122 nsew ground bidirectional
rlabel metal3 s 0 2240 400 2296 6 wb_clk_i
port 123 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 170000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 33973146
string GDS_FILE /home/lucah/gfmpw1-multi/openlane/wrapped_pdp11/runs/25_08_05_14_48/results/signoff/wrapped_pdp11.magic.gds
string GDS_START 315406
<< end >>

