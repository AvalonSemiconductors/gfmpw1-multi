magic
tech gf180mcuD
magscale 1 5
timestamp 1702480270
<< obsm1 >>
rect 672 1359 74312 68305
<< metal2 >>
rect 5152 69600 5208 70000
rect 5488 69600 5544 70000
rect 5824 69600 5880 70000
rect 6160 69600 6216 70000
rect 6496 69600 6552 70000
rect 6832 69600 6888 70000
rect 7168 69600 7224 70000
rect 7504 69600 7560 70000
rect 7840 69600 7896 70000
rect 8176 69600 8232 70000
rect 8512 69600 8568 70000
rect 8848 69600 8904 70000
rect 9184 69600 9240 70000
rect 9520 69600 9576 70000
rect 9856 69600 9912 70000
rect 10192 69600 10248 70000
rect 10528 69600 10584 70000
rect 10864 69600 10920 70000
rect 11200 69600 11256 70000
rect 11536 69600 11592 70000
rect 11872 69600 11928 70000
rect 12208 69600 12264 70000
rect 12544 69600 12600 70000
rect 12880 69600 12936 70000
rect 13216 69600 13272 70000
rect 13552 69600 13608 70000
rect 13888 69600 13944 70000
rect 14224 69600 14280 70000
rect 14560 69600 14616 70000
rect 14896 69600 14952 70000
rect 15232 69600 15288 70000
rect 15568 69600 15624 70000
rect 15904 69600 15960 70000
rect 16240 69600 16296 70000
rect 16576 69600 16632 70000
rect 16912 69600 16968 70000
rect 17248 69600 17304 70000
rect 17584 69600 17640 70000
rect 17920 69600 17976 70000
rect 18256 69600 18312 70000
rect 18592 69600 18648 70000
rect 18928 69600 18984 70000
rect 19264 69600 19320 70000
rect 19600 69600 19656 70000
rect 19936 69600 19992 70000
rect 20272 69600 20328 70000
rect 20608 69600 20664 70000
rect 20944 69600 21000 70000
rect 21280 69600 21336 70000
rect 21616 69600 21672 70000
rect 21952 69600 22008 70000
rect 22288 69600 22344 70000
rect 22624 69600 22680 70000
rect 22960 69600 23016 70000
rect 23296 69600 23352 70000
rect 23632 69600 23688 70000
rect 23968 69600 24024 70000
rect 24304 69600 24360 70000
rect 24640 69600 24696 70000
rect 24976 69600 25032 70000
rect 25312 69600 25368 70000
rect 25648 69600 25704 70000
rect 25984 69600 26040 70000
rect 26320 69600 26376 70000
rect 26656 69600 26712 70000
rect 26992 69600 27048 70000
rect 27328 69600 27384 70000
rect 27664 69600 27720 70000
rect 28000 69600 28056 70000
rect 28336 69600 28392 70000
rect 28672 69600 28728 70000
rect 29008 69600 29064 70000
rect 29344 69600 29400 70000
rect 29680 69600 29736 70000
rect 30016 69600 30072 70000
rect 30352 69600 30408 70000
rect 30688 69600 30744 70000
rect 31024 69600 31080 70000
rect 31360 69600 31416 70000
rect 31696 69600 31752 70000
rect 32032 69600 32088 70000
rect 32368 69600 32424 70000
rect 32704 69600 32760 70000
rect 33040 69600 33096 70000
rect 33376 69600 33432 70000
rect 33712 69600 33768 70000
rect 34048 69600 34104 70000
rect 34384 69600 34440 70000
rect 34720 69600 34776 70000
rect 35056 69600 35112 70000
rect 35392 69600 35448 70000
rect 35728 69600 35784 70000
rect 36064 69600 36120 70000
rect 36400 69600 36456 70000
rect 36736 69600 36792 70000
rect 37072 69600 37128 70000
rect 37408 69600 37464 70000
rect 37744 69600 37800 70000
rect 38080 69600 38136 70000
rect 38416 69600 38472 70000
rect 38752 69600 38808 70000
rect 39088 69600 39144 70000
rect 39424 69600 39480 70000
rect 39760 69600 39816 70000
rect 40096 69600 40152 70000
rect 40432 69600 40488 70000
rect 40768 69600 40824 70000
rect 41104 69600 41160 70000
rect 41440 69600 41496 70000
rect 41776 69600 41832 70000
rect 42112 69600 42168 70000
rect 42448 69600 42504 70000
rect 42784 69600 42840 70000
rect 43120 69600 43176 70000
rect 43456 69600 43512 70000
rect 43792 69600 43848 70000
rect 44128 69600 44184 70000
rect 44464 69600 44520 70000
rect 44800 69600 44856 70000
rect 45136 69600 45192 70000
rect 45472 69600 45528 70000
rect 45808 69600 45864 70000
rect 46144 69600 46200 70000
rect 46480 69600 46536 70000
rect 46816 69600 46872 70000
rect 47152 69600 47208 70000
rect 47488 69600 47544 70000
rect 47824 69600 47880 70000
rect 48160 69600 48216 70000
rect 48496 69600 48552 70000
rect 48832 69600 48888 70000
rect 49168 69600 49224 70000
rect 49504 69600 49560 70000
rect 49840 69600 49896 70000
rect 50176 69600 50232 70000
rect 50512 69600 50568 70000
rect 50848 69600 50904 70000
rect 51184 69600 51240 70000
rect 51520 69600 51576 70000
rect 51856 69600 51912 70000
rect 52192 69600 52248 70000
rect 52528 69600 52584 70000
rect 52864 69600 52920 70000
rect 53200 69600 53256 70000
rect 53536 69600 53592 70000
rect 53872 69600 53928 70000
rect 54208 69600 54264 70000
rect 54544 69600 54600 70000
rect 54880 69600 54936 70000
rect 55216 69600 55272 70000
rect 55552 69600 55608 70000
rect 55888 69600 55944 70000
rect 56224 69600 56280 70000
rect 56560 69600 56616 70000
rect 56896 69600 56952 70000
rect 57232 69600 57288 70000
rect 57568 69600 57624 70000
rect 57904 69600 57960 70000
rect 58240 69600 58296 70000
rect 58576 69600 58632 70000
rect 58912 69600 58968 70000
rect 59248 69600 59304 70000
rect 59584 69600 59640 70000
rect 59920 69600 59976 70000
rect 60256 69600 60312 70000
rect 60592 69600 60648 70000
rect 60928 69600 60984 70000
rect 61264 69600 61320 70000
rect 61600 69600 61656 70000
rect 61936 69600 61992 70000
rect 62272 69600 62328 70000
rect 62608 69600 62664 70000
rect 62944 69600 63000 70000
rect 63280 69600 63336 70000
rect 63616 69600 63672 70000
rect 63952 69600 64008 70000
rect 64288 69600 64344 70000
rect 64624 69600 64680 70000
rect 64960 69600 65016 70000
rect 65296 69600 65352 70000
rect 65632 69600 65688 70000
rect 65968 69600 66024 70000
rect 66304 69600 66360 70000
rect 66640 69600 66696 70000
rect 66976 69600 67032 70000
rect 67312 69600 67368 70000
rect 67648 69600 67704 70000
rect 67984 69600 68040 70000
rect 68320 69600 68376 70000
rect 68656 69600 68712 70000
rect 68992 69600 69048 70000
rect 69328 69600 69384 70000
rect 69664 69600 69720 70000
rect 2464 0 2520 400
rect 2912 0 2968 400
rect 3360 0 3416 400
rect 3808 0 3864 400
rect 4256 0 4312 400
rect 4704 0 4760 400
rect 5152 0 5208 400
rect 5600 0 5656 400
rect 6048 0 6104 400
rect 6496 0 6552 400
rect 6944 0 7000 400
rect 7392 0 7448 400
rect 7840 0 7896 400
rect 8288 0 8344 400
rect 8736 0 8792 400
rect 9184 0 9240 400
rect 9632 0 9688 400
rect 10080 0 10136 400
rect 10528 0 10584 400
rect 10976 0 11032 400
rect 11424 0 11480 400
rect 11872 0 11928 400
rect 12320 0 12376 400
rect 12768 0 12824 400
rect 13216 0 13272 400
rect 13664 0 13720 400
rect 14112 0 14168 400
rect 14560 0 14616 400
rect 15008 0 15064 400
rect 15456 0 15512 400
rect 15904 0 15960 400
rect 16352 0 16408 400
rect 16800 0 16856 400
rect 17248 0 17304 400
rect 17696 0 17752 400
rect 18144 0 18200 400
rect 18592 0 18648 400
rect 19040 0 19096 400
rect 19488 0 19544 400
rect 19936 0 19992 400
rect 20384 0 20440 400
rect 20832 0 20888 400
rect 21280 0 21336 400
rect 21728 0 21784 400
rect 22176 0 22232 400
rect 22624 0 22680 400
rect 23072 0 23128 400
rect 23520 0 23576 400
rect 23968 0 24024 400
rect 24416 0 24472 400
rect 24864 0 24920 400
rect 25312 0 25368 400
rect 25760 0 25816 400
rect 26208 0 26264 400
rect 26656 0 26712 400
rect 27104 0 27160 400
rect 27552 0 27608 400
rect 28000 0 28056 400
rect 28448 0 28504 400
rect 28896 0 28952 400
rect 29344 0 29400 400
rect 29792 0 29848 400
rect 30240 0 30296 400
rect 30688 0 30744 400
rect 31136 0 31192 400
rect 31584 0 31640 400
rect 32032 0 32088 400
rect 32480 0 32536 400
rect 32928 0 32984 400
rect 33376 0 33432 400
rect 33824 0 33880 400
rect 34272 0 34328 400
rect 34720 0 34776 400
rect 35168 0 35224 400
rect 35616 0 35672 400
rect 36064 0 36120 400
rect 36512 0 36568 400
rect 36960 0 37016 400
rect 37408 0 37464 400
rect 37856 0 37912 400
rect 38304 0 38360 400
rect 38752 0 38808 400
rect 39200 0 39256 400
rect 39648 0 39704 400
rect 40096 0 40152 400
rect 40544 0 40600 400
rect 40992 0 41048 400
rect 41440 0 41496 400
rect 41888 0 41944 400
rect 42336 0 42392 400
rect 42784 0 42840 400
rect 43232 0 43288 400
rect 43680 0 43736 400
rect 44128 0 44184 400
rect 44576 0 44632 400
rect 45024 0 45080 400
rect 45472 0 45528 400
rect 45920 0 45976 400
rect 46368 0 46424 400
rect 46816 0 46872 400
rect 47264 0 47320 400
rect 47712 0 47768 400
rect 48160 0 48216 400
rect 48608 0 48664 400
rect 49056 0 49112 400
rect 49504 0 49560 400
rect 49952 0 50008 400
rect 50400 0 50456 400
rect 50848 0 50904 400
rect 51296 0 51352 400
rect 51744 0 51800 400
rect 52192 0 52248 400
rect 52640 0 52696 400
rect 53088 0 53144 400
rect 53536 0 53592 400
rect 53984 0 54040 400
rect 54432 0 54488 400
rect 54880 0 54936 400
rect 55328 0 55384 400
rect 55776 0 55832 400
rect 56224 0 56280 400
rect 56672 0 56728 400
rect 57120 0 57176 400
rect 57568 0 57624 400
rect 58016 0 58072 400
rect 58464 0 58520 400
rect 58912 0 58968 400
rect 59360 0 59416 400
rect 59808 0 59864 400
rect 60256 0 60312 400
rect 60704 0 60760 400
rect 61152 0 61208 400
rect 61600 0 61656 400
rect 62048 0 62104 400
rect 62496 0 62552 400
rect 62944 0 63000 400
rect 63392 0 63448 400
rect 63840 0 63896 400
rect 64288 0 64344 400
rect 64736 0 64792 400
rect 65184 0 65240 400
rect 65632 0 65688 400
rect 66080 0 66136 400
rect 66528 0 66584 400
rect 66976 0 67032 400
rect 67424 0 67480 400
rect 67872 0 67928 400
rect 68320 0 68376 400
rect 68768 0 68824 400
rect 69216 0 69272 400
rect 69664 0 69720 400
rect 70112 0 70168 400
rect 70560 0 70616 400
rect 71008 0 71064 400
rect 71456 0 71512 400
rect 71904 0 71960 400
rect 72352 0 72408 400
<< obsm2 >>
rect 798 69570 5122 69600
rect 5238 69570 5458 69600
rect 5574 69570 5794 69600
rect 5910 69570 6130 69600
rect 6246 69570 6466 69600
rect 6582 69570 6802 69600
rect 6918 69570 7138 69600
rect 7254 69570 7474 69600
rect 7590 69570 7810 69600
rect 7926 69570 8146 69600
rect 8262 69570 8482 69600
rect 8598 69570 8818 69600
rect 8934 69570 9154 69600
rect 9270 69570 9490 69600
rect 9606 69570 9826 69600
rect 9942 69570 10162 69600
rect 10278 69570 10498 69600
rect 10614 69570 10834 69600
rect 10950 69570 11170 69600
rect 11286 69570 11506 69600
rect 11622 69570 11842 69600
rect 11958 69570 12178 69600
rect 12294 69570 12514 69600
rect 12630 69570 12850 69600
rect 12966 69570 13186 69600
rect 13302 69570 13522 69600
rect 13638 69570 13858 69600
rect 13974 69570 14194 69600
rect 14310 69570 14530 69600
rect 14646 69570 14866 69600
rect 14982 69570 15202 69600
rect 15318 69570 15538 69600
rect 15654 69570 15874 69600
rect 15990 69570 16210 69600
rect 16326 69570 16546 69600
rect 16662 69570 16882 69600
rect 16998 69570 17218 69600
rect 17334 69570 17554 69600
rect 17670 69570 17890 69600
rect 18006 69570 18226 69600
rect 18342 69570 18562 69600
rect 18678 69570 18898 69600
rect 19014 69570 19234 69600
rect 19350 69570 19570 69600
rect 19686 69570 19906 69600
rect 20022 69570 20242 69600
rect 20358 69570 20578 69600
rect 20694 69570 20914 69600
rect 21030 69570 21250 69600
rect 21366 69570 21586 69600
rect 21702 69570 21922 69600
rect 22038 69570 22258 69600
rect 22374 69570 22594 69600
rect 22710 69570 22930 69600
rect 23046 69570 23266 69600
rect 23382 69570 23602 69600
rect 23718 69570 23938 69600
rect 24054 69570 24274 69600
rect 24390 69570 24610 69600
rect 24726 69570 24946 69600
rect 25062 69570 25282 69600
rect 25398 69570 25618 69600
rect 25734 69570 25954 69600
rect 26070 69570 26290 69600
rect 26406 69570 26626 69600
rect 26742 69570 26962 69600
rect 27078 69570 27298 69600
rect 27414 69570 27634 69600
rect 27750 69570 27970 69600
rect 28086 69570 28306 69600
rect 28422 69570 28642 69600
rect 28758 69570 28978 69600
rect 29094 69570 29314 69600
rect 29430 69570 29650 69600
rect 29766 69570 29986 69600
rect 30102 69570 30322 69600
rect 30438 69570 30658 69600
rect 30774 69570 30994 69600
rect 31110 69570 31330 69600
rect 31446 69570 31666 69600
rect 31782 69570 32002 69600
rect 32118 69570 32338 69600
rect 32454 69570 32674 69600
rect 32790 69570 33010 69600
rect 33126 69570 33346 69600
rect 33462 69570 33682 69600
rect 33798 69570 34018 69600
rect 34134 69570 34354 69600
rect 34470 69570 34690 69600
rect 34806 69570 35026 69600
rect 35142 69570 35362 69600
rect 35478 69570 35698 69600
rect 35814 69570 36034 69600
rect 36150 69570 36370 69600
rect 36486 69570 36706 69600
rect 36822 69570 37042 69600
rect 37158 69570 37378 69600
rect 37494 69570 37714 69600
rect 37830 69570 38050 69600
rect 38166 69570 38386 69600
rect 38502 69570 38722 69600
rect 38838 69570 39058 69600
rect 39174 69570 39394 69600
rect 39510 69570 39730 69600
rect 39846 69570 40066 69600
rect 40182 69570 40402 69600
rect 40518 69570 40738 69600
rect 40854 69570 41074 69600
rect 41190 69570 41410 69600
rect 41526 69570 41746 69600
rect 41862 69570 42082 69600
rect 42198 69570 42418 69600
rect 42534 69570 42754 69600
rect 42870 69570 43090 69600
rect 43206 69570 43426 69600
rect 43542 69570 43762 69600
rect 43878 69570 44098 69600
rect 44214 69570 44434 69600
rect 44550 69570 44770 69600
rect 44886 69570 45106 69600
rect 45222 69570 45442 69600
rect 45558 69570 45778 69600
rect 45894 69570 46114 69600
rect 46230 69570 46450 69600
rect 46566 69570 46786 69600
rect 46902 69570 47122 69600
rect 47238 69570 47458 69600
rect 47574 69570 47794 69600
rect 47910 69570 48130 69600
rect 48246 69570 48466 69600
rect 48582 69570 48802 69600
rect 48918 69570 49138 69600
rect 49254 69570 49474 69600
rect 49590 69570 49810 69600
rect 49926 69570 50146 69600
rect 50262 69570 50482 69600
rect 50598 69570 50818 69600
rect 50934 69570 51154 69600
rect 51270 69570 51490 69600
rect 51606 69570 51826 69600
rect 51942 69570 52162 69600
rect 52278 69570 52498 69600
rect 52614 69570 52834 69600
rect 52950 69570 53170 69600
rect 53286 69570 53506 69600
rect 53622 69570 53842 69600
rect 53958 69570 54178 69600
rect 54294 69570 54514 69600
rect 54630 69570 54850 69600
rect 54966 69570 55186 69600
rect 55302 69570 55522 69600
rect 55638 69570 55858 69600
rect 55974 69570 56194 69600
rect 56310 69570 56530 69600
rect 56646 69570 56866 69600
rect 56982 69570 57202 69600
rect 57318 69570 57538 69600
rect 57654 69570 57874 69600
rect 57990 69570 58210 69600
rect 58326 69570 58546 69600
rect 58662 69570 58882 69600
rect 58998 69570 59218 69600
rect 59334 69570 59554 69600
rect 59670 69570 59890 69600
rect 60006 69570 60226 69600
rect 60342 69570 60562 69600
rect 60678 69570 60898 69600
rect 61014 69570 61234 69600
rect 61350 69570 61570 69600
rect 61686 69570 61906 69600
rect 62022 69570 62242 69600
rect 62358 69570 62578 69600
rect 62694 69570 62914 69600
rect 63030 69570 63250 69600
rect 63366 69570 63586 69600
rect 63702 69570 63922 69600
rect 64038 69570 64258 69600
rect 64374 69570 64594 69600
rect 64710 69570 64930 69600
rect 65046 69570 65266 69600
rect 65382 69570 65602 69600
rect 65718 69570 65938 69600
rect 66054 69570 66274 69600
rect 66390 69570 66610 69600
rect 66726 69570 66946 69600
rect 67062 69570 67282 69600
rect 67398 69570 67618 69600
rect 67734 69570 67954 69600
rect 68070 69570 68290 69600
rect 68406 69570 68626 69600
rect 68742 69570 68962 69600
rect 69078 69570 69298 69600
rect 69414 69570 69634 69600
rect 69750 69570 74186 69600
rect 798 430 74186 69570
rect 798 345 2434 430
rect 2550 345 2882 430
rect 2998 345 3330 430
rect 3446 345 3778 430
rect 3894 345 4226 430
rect 4342 345 4674 430
rect 4790 345 5122 430
rect 5238 345 5570 430
rect 5686 345 6018 430
rect 6134 345 6466 430
rect 6582 345 6914 430
rect 7030 345 7362 430
rect 7478 345 7810 430
rect 7926 345 8258 430
rect 8374 345 8706 430
rect 8822 345 9154 430
rect 9270 345 9602 430
rect 9718 345 10050 430
rect 10166 345 10498 430
rect 10614 345 10946 430
rect 11062 345 11394 430
rect 11510 345 11842 430
rect 11958 345 12290 430
rect 12406 345 12738 430
rect 12854 345 13186 430
rect 13302 345 13634 430
rect 13750 345 14082 430
rect 14198 345 14530 430
rect 14646 345 14978 430
rect 15094 345 15426 430
rect 15542 345 15874 430
rect 15990 345 16322 430
rect 16438 345 16770 430
rect 16886 345 17218 430
rect 17334 345 17666 430
rect 17782 345 18114 430
rect 18230 345 18562 430
rect 18678 345 19010 430
rect 19126 345 19458 430
rect 19574 345 19906 430
rect 20022 345 20354 430
rect 20470 345 20802 430
rect 20918 345 21250 430
rect 21366 345 21698 430
rect 21814 345 22146 430
rect 22262 345 22594 430
rect 22710 345 23042 430
rect 23158 345 23490 430
rect 23606 345 23938 430
rect 24054 345 24386 430
rect 24502 345 24834 430
rect 24950 345 25282 430
rect 25398 345 25730 430
rect 25846 345 26178 430
rect 26294 345 26626 430
rect 26742 345 27074 430
rect 27190 345 27522 430
rect 27638 345 27970 430
rect 28086 345 28418 430
rect 28534 345 28866 430
rect 28982 345 29314 430
rect 29430 345 29762 430
rect 29878 345 30210 430
rect 30326 345 30658 430
rect 30774 345 31106 430
rect 31222 345 31554 430
rect 31670 345 32002 430
rect 32118 345 32450 430
rect 32566 345 32898 430
rect 33014 345 33346 430
rect 33462 345 33794 430
rect 33910 345 34242 430
rect 34358 345 34690 430
rect 34806 345 35138 430
rect 35254 345 35586 430
rect 35702 345 36034 430
rect 36150 345 36482 430
rect 36598 345 36930 430
rect 37046 345 37378 430
rect 37494 345 37826 430
rect 37942 345 38274 430
rect 38390 345 38722 430
rect 38838 345 39170 430
rect 39286 345 39618 430
rect 39734 345 40066 430
rect 40182 345 40514 430
rect 40630 345 40962 430
rect 41078 345 41410 430
rect 41526 345 41858 430
rect 41974 345 42306 430
rect 42422 345 42754 430
rect 42870 345 43202 430
rect 43318 345 43650 430
rect 43766 345 44098 430
rect 44214 345 44546 430
rect 44662 345 44994 430
rect 45110 345 45442 430
rect 45558 345 45890 430
rect 46006 345 46338 430
rect 46454 345 46786 430
rect 46902 345 47234 430
rect 47350 345 47682 430
rect 47798 345 48130 430
rect 48246 345 48578 430
rect 48694 345 49026 430
rect 49142 345 49474 430
rect 49590 345 49922 430
rect 50038 345 50370 430
rect 50486 345 50818 430
rect 50934 345 51266 430
rect 51382 345 51714 430
rect 51830 345 52162 430
rect 52278 345 52610 430
rect 52726 345 53058 430
rect 53174 345 53506 430
rect 53622 345 53954 430
rect 54070 345 54402 430
rect 54518 345 54850 430
rect 54966 345 55298 430
rect 55414 345 55746 430
rect 55862 345 56194 430
rect 56310 345 56642 430
rect 56758 345 57090 430
rect 57206 345 57538 430
rect 57654 345 57986 430
rect 58102 345 58434 430
rect 58550 345 58882 430
rect 58998 345 59330 430
rect 59446 345 59778 430
rect 59894 345 60226 430
rect 60342 345 60674 430
rect 60790 345 61122 430
rect 61238 345 61570 430
rect 61686 345 62018 430
rect 62134 345 62466 430
rect 62582 345 62914 430
rect 63030 345 63362 430
rect 63478 345 63810 430
rect 63926 345 64258 430
rect 64374 345 64706 430
rect 64822 345 65154 430
rect 65270 345 65602 430
rect 65718 345 66050 430
rect 66166 345 66498 430
rect 66614 345 66946 430
rect 67062 345 67394 430
rect 67510 345 67842 430
rect 67958 345 68290 430
rect 68406 345 68738 430
rect 68854 345 69186 430
rect 69302 345 69634 430
rect 69750 345 70082 430
rect 70198 345 70530 430
rect 70646 345 70978 430
rect 71094 345 71426 430
rect 71542 345 71874 430
rect 71990 345 72322 430
rect 72438 345 74186 430
<< metal3 >>
rect 74600 66976 75000 67032
rect 74600 66528 75000 66584
rect 74600 66080 75000 66136
rect 74600 65632 75000 65688
rect 74600 65184 75000 65240
rect 74600 64736 75000 64792
rect 0 64288 400 64344
rect 74600 64288 75000 64344
rect 74600 63840 75000 63896
rect 0 63728 400 63784
rect 74600 63392 75000 63448
rect 0 63168 400 63224
rect 74600 62944 75000 63000
rect 0 62608 400 62664
rect 74600 62496 75000 62552
rect 0 62048 400 62104
rect 74600 62048 75000 62104
rect 74600 61600 75000 61656
rect 0 61488 400 61544
rect 74600 61152 75000 61208
rect 0 60928 400 60984
rect 74600 60704 75000 60760
rect 0 60368 400 60424
rect 74600 60256 75000 60312
rect 0 59808 400 59864
rect 74600 59808 75000 59864
rect 74600 59360 75000 59416
rect 0 59248 400 59304
rect 74600 58912 75000 58968
rect 0 58688 400 58744
rect 74600 58464 75000 58520
rect 0 58128 400 58184
rect 74600 58016 75000 58072
rect 0 57568 400 57624
rect 74600 57568 75000 57624
rect 74600 57120 75000 57176
rect 0 57008 400 57064
rect 74600 56672 75000 56728
rect 0 56448 400 56504
rect 74600 56224 75000 56280
rect 0 55888 400 55944
rect 74600 55776 75000 55832
rect 0 55328 400 55384
rect 74600 55328 75000 55384
rect 74600 54880 75000 54936
rect 0 54768 400 54824
rect 74600 54432 75000 54488
rect 0 54208 400 54264
rect 74600 53984 75000 54040
rect 0 53648 400 53704
rect 74600 53536 75000 53592
rect 0 53088 400 53144
rect 74600 53088 75000 53144
rect 74600 52640 75000 52696
rect 0 52528 400 52584
rect 74600 52192 75000 52248
rect 0 51968 400 52024
rect 74600 51744 75000 51800
rect 0 51408 400 51464
rect 74600 51296 75000 51352
rect 0 50848 400 50904
rect 74600 50848 75000 50904
rect 74600 50400 75000 50456
rect 0 50288 400 50344
rect 74600 49952 75000 50008
rect 0 49728 400 49784
rect 74600 49504 75000 49560
rect 0 49168 400 49224
rect 74600 49056 75000 49112
rect 0 48608 400 48664
rect 74600 48608 75000 48664
rect 74600 48160 75000 48216
rect 0 48048 400 48104
rect 74600 47712 75000 47768
rect 0 47488 400 47544
rect 74600 47264 75000 47320
rect 0 46928 400 46984
rect 74600 46816 75000 46872
rect 0 46368 400 46424
rect 74600 46368 75000 46424
rect 74600 45920 75000 45976
rect 0 45808 400 45864
rect 74600 45472 75000 45528
rect 0 45248 400 45304
rect 74600 45024 75000 45080
rect 0 44688 400 44744
rect 74600 44576 75000 44632
rect 0 44128 400 44184
rect 74600 44128 75000 44184
rect 74600 43680 75000 43736
rect 0 43568 400 43624
rect 74600 43232 75000 43288
rect 0 43008 400 43064
rect 74600 42784 75000 42840
rect 0 42448 400 42504
rect 74600 42336 75000 42392
rect 0 41888 400 41944
rect 74600 41888 75000 41944
rect 74600 41440 75000 41496
rect 0 41328 400 41384
rect 74600 40992 75000 41048
rect 0 40768 400 40824
rect 74600 40544 75000 40600
rect 0 40208 400 40264
rect 74600 40096 75000 40152
rect 0 39648 400 39704
rect 74600 39648 75000 39704
rect 74600 39200 75000 39256
rect 0 39088 400 39144
rect 74600 38752 75000 38808
rect 0 38528 400 38584
rect 74600 38304 75000 38360
rect 0 37968 400 38024
rect 74600 37856 75000 37912
rect 0 37408 400 37464
rect 74600 37408 75000 37464
rect 74600 36960 75000 37016
rect 0 36848 400 36904
rect 74600 36512 75000 36568
rect 0 36288 400 36344
rect 74600 36064 75000 36120
rect 0 35728 400 35784
rect 74600 35616 75000 35672
rect 0 35168 400 35224
rect 74600 35168 75000 35224
rect 74600 34720 75000 34776
rect 0 34608 400 34664
rect 74600 34272 75000 34328
rect 0 34048 400 34104
rect 74600 33824 75000 33880
rect 0 33488 400 33544
rect 74600 33376 75000 33432
rect 0 32928 400 32984
rect 74600 32928 75000 32984
rect 74600 32480 75000 32536
rect 0 32368 400 32424
rect 74600 32032 75000 32088
rect 0 31808 400 31864
rect 74600 31584 75000 31640
rect 0 31248 400 31304
rect 74600 31136 75000 31192
rect 0 30688 400 30744
rect 74600 30688 75000 30744
rect 74600 30240 75000 30296
rect 0 30128 400 30184
rect 74600 29792 75000 29848
rect 0 29568 400 29624
rect 74600 29344 75000 29400
rect 0 29008 400 29064
rect 74600 28896 75000 28952
rect 0 28448 400 28504
rect 74600 28448 75000 28504
rect 74600 28000 75000 28056
rect 0 27888 400 27944
rect 74600 27552 75000 27608
rect 0 27328 400 27384
rect 74600 27104 75000 27160
rect 0 26768 400 26824
rect 74600 26656 75000 26712
rect 0 26208 400 26264
rect 74600 26208 75000 26264
rect 74600 25760 75000 25816
rect 0 25648 400 25704
rect 74600 25312 75000 25368
rect 0 25088 400 25144
rect 74600 24864 75000 24920
rect 0 24528 400 24584
rect 74600 24416 75000 24472
rect 0 23968 400 24024
rect 74600 23968 75000 24024
rect 74600 23520 75000 23576
rect 0 23408 400 23464
rect 74600 23072 75000 23128
rect 0 22848 400 22904
rect 74600 22624 75000 22680
rect 0 22288 400 22344
rect 74600 22176 75000 22232
rect 0 21728 400 21784
rect 74600 21728 75000 21784
rect 74600 21280 75000 21336
rect 0 21168 400 21224
rect 74600 20832 75000 20888
rect 0 20608 400 20664
rect 74600 20384 75000 20440
rect 0 20048 400 20104
rect 74600 19936 75000 19992
rect 0 19488 400 19544
rect 74600 19488 75000 19544
rect 74600 19040 75000 19096
rect 0 18928 400 18984
rect 74600 18592 75000 18648
rect 0 18368 400 18424
rect 74600 18144 75000 18200
rect 0 17808 400 17864
rect 74600 17696 75000 17752
rect 0 17248 400 17304
rect 74600 17248 75000 17304
rect 74600 16800 75000 16856
rect 0 16688 400 16744
rect 74600 16352 75000 16408
rect 0 16128 400 16184
rect 74600 15904 75000 15960
rect 0 15568 400 15624
rect 74600 15456 75000 15512
rect 0 15008 400 15064
rect 74600 15008 75000 15064
rect 74600 14560 75000 14616
rect 0 14448 400 14504
rect 74600 14112 75000 14168
rect 0 13888 400 13944
rect 74600 13664 75000 13720
rect 0 13328 400 13384
rect 74600 13216 75000 13272
rect 0 12768 400 12824
rect 74600 12768 75000 12824
rect 74600 12320 75000 12376
rect 0 12208 400 12264
rect 74600 11872 75000 11928
rect 0 11648 400 11704
rect 74600 11424 75000 11480
rect 0 11088 400 11144
rect 74600 10976 75000 11032
rect 0 10528 400 10584
rect 74600 10528 75000 10584
rect 74600 10080 75000 10136
rect 0 9968 400 10024
rect 74600 9632 75000 9688
rect 0 9408 400 9464
rect 74600 9184 75000 9240
rect 0 8848 400 8904
rect 74600 8736 75000 8792
rect 0 8288 400 8344
rect 74600 8288 75000 8344
rect 74600 7840 75000 7896
rect 0 7728 400 7784
rect 74600 7392 75000 7448
rect 0 7168 400 7224
rect 74600 6944 75000 7000
rect 0 6608 400 6664
rect 74600 6496 75000 6552
rect 0 6048 400 6104
rect 74600 6048 75000 6104
rect 74600 5600 75000 5656
rect 0 5488 400 5544
rect 74600 5152 75000 5208
rect 74600 4704 75000 4760
rect 74600 4256 75000 4312
rect 74600 3808 75000 3864
rect 74600 3360 75000 3416
rect 74600 2912 75000 2968
<< obsm3 >>
rect 400 67062 74634 69258
rect 400 66946 74570 67062
rect 400 66614 74634 66946
rect 400 66498 74570 66614
rect 400 66166 74634 66498
rect 400 66050 74570 66166
rect 400 65718 74634 66050
rect 400 65602 74570 65718
rect 400 65270 74634 65602
rect 400 65154 74570 65270
rect 400 64822 74634 65154
rect 400 64706 74570 64822
rect 400 64374 74634 64706
rect 430 64258 74570 64374
rect 400 63926 74634 64258
rect 400 63814 74570 63926
rect 430 63810 74570 63814
rect 430 63698 74634 63810
rect 400 63478 74634 63698
rect 400 63362 74570 63478
rect 400 63254 74634 63362
rect 430 63138 74634 63254
rect 400 63030 74634 63138
rect 400 62914 74570 63030
rect 400 62694 74634 62914
rect 430 62582 74634 62694
rect 430 62578 74570 62582
rect 400 62466 74570 62578
rect 400 62134 74634 62466
rect 430 62018 74570 62134
rect 400 61686 74634 62018
rect 400 61574 74570 61686
rect 430 61570 74570 61574
rect 430 61458 74634 61570
rect 400 61238 74634 61458
rect 400 61122 74570 61238
rect 400 61014 74634 61122
rect 430 60898 74634 61014
rect 400 60790 74634 60898
rect 400 60674 74570 60790
rect 400 60454 74634 60674
rect 430 60342 74634 60454
rect 430 60338 74570 60342
rect 400 60226 74570 60338
rect 400 59894 74634 60226
rect 430 59778 74570 59894
rect 400 59446 74634 59778
rect 400 59334 74570 59446
rect 430 59330 74570 59334
rect 430 59218 74634 59330
rect 400 58998 74634 59218
rect 400 58882 74570 58998
rect 400 58774 74634 58882
rect 430 58658 74634 58774
rect 400 58550 74634 58658
rect 400 58434 74570 58550
rect 400 58214 74634 58434
rect 430 58102 74634 58214
rect 430 58098 74570 58102
rect 400 57986 74570 58098
rect 400 57654 74634 57986
rect 430 57538 74570 57654
rect 400 57206 74634 57538
rect 400 57094 74570 57206
rect 430 57090 74570 57094
rect 430 56978 74634 57090
rect 400 56758 74634 56978
rect 400 56642 74570 56758
rect 400 56534 74634 56642
rect 430 56418 74634 56534
rect 400 56310 74634 56418
rect 400 56194 74570 56310
rect 400 55974 74634 56194
rect 430 55862 74634 55974
rect 430 55858 74570 55862
rect 400 55746 74570 55858
rect 400 55414 74634 55746
rect 430 55298 74570 55414
rect 400 54966 74634 55298
rect 400 54854 74570 54966
rect 430 54850 74570 54854
rect 430 54738 74634 54850
rect 400 54518 74634 54738
rect 400 54402 74570 54518
rect 400 54294 74634 54402
rect 430 54178 74634 54294
rect 400 54070 74634 54178
rect 400 53954 74570 54070
rect 400 53734 74634 53954
rect 430 53622 74634 53734
rect 430 53618 74570 53622
rect 400 53506 74570 53618
rect 400 53174 74634 53506
rect 430 53058 74570 53174
rect 400 52726 74634 53058
rect 400 52614 74570 52726
rect 430 52610 74570 52614
rect 430 52498 74634 52610
rect 400 52278 74634 52498
rect 400 52162 74570 52278
rect 400 52054 74634 52162
rect 430 51938 74634 52054
rect 400 51830 74634 51938
rect 400 51714 74570 51830
rect 400 51494 74634 51714
rect 430 51382 74634 51494
rect 430 51378 74570 51382
rect 400 51266 74570 51378
rect 400 50934 74634 51266
rect 430 50818 74570 50934
rect 400 50486 74634 50818
rect 400 50374 74570 50486
rect 430 50370 74570 50374
rect 430 50258 74634 50370
rect 400 50038 74634 50258
rect 400 49922 74570 50038
rect 400 49814 74634 49922
rect 430 49698 74634 49814
rect 400 49590 74634 49698
rect 400 49474 74570 49590
rect 400 49254 74634 49474
rect 430 49142 74634 49254
rect 430 49138 74570 49142
rect 400 49026 74570 49138
rect 400 48694 74634 49026
rect 430 48578 74570 48694
rect 400 48246 74634 48578
rect 400 48134 74570 48246
rect 430 48130 74570 48134
rect 430 48018 74634 48130
rect 400 47798 74634 48018
rect 400 47682 74570 47798
rect 400 47574 74634 47682
rect 430 47458 74634 47574
rect 400 47350 74634 47458
rect 400 47234 74570 47350
rect 400 47014 74634 47234
rect 430 46902 74634 47014
rect 430 46898 74570 46902
rect 400 46786 74570 46898
rect 400 46454 74634 46786
rect 430 46338 74570 46454
rect 400 46006 74634 46338
rect 400 45894 74570 46006
rect 430 45890 74570 45894
rect 430 45778 74634 45890
rect 400 45558 74634 45778
rect 400 45442 74570 45558
rect 400 45334 74634 45442
rect 430 45218 74634 45334
rect 400 45110 74634 45218
rect 400 44994 74570 45110
rect 400 44774 74634 44994
rect 430 44662 74634 44774
rect 430 44658 74570 44662
rect 400 44546 74570 44658
rect 400 44214 74634 44546
rect 430 44098 74570 44214
rect 400 43766 74634 44098
rect 400 43654 74570 43766
rect 430 43650 74570 43654
rect 430 43538 74634 43650
rect 400 43318 74634 43538
rect 400 43202 74570 43318
rect 400 43094 74634 43202
rect 430 42978 74634 43094
rect 400 42870 74634 42978
rect 400 42754 74570 42870
rect 400 42534 74634 42754
rect 430 42422 74634 42534
rect 430 42418 74570 42422
rect 400 42306 74570 42418
rect 400 41974 74634 42306
rect 430 41858 74570 41974
rect 400 41526 74634 41858
rect 400 41414 74570 41526
rect 430 41410 74570 41414
rect 430 41298 74634 41410
rect 400 41078 74634 41298
rect 400 40962 74570 41078
rect 400 40854 74634 40962
rect 430 40738 74634 40854
rect 400 40630 74634 40738
rect 400 40514 74570 40630
rect 400 40294 74634 40514
rect 430 40182 74634 40294
rect 430 40178 74570 40182
rect 400 40066 74570 40178
rect 400 39734 74634 40066
rect 430 39618 74570 39734
rect 400 39286 74634 39618
rect 400 39174 74570 39286
rect 430 39170 74570 39174
rect 430 39058 74634 39170
rect 400 38838 74634 39058
rect 400 38722 74570 38838
rect 400 38614 74634 38722
rect 430 38498 74634 38614
rect 400 38390 74634 38498
rect 400 38274 74570 38390
rect 400 38054 74634 38274
rect 430 37942 74634 38054
rect 430 37938 74570 37942
rect 400 37826 74570 37938
rect 400 37494 74634 37826
rect 430 37378 74570 37494
rect 400 37046 74634 37378
rect 400 36934 74570 37046
rect 430 36930 74570 36934
rect 430 36818 74634 36930
rect 400 36598 74634 36818
rect 400 36482 74570 36598
rect 400 36374 74634 36482
rect 430 36258 74634 36374
rect 400 36150 74634 36258
rect 400 36034 74570 36150
rect 400 35814 74634 36034
rect 430 35702 74634 35814
rect 430 35698 74570 35702
rect 400 35586 74570 35698
rect 400 35254 74634 35586
rect 430 35138 74570 35254
rect 400 34806 74634 35138
rect 400 34694 74570 34806
rect 430 34690 74570 34694
rect 430 34578 74634 34690
rect 400 34358 74634 34578
rect 400 34242 74570 34358
rect 400 34134 74634 34242
rect 430 34018 74634 34134
rect 400 33910 74634 34018
rect 400 33794 74570 33910
rect 400 33574 74634 33794
rect 430 33462 74634 33574
rect 430 33458 74570 33462
rect 400 33346 74570 33458
rect 400 33014 74634 33346
rect 430 32898 74570 33014
rect 400 32566 74634 32898
rect 400 32454 74570 32566
rect 430 32450 74570 32454
rect 430 32338 74634 32450
rect 400 32118 74634 32338
rect 400 32002 74570 32118
rect 400 31894 74634 32002
rect 430 31778 74634 31894
rect 400 31670 74634 31778
rect 400 31554 74570 31670
rect 400 31334 74634 31554
rect 430 31222 74634 31334
rect 430 31218 74570 31222
rect 400 31106 74570 31218
rect 400 30774 74634 31106
rect 430 30658 74570 30774
rect 400 30326 74634 30658
rect 400 30214 74570 30326
rect 430 30210 74570 30214
rect 430 30098 74634 30210
rect 400 29878 74634 30098
rect 400 29762 74570 29878
rect 400 29654 74634 29762
rect 430 29538 74634 29654
rect 400 29430 74634 29538
rect 400 29314 74570 29430
rect 400 29094 74634 29314
rect 430 28982 74634 29094
rect 430 28978 74570 28982
rect 400 28866 74570 28978
rect 400 28534 74634 28866
rect 430 28418 74570 28534
rect 400 28086 74634 28418
rect 400 27974 74570 28086
rect 430 27970 74570 27974
rect 430 27858 74634 27970
rect 400 27638 74634 27858
rect 400 27522 74570 27638
rect 400 27414 74634 27522
rect 430 27298 74634 27414
rect 400 27190 74634 27298
rect 400 27074 74570 27190
rect 400 26854 74634 27074
rect 430 26742 74634 26854
rect 430 26738 74570 26742
rect 400 26626 74570 26738
rect 400 26294 74634 26626
rect 430 26178 74570 26294
rect 400 25846 74634 26178
rect 400 25734 74570 25846
rect 430 25730 74570 25734
rect 430 25618 74634 25730
rect 400 25398 74634 25618
rect 400 25282 74570 25398
rect 400 25174 74634 25282
rect 430 25058 74634 25174
rect 400 24950 74634 25058
rect 400 24834 74570 24950
rect 400 24614 74634 24834
rect 430 24502 74634 24614
rect 430 24498 74570 24502
rect 400 24386 74570 24498
rect 400 24054 74634 24386
rect 430 23938 74570 24054
rect 400 23606 74634 23938
rect 400 23494 74570 23606
rect 430 23490 74570 23494
rect 430 23378 74634 23490
rect 400 23158 74634 23378
rect 400 23042 74570 23158
rect 400 22934 74634 23042
rect 430 22818 74634 22934
rect 400 22710 74634 22818
rect 400 22594 74570 22710
rect 400 22374 74634 22594
rect 430 22262 74634 22374
rect 430 22258 74570 22262
rect 400 22146 74570 22258
rect 400 21814 74634 22146
rect 430 21698 74570 21814
rect 400 21366 74634 21698
rect 400 21254 74570 21366
rect 430 21250 74570 21254
rect 430 21138 74634 21250
rect 400 20918 74634 21138
rect 400 20802 74570 20918
rect 400 20694 74634 20802
rect 430 20578 74634 20694
rect 400 20470 74634 20578
rect 400 20354 74570 20470
rect 400 20134 74634 20354
rect 430 20022 74634 20134
rect 430 20018 74570 20022
rect 400 19906 74570 20018
rect 400 19574 74634 19906
rect 430 19458 74570 19574
rect 400 19126 74634 19458
rect 400 19014 74570 19126
rect 430 19010 74570 19014
rect 430 18898 74634 19010
rect 400 18678 74634 18898
rect 400 18562 74570 18678
rect 400 18454 74634 18562
rect 430 18338 74634 18454
rect 400 18230 74634 18338
rect 400 18114 74570 18230
rect 400 17894 74634 18114
rect 430 17782 74634 17894
rect 430 17778 74570 17782
rect 400 17666 74570 17778
rect 400 17334 74634 17666
rect 430 17218 74570 17334
rect 400 16886 74634 17218
rect 400 16774 74570 16886
rect 430 16770 74570 16774
rect 430 16658 74634 16770
rect 400 16438 74634 16658
rect 400 16322 74570 16438
rect 400 16214 74634 16322
rect 430 16098 74634 16214
rect 400 15990 74634 16098
rect 400 15874 74570 15990
rect 400 15654 74634 15874
rect 430 15542 74634 15654
rect 430 15538 74570 15542
rect 400 15426 74570 15538
rect 400 15094 74634 15426
rect 430 14978 74570 15094
rect 400 14646 74634 14978
rect 400 14534 74570 14646
rect 430 14530 74570 14534
rect 430 14418 74634 14530
rect 400 14198 74634 14418
rect 400 14082 74570 14198
rect 400 13974 74634 14082
rect 430 13858 74634 13974
rect 400 13750 74634 13858
rect 400 13634 74570 13750
rect 400 13414 74634 13634
rect 430 13302 74634 13414
rect 430 13298 74570 13302
rect 400 13186 74570 13298
rect 400 12854 74634 13186
rect 430 12738 74570 12854
rect 400 12406 74634 12738
rect 400 12294 74570 12406
rect 430 12290 74570 12294
rect 430 12178 74634 12290
rect 400 11958 74634 12178
rect 400 11842 74570 11958
rect 400 11734 74634 11842
rect 430 11618 74634 11734
rect 400 11510 74634 11618
rect 400 11394 74570 11510
rect 400 11174 74634 11394
rect 430 11062 74634 11174
rect 430 11058 74570 11062
rect 400 10946 74570 11058
rect 400 10614 74634 10946
rect 430 10498 74570 10614
rect 400 10166 74634 10498
rect 400 10054 74570 10166
rect 430 10050 74570 10054
rect 430 9938 74634 10050
rect 400 9718 74634 9938
rect 400 9602 74570 9718
rect 400 9494 74634 9602
rect 430 9378 74634 9494
rect 400 9270 74634 9378
rect 400 9154 74570 9270
rect 400 8934 74634 9154
rect 430 8822 74634 8934
rect 430 8818 74570 8822
rect 400 8706 74570 8818
rect 400 8374 74634 8706
rect 430 8258 74570 8374
rect 400 7926 74634 8258
rect 400 7814 74570 7926
rect 430 7810 74570 7814
rect 430 7698 74634 7810
rect 400 7478 74634 7698
rect 400 7362 74570 7478
rect 400 7254 74634 7362
rect 430 7138 74634 7254
rect 400 7030 74634 7138
rect 400 6914 74570 7030
rect 400 6694 74634 6914
rect 430 6582 74634 6694
rect 430 6578 74570 6582
rect 400 6466 74570 6578
rect 400 6134 74634 6466
rect 430 6018 74570 6134
rect 400 5686 74634 6018
rect 400 5574 74570 5686
rect 430 5570 74570 5574
rect 430 5458 74634 5570
rect 400 5238 74634 5458
rect 400 5122 74570 5238
rect 400 4790 74634 5122
rect 400 4674 74570 4790
rect 400 4342 74634 4674
rect 400 4226 74570 4342
rect 400 3894 74634 4226
rect 400 3778 74570 3894
rect 400 3446 74634 3778
rect 400 3330 74570 3446
rect 400 2998 74634 3330
rect 400 2882 74570 2998
rect 400 350 74634 2882
<< metal4 >>
rect 2224 1538 2384 68238
rect 9904 1538 10064 68238
rect 17584 1538 17744 68238
rect 25264 1538 25424 68238
rect 32944 1538 33104 68238
rect 40624 1538 40784 68238
rect 48304 1538 48464 68238
rect 55984 1538 56144 68238
rect 63664 1538 63824 68238
rect 71344 1538 71504 68238
<< obsm4 >>
rect 26278 68268 73850 69263
rect 26278 1508 32914 68268
rect 33134 1508 40594 68268
rect 40814 1508 48274 68268
rect 48494 1508 55954 68268
rect 56174 1508 63634 68268
rect 63854 1508 71314 68268
rect 71534 1508 73850 68268
rect 26278 1073 73850 1508
<< labels >>
rlabel metal2 s 19600 69600 19656 70000 6 ay8913_do[0]
port 1 nsew signal input
rlabel metal2 s 22960 69600 23016 70000 6 ay8913_do[10]
port 2 nsew signal input
rlabel metal2 s 23296 69600 23352 70000 6 ay8913_do[11]
port 3 nsew signal input
rlabel metal2 s 23632 69600 23688 70000 6 ay8913_do[12]
port 4 nsew signal input
rlabel metal2 s 23968 69600 24024 70000 6 ay8913_do[13]
port 5 nsew signal input
rlabel metal2 s 24304 69600 24360 70000 6 ay8913_do[14]
port 6 nsew signal input
rlabel metal2 s 24640 69600 24696 70000 6 ay8913_do[15]
port 7 nsew signal input
rlabel metal2 s 24976 69600 25032 70000 6 ay8913_do[16]
port 8 nsew signal input
rlabel metal2 s 25312 69600 25368 70000 6 ay8913_do[17]
port 9 nsew signal input
rlabel metal2 s 25648 69600 25704 70000 6 ay8913_do[18]
port 10 nsew signal input
rlabel metal2 s 25984 69600 26040 70000 6 ay8913_do[19]
port 11 nsew signal input
rlabel metal2 s 19936 69600 19992 70000 6 ay8913_do[1]
port 12 nsew signal input
rlabel metal2 s 26320 69600 26376 70000 6 ay8913_do[20]
port 13 nsew signal input
rlabel metal2 s 26656 69600 26712 70000 6 ay8913_do[21]
port 14 nsew signal input
rlabel metal2 s 26992 69600 27048 70000 6 ay8913_do[22]
port 15 nsew signal input
rlabel metal2 s 27328 69600 27384 70000 6 ay8913_do[23]
port 16 nsew signal input
rlabel metal2 s 27664 69600 27720 70000 6 ay8913_do[24]
port 17 nsew signal input
rlabel metal2 s 28000 69600 28056 70000 6 ay8913_do[25]
port 18 nsew signal input
rlabel metal2 s 28336 69600 28392 70000 6 ay8913_do[26]
port 19 nsew signal input
rlabel metal2 s 28672 69600 28728 70000 6 ay8913_do[27]
port 20 nsew signal input
rlabel metal2 s 20272 69600 20328 70000 6 ay8913_do[2]
port 21 nsew signal input
rlabel metal2 s 20608 69600 20664 70000 6 ay8913_do[3]
port 22 nsew signal input
rlabel metal2 s 20944 69600 21000 70000 6 ay8913_do[4]
port 23 nsew signal input
rlabel metal2 s 21280 69600 21336 70000 6 ay8913_do[5]
port 24 nsew signal input
rlabel metal2 s 21616 69600 21672 70000 6 ay8913_do[6]
port 25 nsew signal input
rlabel metal2 s 21952 69600 22008 70000 6 ay8913_do[7]
port 26 nsew signal input
rlabel metal2 s 22288 69600 22344 70000 6 ay8913_do[8]
port 27 nsew signal input
rlabel metal2 s 22624 69600 22680 70000 6 ay8913_do[9]
port 28 nsew signal input
rlabel metal3 s 0 63168 400 63224 6 blinker_do[0]
port 29 nsew signal input
rlabel metal3 s 0 63728 400 63784 6 blinker_do[1]
port 30 nsew signal input
rlabel metal3 s 0 64288 400 64344 6 blinker_do[2]
port 31 nsew signal input
rlabel metal3 s 74600 19040 75000 19096 6 custom_settings[0]
port 32 nsew signal output
rlabel metal3 s 74600 23520 75000 23576 6 custom_settings[10]
port 33 nsew signal output
rlabel metal3 s 74600 23968 75000 24024 6 custom_settings[11]
port 34 nsew signal output
rlabel metal3 s 74600 24416 75000 24472 6 custom_settings[12]
port 35 nsew signal output
rlabel metal3 s 74600 24864 75000 24920 6 custom_settings[13]
port 36 nsew signal output
rlabel metal3 s 74600 25312 75000 25368 6 custom_settings[14]
port 37 nsew signal output
rlabel metal3 s 74600 25760 75000 25816 6 custom_settings[15]
port 38 nsew signal output
rlabel metal3 s 74600 26208 75000 26264 6 custom_settings[16]
port 39 nsew signal output
rlabel metal3 s 74600 26656 75000 26712 6 custom_settings[17]
port 40 nsew signal output
rlabel metal3 s 74600 27104 75000 27160 6 custom_settings[18]
port 41 nsew signal output
rlabel metal3 s 74600 27552 75000 27608 6 custom_settings[19]
port 42 nsew signal output
rlabel metal3 s 74600 19488 75000 19544 6 custom_settings[1]
port 43 nsew signal output
rlabel metal3 s 74600 28000 75000 28056 6 custom_settings[20]
port 44 nsew signal output
rlabel metal3 s 74600 28448 75000 28504 6 custom_settings[21]
port 45 nsew signal output
rlabel metal3 s 74600 28896 75000 28952 6 custom_settings[22]
port 46 nsew signal output
rlabel metal3 s 74600 29344 75000 29400 6 custom_settings[23]
port 47 nsew signal output
rlabel metal3 s 74600 29792 75000 29848 6 custom_settings[24]
port 48 nsew signal output
rlabel metal3 s 74600 30240 75000 30296 6 custom_settings[25]
port 49 nsew signal output
rlabel metal3 s 74600 30688 75000 30744 6 custom_settings[26]
port 50 nsew signal output
rlabel metal3 s 74600 31136 75000 31192 6 custom_settings[27]
port 51 nsew signal output
rlabel metal3 s 74600 31584 75000 31640 6 custom_settings[28]
port 52 nsew signal output
rlabel metal3 s 74600 32032 75000 32088 6 custom_settings[29]
port 53 nsew signal output
rlabel metal3 s 74600 19936 75000 19992 6 custom_settings[2]
port 54 nsew signal output
rlabel metal3 s 74600 32480 75000 32536 6 custom_settings[30]
port 55 nsew signal output
rlabel metal3 s 74600 32928 75000 32984 6 custom_settings[31]
port 56 nsew signal output
rlabel metal3 s 74600 20384 75000 20440 6 custom_settings[3]
port 57 nsew signal output
rlabel metal3 s 74600 20832 75000 20888 6 custom_settings[4]
port 58 nsew signal output
rlabel metal3 s 74600 21280 75000 21336 6 custom_settings[5]
port 59 nsew signal output
rlabel metal3 s 74600 21728 75000 21784 6 custom_settings[6]
port 60 nsew signal output
rlabel metal3 s 74600 22176 75000 22232 6 custom_settings[7]
port 61 nsew signal output
rlabel metal3 s 74600 22624 75000 22680 6 custom_settings[8]
port 62 nsew signal output
rlabel metal3 s 74600 23072 75000 23128 6 custom_settings[9]
port 63 nsew signal output
rlabel metal2 s 62944 69600 63000 70000 6 diceroll_do[0]
port 64 nsew signal input
rlabel metal2 s 63280 69600 63336 70000 6 diceroll_do[1]
port 65 nsew signal input
rlabel metal2 s 63616 69600 63672 70000 6 diceroll_do[2]
port 66 nsew signal input
rlabel metal2 s 63952 69600 64008 70000 6 diceroll_do[3]
port 67 nsew signal input
rlabel metal2 s 64288 69600 64344 70000 6 diceroll_do[4]
port 68 nsew signal input
rlabel metal2 s 64624 69600 64680 70000 6 diceroll_do[5]
port 69 nsew signal input
rlabel metal2 s 64960 69600 65016 70000 6 diceroll_do[6]
port 70 nsew signal input
rlabel metal2 s 65296 69600 65352 70000 6 diceroll_do[7]
port 71 nsew signal input
rlabel metal2 s 65632 69600 65688 70000 6 diceroll_do[8]
port 72 nsew signal input
rlabel metal3 s 0 58688 400 58744 6 hellorld_do
port 73 nsew signal input
rlabel metal2 s 5152 69600 5208 70000 6 io_in_0
port 74 nsew signal input
rlabel metal3 s 0 5488 400 5544 6 io_oeb[0]
port 75 nsew signal output
rlabel metal3 s 0 11088 400 11144 6 io_oeb[10]
port 76 nsew signal output
rlabel metal3 s 0 11648 400 11704 6 io_oeb[11]
port 77 nsew signal output
rlabel metal3 s 0 12208 400 12264 6 io_oeb[12]
port 78 nsew signal output
rlabel metal3 s 0 12768 400 12824 6 io_oeb[13]
port 79 nsew signal output
rlabel metal3 s 0 13328 400 13384 6 io_oeb[14]
port 80 nsew signal output
rlabel metal3 s 0 13888 400 13944 6 io_oeb[15]
port 81 nsew signal output
rlabel metal3 s 0 14448 400 14504 6 io_oeb[16]
port 82 nsew signal output
rlabel metal3 s 0 15008 400 15064 6 io_oeb[17]
port 83 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 io_oeb[18]
port 84 nsew signal output
rlabel metal3 s 0 16128 400 16184 6 io_oeb[19]
port 85 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 io_oeb[1]
port 86 nsew signal output
rlabel metal3 s 0 16688 400 16744 6 io_oeb[20]
port 87 nsew signal output
rlabel metal3 s 0 17248 400 17304 6 io_oeb[21]
port 88 nsew signal output
rlabel metal3 s 0 17808 400 17864 6 io_oeb[22]
port 89 nsew signal output
rlabel metal3 s 0 18368 400 18424 6 io_oeb[23]
port 90 nsew signal output
rlabel metal3 s 0 18928 400 18984 6 io_oeb[24]
port 91 nsew signal output
rlabel metal3 s 0 19488 400 19544 6 io_oeb[25]
port 92 nsew signal output
rlabel metal3 s 0 20048 400 20104 6 io_oeb[26]
port 93 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 io_oeb[27]
port 94 nsew signal output
rlabel metal3 s 0 21168 400 21224 6 io_oeb[28]
port 95 nsew signal output
rlabel metal3 s 0 21728 400 21784 6 io_oeb[29]
port 96 nsew signal output
rlabel metal3 s 0 6608 400 6664 6 io_oeb[2]
port 97 nsew signal output
rlabel metal3 s 0 22288 400 22344 6 io_oeb[30]
port 98 nsew signal output
rlabel metal3 s 0 22848 400 22904 6 io_oeb[31]
port 99 nsew signal output
rlabel metal3 s 0 23408 400 23464 6 io_oeb[32]
port 100 nsew signal output
rlabel metal3 s 0 23968 400 24024 6 io_oeb[33]
port 101 nsew signal output
rlabel metal3 s 0 24528 400 24584 6 io_oeb[34]
port 102 nsew signal output
rlabel metal3 s 0 25088 400 25144 6 io_oeb[35]
port 103 nsew signal output
rlabel metal3 s 0 25648 400 25704 6 io_oeb[36]
port 104 nsew signal output
rlabel metal3 s 0 26208 400 26264 6 io_oeb[37]
port 105 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 io_oeb[3]
port 106 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 io_oeb[4]
port 107 nsew signal output
rlabel metal3 s 0 8288 400 8344 6 io_oeb[5]
port 108 nsew signal output
rlabel metal3 s 0 8848 400 8904 6 io_oeb[6]
port 109 nsew signal output
rlabel metal3 s 0 9408 400 9464 6 io_oeb[7]
port 110 nsew signal output
rlabel metal3 s 0 9968 400 10024 6 io_oeb[8]
port 111 nsew signal output
rlabel metal3 s 0 10528 400 10584 6 io_oeb[9]
port 112 nsew signal output
rlabel metal2 s 5488 69600 5544 70000 6 io_out[0]
port 113 nsew signal output
rlabel metal2 s 8848 69600 8904 70000 6 io_out[10]
port 114 nsew signal output
rlabel metal2 s 9184 69600 9240 70000 6 io_out[11]
port 115 nsew signal output
rlabel metal2 s 9520 69600 9576 70000 6 io_out[12]
port 116 nsew signal output
rlabel metal2 s 9856 69600 9912 70000 6 io_out[13]
port 117 nsew signal output
rlabel metal2 s 10192 69600 10248 70000 6 io_out[14]
port 118 nsew signal output
rlabel metal2 s 10528 69600 10584 70000 6 io_out[15]
port 119 nsew signal output
rlabel metal2 s 10864 69600 10920 70000 6 io_out[16]
port 120 nsew signal output
rlabel metal2 s 11200 69600 11256 70000 6 io_out[17]
port 121 nsew signal output
rlabel metal2 s 11536 69600 11592 70000 6 io_out[18]
port 122 nsew signal output
rlabel metal2 s 11872 69600 11928 70000 6 io_out[19]
port 123 nsew signal output
rlabel metal2 s 5824 69600 5880 70000 6 io_out[1]
port 124 nsew signal output
rlabel metal2 s 12208 69600 12264 70000 6 io_out[20]
port 125 nsew signal output
rlabel metal2 s 12544 69600 12600 70000 6 io_out[21]
port 126 nsew signal output
rlabel metal2 s 12880 69600 12936 70000 6 io_out[22]
port 127 nsew signal output
rlabel metal2 s 13216 69600 13272 70000 6 io_out[23]
port 128 nsew signal output
rlabel metal2 s 13552 69600 13608 70000 6 io_out[24]
port 129 nsew signal output
rlabel metal2 s 13888 69600 13944 70000 6 io_out[25]
port 130 nsew signal output
rlabel metal2 s 14224 69600 14280 70000 6 io_out[26]
port 131 nsew signal output
rlabel metal2 s 14560 69600 14616 70000 6 io_out[27]
port 132 nsew signal output
rlabel metal2 s 14896 69600 14952 70000 6 io_out[28]
port 133 nsew signal output
rlabel metal2 s 15232 69600 15288 70000 6 io_out[29]
port 134 nsew signal output
rlabel metal2 s 6160 69600 6216 70000 6 io_out[2]
port 135 nsew signal output
rlabel metal2 s 15568 69600 15624 70000 6 io_out[30]
port 136 nsew signal output
rlabel metal2 s 15904 69600 15960 70000 6 io_out[31]
port 137 nsew signal output
rlabel metal2 s 16240 69600 16296 70000 6 io_out[32]
port 138 nsew signal output
rlabel metal2 s 16576 69600 16632 70000 6 io_out[33]
port 139 nsew signal output
rlabel metal2 s 16912 69600 16968 70000 6 io_out[34]
port 140 nsew signal output
rlabel metal2 s 17248 69600 17304 70000 6 io_out[35]
port 141 nsew signal output
rlabel metal2 s 17584 69600 17640 70000 6 io_out[36]
port 142 nsew signal output
rlabel metal2 s 17920 69600 17976 70000 6 io_out[37]
port 143 nsew signal output
rlabel metal2 s 6496 69600 6552 70000 6 io_out[3]
port 144 nsew signal output
rlabel metal2 s 6832 69600 6888 70000 6 io_out[4]
port 145 nsew signal output
rlabel metal2 s 7168 69600 7224 70000 6 io_out[5]
port 146 nsew signal output
rlabel metal2 s 7504 69600 7560 70000 6 io_out[6]
port 147 nsew signal output
rlabel metal2 s 7840 69600 7896 70000 6 io_out[7]
port 148 nsew signal output
rlabel metal2 s 8176 69600 8232 70000 6 io_out[8]
port 149 nsew signal output
rlabel metal2 s 8512 69600 8568 70000 6 io_out[9]
port 150 nsew signal output
rlabel metal2 s 18256 69600 18312 70000 6 irq[0]
port 151 nsew signal output
rlabel metal2 s 18592 69600 18648 70000 6 irq[1]
port 152 nsew signal output
rlabel metal2 s 18928 69600 18984 70000 6 irq[2]
port 153 nsew signal output
rlabel metal3 s 0 40768 400 40824 6 mc14500_do[0]
port 154 nsew signal input
rlabel metal3 s 0 46368 400 46424 6 mc14500_do[10]
port 155 nsew signal input
rlabel metal3 s 0 46928 400 46984 6 mc14500_do[11]
port 156 nsew signal input
rlabel metal3 s 0 47488 400 47544 6 mc14500_do[12]
port 157 nsew signal input
rlabel metal3 s 0 48048 400 48104 6 mc14500_do[13]
port 158 nsew signal input
rlabel metal3 s 0 48608 400 48664 6 mc14500_do[14]
port 159 nsew signal input
rlabel metal3 s 0 49168 400 49224 6 mc14500_do[15]
port 160 nsew signal input
rlabel metal3 s 0 49728 400 49784 6 mc14500_do[16]
port 161 nsew signal input
rlabel metal3 s 0 50288 400 50344 6 mc14500_do[17]
port 162 nsew signal input
rlabel metal3 s 0 50848 400 50904 6 mc14500_do[18]
port 163 nsew signal input
rlabel metal3 s 0 51408 400 51464 6 mc14500_do[19]
port 164 nsew signal input
rlabel metal3 s 0 41328 400 41384 6 mc14500_do[1]
port 165 nsew signal input
rlabel metal3 s 0 51968 400 52024 6 mc14500_do[20]
port 166 nsew signal input
rlabel metal3 s 0 52528 400 52584 6 mc14500_do[21]
port 167 nsew signal input
rlabel metal3 s 0 53088 400 53144 6 mc14500_do[22]
port 168 nsew signal input
rlabel metal3 s 0 53648 400 53704 6 mc14500_do[23]
port 169 nsew signal input
rlabel metal3 s 0 54208 400 54264 6 mc14500_do[24]
port 170 nsew signal input
rlabel metal3 s 0 54768 400 54824 6 mc14500_do[25]
port 171 nsew signal input
rlabel metal3 s 0 55328 400 55384 6 mc14500_do[26]
port 172 nsew signal input
rlabel metal3 s 0 55888 400 55944 6 mc14500_do[27]
port 173 nsew signal input
rlabel metal3 s 0 56448 400 56504 6 mc14500_do[28]
port 174 nsew signal input
rlabel metal3 s 0 57008 400 57064 6 mc14500_do[29]
port 175 nsew signal input
rlabel metal3 s 0 41888 400 41944 6 mc14500_do[2]
port 176 nsew signal input
rlabel metal3 s 0 57568 400 57624 6 mc14500_do[30]
port 177 nsew signal input
rlabel metal3 s 0 42448 400 42504 6 mc14500_do[3]
port 178 nsew signal input
rlabel metal3 s 0 43008 400 43064 6 mc14500_do[4]
port 179 nsew signal input
rlabel metal3 s 0 43568 400 43624 6 mc14500_do[5]
port 180 nsew signal input
rlabel metal3 s 0 44128 400 44184 6 mc14500_do[6]
port 181 nsew signal input
rlabel metal3 s 0 44688 400 44744 6 mc14500_do[7]
port 182 nsew signal input
rlabel metal3 s 0 45248 400 45304 6 mc14500_do[8]
port 183 nsew signal input
rlabel metal3 s 0 45808 400 45864 6 mc14500_do[9]
port 184 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 mc14500_sram_addr[0]
port 185 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 mc14500_sram_addr[1]
port 186 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 mc14500_sram_addr[2]
port 187 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 mc14500_sram_addr[3]
port 188 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 mc14500_sram_addr[4]
port 189 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 mc14500_sram_addr[5]
port 190 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 mc14500_sram_gwe
port 191 nsew signal input
rlabel metal2 s 68768 0 68824 400 6 mc14500_sram_in[0]
port 192 nsew signal input
rlabel metal2 s 69216 0 69272 400 6 mc14500_sram_in[1]
port 193 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 mc14500_sram_in[2]
port 194 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 mc14500_sram_in[3]
port 195 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 mc14500_sram_in[4]
port 196 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 mc14500_sram_in[5]
port 197 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 mc14500_sram_in[6]
port 198 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 mc14500_sram_in[7]
port 199 nsew signal input
rlabel metal2 s 29008 69600 29064 70000 6 pdp11_do[0]
port 200 nsew signal input
rlabel metal2 s 35728 69600 35784 70000 6 pdp11_do[10]
port 201 nsew signal input
rlabel metal2 s 36400 69600 36456 70000 6 pdp11_do[11]
port 202 nsew signal input
rlabel metal2 s 37072 69600 37128 70000 6 pdp11_do[12]
port 203 nsew signal input
rlabel metal2 s 37744 69600 37800 70000 6 pdp11_do[13]
port 204 nsew signal input
rlabel metal2 s 38416 69600 38472 70000 6 pdp11_do[14]
port 205 nsew signal input
rlabel metal2 s 39088 69600 39144 70000 6 pdp11_do[15]
port 206 nsew signal input
rlabel metal2 s 39760 69600 39816 70000 6 pdp11_do[16]
port 207 nsew signal input
rlabel metal2 s 40432 69600 40488 70000 6 pdp11_do[17]
port 208 nsew signal input
rlabel metal2 s 41104 69600 41160 70000 6 pdp11_do[18]
port 209 nsew signal input
rlabel metal2 s 41776 69600 41832 70000 6 pdp11_do[19]
port 210 nsew signal input
rlabel metal2 s 29680 69600 29736 70000 6 pdp11_do[1]
port 211 nsew signal input
rlabel metal2 s 42448 69600 42504 70000 6 pdp11_do[20]
port 212 nsew signal input
rlabel metal2 s 43120 69600 43176 70000 6 pdp11_do[21]
port 213 nsew signal input
rlabel metal2 s 43792 69600 43848 70000 6 pdp11_do[22]
port 214 nsew signal input
rlabel metal2 s 44464 69600 44520 70000 6 pdp11_do[23]
port 215 nsew signal input
rlabel metal2 s 45136 69600 45192 70000 6 pdp11_do[24]
port 216 nsew signal input
rlabel metal2 s 45808 69600 45864 70000 6 pdp11_do[25]
port 217 nsew signal input
rlabel metal2 s 46480 69600 46536 70000 6 pdp11_do[26]
port 218 nsew signal input
rlabel metal2 s 47152 69600 47208 70000 6 pdp11_do[27]
port 219 nsew signal input
rlabel metal2 s 47824 69600 47880 70000 6 pdp11_do[28]
port 220 nsew signal input
rlabel metal2 s 48496 69600 48552 70000 6 pdp11_do[29]
port 221 nsew signal input
rlabel metal2 s 30352 69600 30408 70000 6 pdp11_do[2]
port 222 nsew signal input
rlabel metal2 s 49168 69600 49224 70000 6 pdp11_do[30]
port 223 nsew signal input
rlabel metal2 s 49840 69600 49896 70000 6 pdp11_do[31]
port 224 nsew signal input
rlabel metal2 s 50512 69600 50568 70000 6 pdp11_do[32]
port 225 nsew signal input
rlabel metal2 s 31024 69600 31080 70000 6 pdp11_do[3]
port 226 nsew signal input
rlabel metal2 s 31696 69600 31752 70000 6 pdp11_do[4]
port 227 nsew signal input
rlabel metal2 s 32368 69600 32424 70000 6 pdp11_do[5]
port 228 nsew signal input
rlabel metal2 s 33040 69600 33096 70000 6 pdp11_do[6]
port 229 nsew signal input
rlabel metal2 s 33712 69600 33768 70000 6 pdp11_do[7]
port 230 nsew signal input
rlabel metal2 s 34384 69600 34440 70000 6 pdp11_do[8]
port 231 nsew signal input
rlabel metal2 s 35056 69600 35112 70000 6 pdp11_do[9]
port 232 nsew signal input
rlabel metal2 s 29344 69600 29400 70000 6 pdp11_oeb[0]
port 233 nsew signal input
rlabel metal2 s 36064 69600 36120 70000 6 pdp11_oeb[10]
port 234 nsew signal input
rlabel metal2 s 36736 69600 36792 70000 6 pdp11_oeb[11]
port 235 nsew signal input
rlabel metal2 s 37408 69600 37464 70000 6 pdp11_oeb[12]
port 236 nsew signal input
rlabel metal2 s 38080 69600 38136 70000 6 pdp11_oeb[13]
port 237 nsew signal input
rlabel metal2 s 38752 69600 38808 70000 6 pdp11_oeb[14]
port 238 nsew signal input
rlabel metal2 s 39424 69600 39480 70000 6 pdp11_oeb[15]
port 239 nsew signal input
rlabel metal2 s 40096 69600 40152 70000 6 pdp11_oeb[16]
port 240 nsew signal input
rlabel metal2 s 40768 69600 40824 70000 6 pdp11_oeb[17]
port 241 nsew signal input
rlabel metal2 s 41440 69600 41496 70000 6 pdp11_oeb[18]
port 242 nsew signal input
rlabel metal2 s 42112 69600 42168 70000 6 pdp11_oeb[19]
port 243 nsew signal input
rlabel metal2 s 30016 69600 30072 70000 6 pdp11_oeb[1]
port 244 nsew signal input
rlabel metal2 s 42784 69600 42840 70000 6 pdp11_oeb[20]
port 245 nsew signal input
rlabel metal2 s 43456 69600 43512 70000 6 pdp11_oeb[21]
port 246 nsew signal input
rlabel metal2 s 44128 69600 44184 70000 6 pdp11_oeb[22]
port 247 nsew signal input
rlabel metal2 s 44800 69600 44856 70000 6 pdp11_oeb[23]
port 248 nsew signal input
rlabel metal2 s 45472 69600 45528 70000 6 pdp11_oeb[24]
port 249 nsew signal input
rlabel metal2 s 46144 69600 46200 70000 6 pdp11_oeb[25]
port 250 nsew signal input
rlabel metal2 s 46816 69600 46872 70000 6 pdp11_oeb[26]
port 251 nsew signal input
rlabel metal2 s 47488 69600 47544 70000 6 pdp11_oeb[27]
port 252 nsew signal input
rlabel metal2 s 48160 69600 48216 70000 6 pdp11_oeb[28]
port 253 nsew signal input
rlabel metal2 s 48832 69600 48888 70000 6 pdp11_oeb[29]
port 254 nsew signal input
rlabel metal2 s 30688 69600 30744 70000 6 pdp11_oeb[2]
port 255 nsew signal input
rlabel metal2 s 49504 69600 49560 70000 6 pdp11_oeb[30]
port 256 nsew signal input
rlabel metal2 s 50176 69600 50232 70000 6 pdp11_oeb[31]
port 257 nsew signal input
rlabel metal2 s 50848 69600 50904 70000 6 pdp11_oeb[32]
port 258 nsew signal input
rlabel metal2 s 31360 69600 31416 70000 6 pdp11_oeb[3]
port 259 nsew signal input
rlabel metal2 s 32032 69600 32088 70000 6 pdp11_oeb[4]
port 260 nsew signal input
rlabel metal2 s 32704 69600 32760 70000 6 pdp11_oeb[5]
port 261 nsew signal input
rlabel metal2 s 33376 69600 33432 70000 6 pdp11_oeb[6]
port 262 nsew signal input
rlabel metal2 s 34048 69600 34104 70000 6 pdp11_oeb[7]
port 263 nsew signal input
rlabel metal2 s 34720 69600 34776 70000 6 pdp11_oeb[8]
port 264 nsew signal input
rlabel metal2 s 35392 69600 35448 70000 6 pdp11_oeb[9]
port 265 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 qcpu_do[0]
port 266 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 qcpu_do[10]
port 267 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 qcpu_do[11]
port 268 nsew signal input
rlabel metal2 s 49952 0 50008 400 6 qcpu_do[12]
port 269 nsew signal input
rlabel metal2 s 50400 0 50456 400 6 qcpu_do[13]
port 270 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 qcpu_do[14]
port 271 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 qcpu_do[15]
port 272 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 qcpu_do[16]
port 273 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 qcpu_do[17]
port 274 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 qcpu_do[18]
port 275 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 qcpu_do[19]
port 276 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 qcpu_do[1]
port 277 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 qcpu_do[20]
port 278 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 qcpu_do[21]
port 279 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 qcpu_do[22]
port 280 nsew signal input
rlabel metal2 s 54880 0 54936 400 6 qcpu_do[23]
port 281 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 qcpu_do[24]
port 282 nsew signal input
rlabel metal2 s 55776 0 55832 400 6 qcpu_do[25]
port 283 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 qcpu_do[26]
port 284 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 qcpu_do[27]
port 285 nsew signal input
rlabel metal2 s 57120 0 57176 400 6 qcpu_do[28]
port 286 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 qcpu_do[29]
port 287 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 qcpu_do[2]
port 288 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 qcpu_do[30]
port 289 nsew signal input
rlabel metal2 s 58464 0 58520 400 6 qcpu_do[31]
port 290 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 qcpu_do[32]
port 291 nsew signal input
rlabel metal2 s 45920 0 45976 400 6 qcpu_do[3]
port 292 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 qcpu_do[4]
port 293 nsew signal input
rlabel metal2 s 46816 0 46872 400 6 qcpu_do[5]
port 294 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 qcpu_do[6]
port 295 nsew signal input
rlabel metal2 s 47712 0 47768 400 6 qcpu_do[7]
port 296 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 qcpu_do[8]
port 297 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 qcpu_do[9]
port 298 nsew signal input
rlabel metal3 s 74600 33376 75000 33432 6 qcpu_oeb[0]
port 299 nsew signal input
rlabel metal3 s 74600 37856 75000 37912 6 qcpu_oeb[10]
port 300 nsew signal input
rlabel metal3 s 74600 38304 75000 38360 6 qcpu_oeb[11]
port 301 nsew signal input
rlabel metal3 s 74600 38752 75000 38808 6 qcpu_oeb[12]
port 302 nsew signal input
rlabel metal3 s 74600 39200 75000 39256 6 qcpu_oeb[13]
port 303 nsew signal input
rlabel metal3 s 74600 39648 75000 39704 6 qcpu_oeb[14]
port 304 nsew signal input
rlabel metal3 s 74600 40096 75000 40152 6 qcpu_oeb[15]
port 305 nsew signal input
rlabel metal3 s 74600 40544 75000 40600 6 qcpu_oeb[16]
port 306 nsew signal input
rlabel metal3 s 74600 40992 75000 41048 6 qcpu_oeb[17]
port 307 nsew signal input
rlabel metal3 s 74600 41440 75000 41496 6 qcpu_oeb[18]
port 308 nsew signal input
rlabel metal3 s 74600 41888 75000 41944 6 qcpu_oeb[19]
port 309 nsew signal input
rlabel metal3 s 74600 33824 75000 33880 6 qcpu_oeb[1]
port 310 nsew signal input
rlabel metal3 s 74600 42336 75000 42392 6 qcpu_oeb[20]
port 311 nsew signal input
rlabel metal3 s 74600 42784 75000 42840 6 qcpu_oeb[21]
port 312 nsew signal input
rlabel metal3 s 74600 43232 75000 43288 6 qcpu_oeb[22]
port 313 nsew signal input
rlabel metal3 s 74600 43680 75000 43736 6 qcpu_oeb[23]
port 314 nsew signal input
rlabel metal3 s 74600 44128 75000 44184 6 qcpu_oeb[24]
port 315 nsew signal input
rlabel metal3 s 74600 44576 75000 44632 6 qcpu_oeb[25]
port 316 nsew signal input
rlabel metal3 s 74600 45024 75000 45080 6 qcpu_oeb[26]
port 317 nsew signal input
rlabel metal3 s 74600 45472 75000 45528 6 qcpu_oeb[27]
port 318 nsew signal input
rlabel metal3 s 74600 45920 75000 45976 6 qcpu_oeb[28]
port 319 nsew signal input
rlabel metal3 s 74600 46368 75000 46424 6 qcpu_oeb[29]
port 320 nsew signal input
rlabel metal3 s 74600 34272 75000 34328 6 qcpu_oeb[2]
port 321 nsew signal input
rlabel metal3 s 74600 46816 75000 46872 6 qcpu_oeb[30]
port 322 nsew signal input
rlabel metal3 s 74600 47264 75000 47320 6 qcpu_oeb[31]
port 323 nsew signal input
rlabel metal3 s 74600 47712 75000 47768 6 qcpu_oeb[32]
port 324 nsew signal input
rlabel metal3 s 74600 34720 75000 34776 6 qcpu_oeb[3]
port 325 nsew signal input
rlabel metal3 s 74600 35168 75000 35224 6 qcpu_oeb[4]
port 326 nsew signal input
rlabel metal3 s 74600 35616 75000 35672 6 qcpu_oeb[5]
port 327 nsew signal input
rlabel metal3 s 74600 36064 75000 36120 6 qcpu_oeb[6]
port 328 nsew signal input
rlabel metal3 s 74600 36512 75000 36568 6 qcpu_oeb[7]
port 329 nsew signal input
rlabel metal3 s 74600 36960 75000 37016 6 qcpu_oeb[8]
port 330 nsew signal input
rlabel metal3 s 74600 37408 75000 37464 6 qcpu_oeb[9]
port 331 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 qcpu_sram_addr[0]
port 332 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 qcpu_sram_addr[1]
port 333 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 qcpu_sram_addr[2]
port 334 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 qcpu_sram_addr[3]
port 335 nsew signal input
rlabel metal2 s 61152 0 61208 400 6 qcpu_sram_addr[4]
port 336 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 qcpu_sram_addr[5]
port 337 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 qcpu_sram_gwe
port 338 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 qcpu_sram_in[0]
port 339 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 qcpu_sram_in[1]
port 340 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 qcpu_sram_in[2]
port 341 nsew signal input
rlabel metal2 s 63840 0 63896 400 6 qcpu_sram_in[3]
port 342 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 qcpu_sram_in[4]
port 343 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 qcpu_sram_in[5]
port 344 nsew signal input
rlabel metal2 s 65184 0 65240 400 6 qcpu_sram_in[6]
port 345 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 qcpu_sram_in[7]
port 346 nsew signal input
rlabel metal3 s 74600 48160 75000 48216 6 qcpu_sram_out[0]
port 347 nsew signal output
rlabel metal3 s 74600 48608 75000 48664 6 qcpu_sram_out[1]
port 348 nsew signal output
rlabel metal3 s 74600 49056 75000 49112 6 qcpu_sram_out[2]
port 349 nsew signal output
rlabel metal3 s 74600 49504 75000 49560 6 qcpu_sram_out[3]
port 350 nsew signal output
rlabel metal3 s 74600 49952 75000 50008 6 qcpu_sram_out[4]
port 351 nsew signal output
rlabel metal3 s 74600 50400 75000 50456 6 qcpu_sram_out[5]
port 352 nsew signal output
rlabel metal3 s 74600 50848 75000 50904 6 qcpu_sram_out[6]
port 353 nsew signal output
rlabel metal3 s 74600 51296 75000 51352 6 qcpu_sram_out[7]
port 354 nsew signal output
rlabel metal3 s 74600 51744 75000 51800 6 rst_ay8913
port 355 nsew signal output
rlabel metal3 s 0 62608 400 62664 6 rst_blinker
port 356 nsew signal output
rlabel metal2 s 62608 69600 62664 70000 6 rst_diceroll
port 357 nsew signal output
rlabel metal3 s 0 58128 400 58184 6 rst_hellorld
port 358 nsew signal output
rlabel metal3 s 0 40208 400 40264 6 rst_mc14500
port 359 nsew signal output
rlabel metal3 s 74600 52192 75000 52248 6 rst_pdp11
port 360 nsew signal output
rlabel metal3 s 0 39648 400 39704 6 rst_qcpu
port 361 nsew signal output
rlabel metal3 s 0 26768 400 26824 6 rst_sid
port 362 nsew signal output
rlabel metal2 s 19264 69600 19320 70000 6 rst_sn76489
port 363 nsew signal output
rlabel metal3 s 0 59248 400 59304 6 rst_tbb1143
port 364 nsew signal output
rlabel metal2 s 51184 69600 51240 70000 6 rst_tholin_riscv
port 365 nsew signal output
rlabel metal2 s 65968 69600 66024 70000 6 rst_ue1
port 366 nsew signal output
rlabel metal3 s 0 27328 400 27384 6 sid_do[0]
port 367 nsew signal input
rlabel metal3 s 0 32928 400 32984 6 sid_do[10]
port 368 nsew signal input
rlabel metal3 s 0 33488 400 33544 6 sid_do[11]
port 369 nsew signal input
rlabel metal3 s 0 34048 400 34104 6 sid_do[12]
port 370 nsew signal input
rlabel metal3 s 0 34608 400 34664 6 sid_do[13]
port 371 nsew signal input
rlabel metal3 s 0 35168 400 35224 6 sid_do[14]
port 372 nsew signal input
rlabel metal3 s 0 35728 400 35784 6 sid_do[15]
port 373 nsew signal input
rlabel metal3 s 0 36288 400 36344 6 sid_do[16]
port 374 nsew signal input
rlabel metal3 s 0 36848 400 36904 6 sid_do[17]
port 375 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 sid_do[18]
port 376 nsew signal input
rlabel metal3 s 0 37968 400 38024 6 sid_do[19]
port 377 nsew signal input
rlabel metal3 s 0 27888 400 27944 6 sid_do[1]
port 378 nsew signal input
rlabel metal3 s 0 38528 400 38584 6 sid_do[20]
port 379 nsew signal input
rlabel metal3 s 0 28448 400 28504 6 sid_do[2]
port 380 nsew signal input
rlabel metal3 s 0 29008 400 29064 6 sid_do[3]
port 381 nsew signal input
rlabel metal3 s 0 29568 400 29624 6 sid_do[4]
port 382 nsew signal input
rlabel metal3 s 0 30128 400 30184 6 sid_do[5]
port 383 nsew signal input
rlabel metal3 s 0 30688 400 30744 6 sid_do[6]
port 384 nsew signal input
rlabel metal3 s 0 31248 400 31304 6 sid_do[7]
port 385 nsew signal input
rlabel metal3 s 0 31808 400 31864 6 sid_do[8]
port 386 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 sid_do[9]
port 387 nsew signal input
rlabel metal3 s 0 39088 400 39144 6 sid_oeb
port 388 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 sn76489_do[0]
port 389 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 sn76489_do[10]
port 390 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 sn76489_do[11]
port 391 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 sn76489_do[12]
port 392 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 sn76489_do[13]
port 393 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 sn76489_do[14]
port 394 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 sn76489_do[15]
port 395 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 sn76489_do[16]
port 396 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 sn76489_do[17]
port 397 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 sn76489_do[18]
port 398 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 sn76489_do[19]
port 399 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 sn76489_do[1]
port 400 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 sn76489_do[20]
port 401 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 sn76489_do[21]
port 402 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 sn76489_do[22]
port 403 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 sn76489_do[23]
port 404 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 sn76489_do[24]
port 405 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 sn76489_do[25]
port 406 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 sn76489_do[26]
port 407 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 sn76489_do[27]
port 408 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 sn76489_do[2]
port 409 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 sn76489_do[3]
port 410 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 sn76489_do[4]
port 411 nsew signal input
rlabel metal2 s 34272 0 34328 400 6 sn76489_do[5]
port 412 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 sn76489_do[6]
port 413 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 sn76489_do[7]
port 414 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 sn76489_do[8]
port 415 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 sn76489_do[9]
port 416 nsew signal input
rlabel metal3 s 0 59808 400 59864 6 tbb1143_do[0]
port 417 nsew signal input
rlabel metal3 s 0 60368 400 60424 6 tbb1143_do[1]
port 418 nsew signal input
rlabel metal3 s 0 60928 400 60984 6 tbb1143_do[2]
port 419 nsew signal input
rlabel metal3 s 0 61488 400 61544 6 tbb1143_do[3]
port 420 nsew signal input
rlabel metal3 s 0 62048 400 62104 6 tbb1143_do[4]
port 421 nsew signal input
rlabel metal3 s 74600 52640 75000 52696 6 tholin_riscv_do[0]
port 422 nsew signal input
rlabel metal3 s 74600 57120 75000 57176 6 tholin_riscv_do[10]
port 423 nsew signal input
rlabel metal3 s 74600 57568 75000 57624 6 tholin_riscv_do[11]
port 424 nsew signal input
rlabel metal3 s 74600 58016 75000 58072 6 tholin_riscv_do[12]
port 425 nsew signal input
rlabel metal3 s 74600 58464 75000 58520 6 tholin_riscv_do[13]
port 426 nsew signal input
rlabel metal3 s 74600 58912 75000 58968 6 tholin_riscv_do[14]
port 427 nsew signal input
rlabel metal3 s 74600 59360 75000 59416 6 tholin_riscv_do[15]
port 428 nsew signal input
rlabel metal3 s 74600 59808 75000 59864 6 tholin_riscv_do[16]
port 429 nsew signal input
rlabel metal3 s 74600 60256 75000 60312 6 tholin_riscv_do[17]
port 430 nsew signal input
rlabel metal3 s 74600 60704 75000 60760 6 tholin_riscv_do[18]
port 431 nsew signal input
rlabel metal3 s 74600 61152 75000 61208 6 tholin_riscv_do[19]
port 432 nsew signal input
rlabel metal3 s 74600 53088 75000 53144 6 tholin_riscv_do[1]
port 433 nsew signal input
rlabel metal3 s 74600 61600 75000 61656 6 tholin_riscv_do[20]
port 434 nsew signal input
rlabel metal3 s 74600 62048 75000 62104 6 tholin_riscv_do[21]
port 435 nsew signal input
rlabel metal3 s 74600 62496 75000 62552 6 tholin_riscv_do[22]
port 436 nsew signal input
rlabel metal3 s 74600 62944 75000 63000 6 tholin_riscv_do[23]
port 437 nsew signal input
rlabel metal3 s 74600 63392 75000 63448 6 tholin_riscv_do[24]
port 438 nsew signal input
rlabel metal3 s 74600 63840 75000 63896 6 tholin_riscv_do[25]
port 439 nsew signal input
rlabel metal3 s 74600 64288 75000 64344 6 tholin_riscv_do[26]
port 440 nsew signal input
rlabel metal3 s 74600 64736 75000 64792 6 tholin_riscv_do[27]
port 441 nsew signal input
rlabel metal3 s 74600 65184 75000 65240 6 tholin_riscv_do[28]
port 442 nsew signal input
rlabel metal3 s 74600 65632 75000 65688 6 tholin_riscv_do[29]
port 443 nsew signal input
rlabel metal3 s 74600 53536 75000 53592 6 tholin_riscv_do[2]
port 444 nsew signal input
rlabel metal3 s 74600 66080 75000 66136 6 tholin_riscv_do[30]
port 445 nsew signal input
rlabel metal3 s 74600 66528 75000 66584 6 tholin_riscv_do[31]
port 446 nsew signal input
rlabel metal3 s 74600 66976 75000 67032 6 tholin_riscv_do[32]
port 447 nsew signal input
rlabel metal3 s 74600 53984 75000 54040 6 tholin_riscv_do[3]
port 448 nsew signal input
rlabel metal3 s 74600 54432 75000 54488 6 tholin_riscv_do[4]
port 449 nsew signal input
rlabel metal3 s 74600 54880 75000 54936 6 tholin_riscv_do[5]
port 450 nsew signal input
rlabel metal3 s 74600 55328 75000 55384 6 tholin_riscv_do[6]
port 451 nsew signal input
rlabel metal3 s 74600 55776 75000 55832 6 tholin_riscv_do[7]
port 452 nsew signal input
rlabel metal3 s 74600 56224 75000 56280 6 tholin_riscv_do[8]
port 453 nsew signal input
rlabel metal3 s 74600 56672 75000 56728 6 tholin_riscv_do[9]
port 454 nsew signal input
rlabel metal2 s 51520 69600 51576 70000 6 tholin_riscv_oeb[0]
port 455 nsew signal input
rlabel metal2 s 54880 69600 54936 70000 6 tholin_riscv_oeb[10]
port 456 nsew signal input
rlabel metal2 s 55216 69600 55272 70000 6 tholin_riscv_oeb[11]
port 457 nsew signal input
rlabel metal2 s 55552 69600 55608 70000 6 tholin_riscv_oeb[12]
port 458 nsew signal input
rlabel metal2 s 55888 69600 55944 70000 6 tholin_riscv_oeb[13]
port 459 nsew signal input
rlabel metal2 s 56224 69600 56280 70000 6 tholin_riscv_oeb[14]
port 460 nsew signal input
rlabel metal2 s 56560 69600 56616 70000 6 tholin_riscv_oeb[15]
port 461 nsew signal input
rlabel metal2 s 56896 69600 56952 70000 6 tholin_riscv_oeb[16]
port 462 nsew signal input
rlabel metal2 s 57232 69600 57288 70000 6 tholin_riscv_oeb[17]
port 463 nsew signal input
rlabel metal2 s 57568 69600 57624 70000 6 tholin_riscv_oeb[18]
port 464 nsew signal input
rlabel metal2 s 57904 69600 57960 70000 6 tholin_riscv_oeb[19]
port 465 nsew signal input
rlabel metal2 s 51856 69600 51912 70000 6 tholin_riscv_oeb[1]
port 466 nsew signal input
rlabel metal2 s 58240 69600 58296 70000 6 tholin_riscv_oeb[20]
port 467 nsew signal input
rlabel metal2 s 58576 69600 58632 70000 6 tholin_riscv_oeb[21]
port 468 nsew signal input
rlabel metal2 s 58912 69600 58968 70000 6 tholin_riscv_oeb[22]
port 469 nsew signal input
rlabel metal2 s 59248 69600 59304 70000 6 tholin_riscv_oeb[23]
port 470 nsew signal input
rlabel metal2 s 59584 69600 59640 70000 6 tholin_riscv_oeb[24]
port 471 nsew signal input
rlabel metal2 s 59920 69600 59976 70000 6 tholin_riscv_oeb[25]
port 472 nsew signal input
rlabel metal2 s 60256 69600 60312 70000 6 tholin_riscv_oeb[26]
port 473 nsew signal input
rlabel metal2 s 60592 69600 60648 70000 6 tholin_riscv_oeb[27]
port 474 nsew signal input
rlabel metal2 s 60928 69600 60984 70000 6 tholin_riscv_oeb[28]
port 475 nsew signal input
rlabel metal2 s 61264 69600 61320 70000 6 tholin_riscv_oeb[29]
port 476 nsew signal input
rlabel metal2 s 52192 69600 52248 70000 6 tholin_riscv_oeb[2]
port 477 nsew signal input
rlabel metal2 s 61600 69600 61656 70000 6 tholin_riscv_oeb[30]
port 478 nsew signal input
rlabel metal2 s 61936 69600 61992 70000 6 tholin_riscv_oeb[31]
port 479 nsew signal input
rlabel metal2 s 62272 69600 62328 70000 6 tholin_riscv_oeb[32]
port 480 nsew signal input
rlabel metal2 s 52528 69600 52584 70000 6 tholin_riscv_oeb[3]
port 481 nsew signal input
rlabel metal2 s 52864 69600 52920 70000 6 tholin_riscv_oeb[4]
port 482 nsew signal input
rlabel metal2 s 53200 69600 53256 70000 6 tholin_riscv_oeb[5]
port 483 nsew signal input
rlabel metal2 s 53536 69600 53592 70000 6 tholin_riscv_oeb[6]
port 484 nsew signal input
rlabel metal2 s 53872 69600 53928 70000 6 tholin_riscv_oeb[7]
port 485 nsew signal input
rlabel metal2 s 54208 69600 54264 70000 6 tholin_riscv_oeb[8]
port 486 nsew signal input
rlabel metal2 s 54544 69600 54600 70000 6 tholin_riscv_oeb[9]
port 487 nsew signal input
rlabel metal2 s 66640 69600 66696 70000 6 ue1_do[0]
port 488 nsew signal input
rlabel metal2 s 66976 69600 67032 70000 6 ue1_do[1]
port 489 nsew signal input
rlabel metal2 s 67312 69600 67368 70000 6 ue1_do[2]
port 490 nsew signal input
rlabel metal2 s 67648 69600 67704 70000 6 ue1_do[3]
port 491 nsew signal input
rlabel metal2 s 67984 69600 68040 70000 6 ue1_do[4]
port 492 nsew signal input
rlabel metal2 s 68320 69600 68376 70000 6 ue1_do[5]
port 493 nsew signal input
rlabel metal2 s 68656 69600 68712 70000 6 ue1_do[6]
port 494 nsew signal input
rlabel metal2 s 68992 69600 69048 70000 6 ue1_do[7]
port 495 nsew signal input
rlabel metal2 s 69328 69600 69384 70000 6 ue1_do[8]
port 496 nsew signal input
rlabel metal2 s 69664 69600 69720 70000 6 ue1_do[9]
port 497 nsew signal input
rlabel metal2 s 66304 69600 66360 70000 6 ue1_oeb
port 498 nsew signal input
rlabel metal4 s 2224 1538 2384 68238 6 vdd
port 499 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 68238 6 vdd
port 499 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 68238 6 vdd
port 499 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 68238 6 vdd
port 499 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 68238 6 vdd
port 499 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 68238 6 vss
port 500 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 68238 6 vss
port 500 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 68238 6 vss
port 500 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 68238 6 vss
port 500 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 68238 6 vss
port 500 nsew ground bidirectional
rlabel metal2 s 2464 0 2520 400 6 wb_clk_i
port 501 nsew signal input
rlabel metal2 s 2912 0 2968 400 6 wb_rst_i
port 502 nsew signal input
rlabel metal3 s 74600 18592 75000 18648 6 wbs_ack_o
port 503 nsew signal output
rlabel metal2 s 3360 0 3416 400 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal2 s 9184 0 9240 400 6 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal2 s 17248 0 17304 400 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal3 s 74600 17696 75000 17752 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal2 s 28896 0 28952 400 6 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal3 s 74600 2912 75000 2968 6 wbs_dat_o[0]
port 569 nsew signal output
rlabel metal3 s 74600 7392 75000 7448 6 wbs_dat_o[10]
port 570 nsew signal output
rlabel metal3 s 74600 7840 75000 7896 6 wbs_dat_o[11]
port 571 nsew signal output
rlabel metal3 s 74600 8288 75000 8344 6 wbs_dat_o[12]
port 572 nsew signal output
rlabel metal3 s 74600 8736 75000 8792 6 wbs_dat_o[13]
port 573 nsew signal output
rlabel metal3 s 74600 9184 75000 9240 6 wbs_dat_o[14]
port 574 nsew signal output
rlabel metal3 s 74600 9632 75000 9688 6 wbs_dat_o[15]
port 575 nsew signal output
rlabel metal3 s 74600 10080 75000 10136 6 wbs_dat_o[16]
port 576 nsew signal output
rlabel metal3 s 74600 10528 75000 10584 6 wbs_dat_o[17]
port 577 nsew signal output
rlabel metal3 s 74600 10976 75000 11032 6 wbs_dat_o[18]
port 578 nsew signal output
rlabel metal3 s 74600 11424 75000 11480 6 wbs_dat_o[19]
port 579 nsew signal output
rlabel metal3 s 74600 3360 75000 3416 6 wbs_dat_o[1]
port 580 nsew signal output
rlabel metal3 s 74600 11872 75000 11928 6 wbs_dat_o[20]
port 581 nsew signal output
rlabel metal3 s 74600 12320 75000 12376 6 wbs_dat_o[21]
port 582 nsew signal output
rlabel metal3 s 74600 12768 75000 12824 6 wbs_dat_o[22]
port 583 nsew signal output
rlabel metal3 s 74600 13216 75000 13272 6 wbs_dat_o[23]
port 584 nsew signal output
rlabel metal3 s 74600 13664 75000 13720 6 wbs_dat_o[24]
port 585 nsew signal output
rlabel metal3 s 74600 14112 75000 14168 6 wbs_dat_o[25]
port 586 nsew signal output
rlabel metal3 s 74600 14560 75000 14616 6 wbs_dat_o[26]
port 587 nsew signal output
rlabel metal3 s 74600 15008 75000 15064 6 wbs_dat_o[27]
port 588 nsew signal output
rlabel metal3 s 74600 15456 75000 15512 6 wbs_dat_o[28]
port 589 nsew signal output
rlabel metal3 s 74600 15904 75000 15960 6 wbs_dat_o[29]
port 590 nsew signal output
rlabel metal3 s 74600 3808 75000 3864 6 wbs_dat_o[2]
port 591 nsew signal output
rlabel metal3 s 74600 16352 75000 16408 6 wbs_dat_o[30]
port 592 nsew signal output
rlabel metal3 s 74600 16800 75000 16856 6 wbs_dat_o[31]
port 593 nsew signal output
rlabel metal3 s 74600 4256 75000 4312 6 wbs_dat_o[3]
port 594 nsew signal output
rlabel metal3 s 74600 4704 75000 4760 6 wbs_dat_o[4]
port 595 nsew signal output
rlabel metal3 s 74600 5152 75000 5208 6 wbs_dat_o[5]
port 596 nsew signal output
rlabel metal3 s 74600 5600 75000 5656 6 wbs_dat_o[6]
port 597 nsew signal output
rlabel metal3 s 74600 6048 75000 6104 6 wbs_dat_o[7]
port 598 nsew signal output
rlabel metal3 s 74600 6496 75000 6552 6 wbs_dat_o[8]
port 599 nsew signal output
rlabel metal3 s 74600 6944 75000 7000 6 wbs_dat_o[9]
port 600 nsew signal output
rlabel metal3 s 74600 18144 75000 18200 6 wbs_stb_i
port 601 nsew signal input
rlabel metal3 s 74600 17248 75000 17304 6 wbs_we_i
port 602 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 75000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9738112
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/Multiplexer/runs/23_12_13_16_01/results/signoff/multiplexer.magic.gds
string GDS_START 407388
<< end >>

