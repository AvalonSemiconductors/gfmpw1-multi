magic
tech gf180mcuD
magscale 1 5
timestamp 1700060047
<< obsm1 >>
rect 672 1415 64288 64105
<< metal2 >>
rect 4144 64600 4200 65000
rect 4592 64600 4648 65000
rect 5040 64600 5096 65000
rect 5488 64600 5544 65000
rect 5936 64600 5992 65000
rect 6384 64600 6440 65000
rect 6832 64600 6888 65000
rect 7280 64600 7336 65000
rect 7728 64600 7784 65000
rect 8176 64600 8232 65000
rect 8624 64600 8680 65000
rect 9072 64600 9128 65000
rect 9520 64600 9576 65000
rect 9968 64600 10024 65000
rect 10416 64600 10472 65000
rect 10864 64600 10920 65000
rect 11312 64600 11368 65000
rect 11760 64600 11816 65000
rect 12208 64600 12264 65000
rect 12656 64600 12712 65000
rect 13104 64600 13160 65000
rect 13552 64600 13608 65000
rect 14000 64600 14056 65000
rect 14448 64600 14504 65000
rect 14896 64600 14952 65000
rect 15344 64600 15400 65000
rect 15792 64600 15848 65000
rect 16240 64600 16296 65000
rect 16688 64600 16744 65000
rect 17136 64600 17192 65000
rect 17584 64600 17640 65000
rect 18032 64600 18088 65000
rect 18480 64600 18536 65000
rect 18928 64600 18984 65000
rect 19376 64600 19432 65000
rect 19824 64600 19880 65000
rect 20272 64600 20328 65000
rect 20720 64600 20776 65000
rect 21168 64600 21224 65000
rect 21616 64600 21672 65000
rect 22064 64600 22120 65000
rect 22512 64600 22568 65000
rect 22960 64600 23016 65000
rect 23408 64600 23464 65000
rect 23856 64600 23912 65000
rect 24304 64600 24360 65000
rect 24752 64600 24808 65000
rect 25200 64600 25256 65000
rect 25648 64600 25704 65000
rect 26096 64600 26152 65000
rect 26544 64600 26600 65000
rect 26992 64600 27048 65000
rect 27440 64600 27496 65000
rect 27888 64600 27944 65000
rect 28336 64600 28392 65000
rect 28784 64600 28840 65000
rect 29232 64600 29288 65000
rect 29680 64600 29736 65000
rect 30128 64600 30184 65000
rect 30576 64600 30632 65000
rect 31024 64600 31080 65000
rect 31472 64600 31528 65000
rect 31920 64600 31976 65000
rect 32368 64600 32424 65000
rect 32816 64600 32872 65000
rect 33264 64600 33320 65000
rect 33712 64600 33768 65000
rect 34160 64600 34216 65000
rect 34608 64600 34664 65000
rect 35056 64600 35112 65000
rect 35504 64600 35560 65000
rect 35952 64600 36008 65000
rect 36400 64600 36456 65000
rect 36848 64600 36904 65000
rect 37296 64600 37352 65000
rect 37744 64600 37800 65000
rect 38192 64600 38248 65000
rect 38640 64600 38696 65000
rect 39088 64600 39144 65000
rect 39536 64600 39592 65000
rect 39984 64600 40040 65000
rect 40432 64600 40488 65000
rect 40880 64600 40936 65000
rect 41328 64600 41384 65000
rect 41776 64600 41832 65000
rect 42224 64600 42280 65000
rect 42672 64600 42728 65000
rect 43120 64600 43176 65000
rect 43568 64600 43624 65000
rect 44016 64600 44072 65000
rect 44464 64600 44520 65000
rect 44912 64600 44968 65000
rect 45360 64600 45416 65000
rect 45808 64600 45864 65000
rect 46256 64600 46312 65000
rect 46704 64600 46760 65000
rect 47152 64600 47208 65000
rect 47600 64600 47656 65000
rect 48048 64600 48104 65000
rect 48496 64600 48552 65000
rect 48944 64600 49000 65000
rect 49392 64600 49448 65000
rect 49840 64600 49896 65000
rect 50288 64600 50344 65000
rect 50736 64600 50792 65000
rect 51184 64600 51240 65000
rect 51632 64600 51688 65000
rect 52080 64600 52136 65000
rect 52528 64600 52584 65000
rect 52976 64600 53032 65000
rect 53424 64600 53480 65000
rect 53872 64600 53928 65000
rect 54320 64600 54376 65000
rect 54768 64600 54824 65000
rect 55216 64600 55272 65000
rect 55664 64600 55720 65000
rect 56112 64600 56168 65000
rect 56560 64600 56616 65000
rect 57008 64600 57064 65000
rect 57456 64600 57512 65000
rect 57904 64600 57960 65000
rect 58352 64600 58408 65000
rect 58800 64600 58856 65000
rect 59248 64600 59304 65000
rect 59696 64600 59752 65000
rect 60144 64600 60200 65000
rect 60592 64600 60648 65000
rect 2576 0 2632 400
rect 3024 0 3080 400
rect 3472 0 3528 400
rect 3920 0 3976 400
rect 4368 0 4424 400
rect 4816 0 4872 400
rect 5264 0 5320 400
rect 5712 0 5768 400
rect 6160 0 6216 400
rect 6608 0 6664 400
rect 7056 0 7112 400
rect 7504 0 7560 400
rect 7952 0 8008 400
rect 8400 0 8456 400
rect 8848 0 8904 400
rect 9296 0 9352 400
rect 9744 0 9800 400
rect 10192 0 10248 400
rect 10640 0 10696 400
rect 11088 0 11144 400
rect 11536 0 11592 400
rect 11984 0 12040 400
rect 12432 0 12488 400
rect 12880 0 12936 400
rect 13328 0 13384 400
rect 13776 0 13832 400
rect 14224 0 14280 400
rect 14672 0 14728 400
rect 15120 0 15176 400
rect 15568 0 15624 400
rect 16016 0 16072 400
rect 16464 0 16520 400
rect 16912 0 16968 400
rect 17360 0 17416 400
rect 17808 0 17864 400
rect 18256 0 18312 400
rect 18704 0 18760 400
rect 19152 0 19208 400
rect 19600 0 19656 400
rect 20048 0 20104 400
rect 20496 0 20552 400
rect 20944 0 21000 400
rect 21392 0 21448 400
rect 21840 0 21896 400
rect 22288 0 22344 400
rect 22736 0 22792 400
rect 23184 0 23240 400
rect 23632 0 23688 400
rect 24080 0 24136 400
rect 24528 0 24584 400
rect 24976 0 25032 400
rect 25424 0 25480 400
rect 25872 0 25928 400
rect 26320 0 26376 400
rect 26768 0 26824 400
rect 27216 0 27272 400
rect 27664 0 27720 400
rect 28112 0 28168 400
rect 28560 0 28616 400
rect 29008 0 29064 400
rect 29456 0 29512 400
rect 29904 0 29960 400
rect 30352 0 30408 400
rect 30800 0 30856 400
rect 31248 0 31304 400
rect 31696 0 31752 400
rect 32144 0 32200 400
rect 32592 0 32648 400
rect 33040 0 33096 400
rect 33488 0 33544 400
rect 33936 0 33992 400
rect 34384 0 34440 400
rect 34832 0 34888 400
rect 35280 0 35336 400
rect 35728 0 35784 400
rect 36176 0 36232 400
rect 36624 0 36680 400
rect 37072 0 37128 400
rect 37520 0 37576 400
rect 37968 0 38024 400
rect 38416 0 38472 400
rect 38864 0 38920 400
rect 39312 0 39368 400
rect 39760 0 39816 400
rect 40208 0 40264 400
rect 40656 0 40712 400
rect 41104 0 41160 400
rect 41552 0 41608 400
rect 42000 0 42056 400
rect 42448 0 42504 400
rect 42896 0 42952 400
rect 43344 0 43400 400
rect 43792 0 43848 400
rect 44240 0 44296 400
rect 44688 0 44744 400
rect 45136 0 45192 400
rect 45584 0 45640 400
rect 46032 0 46088 400
rect 46480 0 46536 400
rect 46928 0 46984 400
rect 47376 0 47432 400
rect 47824 0 47880 400
rect 48272 0 48328 400
rect 48720 0 48776 400
rect 49168 0 49224 400
rect 49616 0 49672 400
rect 50064 0 50120 400
rect 50512 0 50568 400
rect 50960 0 51016 400
rect 51408 0 51464 400
rect 51856 0 51912 400
rect 52304 0 52360 400
rect 52752 0 52808 400
rect 53200 0 53256 400
rect 53648 0 53704 400
rect 54096 0 54152 400
rect 54544 0 54600 400
rect 54992 0 55048 400
rect 55440 0 55496 400
rect 55888 0 55944 400
rect 56336 0 56392 400
rect 56784 0 56840 400
rect 57232 0 57288 400
rect 57680 0 57736 400
rect 58128 0 58184 400
rect 58576 0 58632 400
rect 59024 0 59080 400
rect 59472 0 59528 400
rect 59920 0 59976 400
rect 60368 0 60424 400
rect 60816 0 60872 400
rect 61264 0 61320 400
rect 61712 0 61768 400
rect 62160 0 62216 400
<< obsm2 >>
rect 742 64570 4114 64666
rect 4230 64570 4562 64666
rect 4678 64570 5010 64666
rect 5126 64570 5458 64666
rect 5574 64570 5906 64666
rect 6022 64570 6354 64666
rect 6470 64570 6802 64666
rect 6918 64570 7250 64666
rect 7366 64570 7698 64666
rect 7814 64570 8146 64666
rect 8262 64570 8594 64666
rect 8710 64570 9042 64666
rect 9158 64570 9490 64666
rect 9606 64570 9938 64666
rect 10054 64570 10386 64666
rect 10502 64570 10834 64666
rect 10950 64570 11282 64666
rect 11398 64570 11730 64666
rect 11846 64570 12178 64666
rect 12294 64570 12626 64666
rect 12742 64570 13074 64666
rect 13190 64570 13522 64666
rect 13638 64570 13970 64666
rect 14086 64570 14418 64666
rect 14534 64570 14866 64666
rect 14982 64570 15314 64666
rect 15430 64570 15762 64666
rect 15878 64570 16210 64666
rect 16326 64570 16658 64666
rect 16774 64570 17106 64666
rect 17222 64570 17554 64666
rect 17670 64570 18002 64666
rect 18118 64570 18450 64666
rect 18566 64570 18898 64666
rect 19014 64570 19346 64666
rect 19462 64570 19794 64666
rect 19910 64570 20242 64666
rect 20358 64570 20690 64666
rect 20806 64570 21138 64666
rect 21254 64570 21586 64666
rect 21702 64570 22034 64666
rect 22150 64570 22482 64666
rect 22598 64570 22930 64666
rect 23046 64570 23378 64666
rect 23494 64570 23826 64666
rect 23942 64570 24274 64666
rect 24390 64570 24722 64666
rect 24838 64570 25170 64666
rect 25286 64570 25618 64666
rect 25734 64570 26066 64666
rect 26182 64570 26514 64666
rect 26630 64570 26962 64666
rect 27078 64570 27410 64666
rect 27526 64570 27858 64666
rect 27974 64570 28306 64666
rect 28422 64570 28754 64666
rect 28870 64570 29202 64666
rect 29318 64570 29650 64666
rect 29766 64570 30098 64666
rect 30214 64570 30546 64666
rect 30662 64570 30994 64666
rect 31110 64570 31442 64666
rect 31558 64570 31890 64666
rect 32006 64570 32338 64666
rect 32454 64570 32786 64666
rect 32902 64570 33234 64666
rect 33350 64570 33682 64666
rect 33798 64570 34130 64666
rect 34246 64570 34578 64666
rect 34694 64570 35026 64666
rect 35142 64570 35474 64666
rect 35590 64570 35922 64666
rect 36038 64570 36370 64666
rect 36486 64570 36818 64666
rect 36934 64570 37266 64666
rect 37382 64570 37714 64666
rect 37830 64570 38162 64666
rect 38278 64570 38610 64666
rect 38726 64570 39058 64666
rect 39174 64570 39506 64666
rect 39622 64570 39954 64666
rect 40070 64570 40402 64666
rect 40518 64570 40850 64666
rect 40966 64570 41298 64666
rect 41414 64570 41746 64666
rect 41862 64570 42194 64666
rect 42310 64570 42642 64666
rect 42758 64570 43090 64666
rect 43206 64570 43538 64666
rect 43654 64570 43986 64666
rect 44102 64570 44434 64666
rect 44550 64570 44882 64666
rect 44998 64570 45330 64666
rect 45446 64570 45778 64666
rect 45894 64570 46226 64666
rect 46342 64570 46674 64666
rect 46790 64570 47122 64666
rect 47238 64570 47570 64666
rect 47686 64570 48018 64666
rect 48134 64570 48466 64666
rect 48582 64570 48914 64666
rect 49030 64570 49362 64666
rect 49478 64570 49810 64666
rect 49926 64570 50258 64666
rect 50374 64570 50706 64666
rect 50822 64570 51154 64666
rect 51270 64570 51602 64666
rect 51718 64570 52050 64666
rect 52166 64570 52498 64666
rect 52614 64570 52946 64666
rect 53062 64570 53394 64666
rect 53510 64570 53842 64666
rect 53958 64570 54290 64666
rect 54406 64570 54738 64666
rect 54854 64570 55186 64666
rect 55302 64570 55634 64666
rect 55750 64570 56082 64666
rect 56198 64570 56530 64666
rect 56646 64570 56978 64666
rect 57094 64570 57426 64666
rect 57542 64570 57874 64666
rect 57990 64570 58322 64666
rect 58438 64570 58770 64666
rect 58886 64570 59218 64666
rect 59334 64570 59666 64666
rect 59782 64570 60114 64666
rect 60230 64570 60562 64666
rect 60678 64570 64610 64666
rect 742 430 64610 64570
rect 742 350 2546 430
rect 2662 350 2994 430
rect 3110 350 3442 430
rect 3558 350 3890 430
rect 4006 350 4338 430
rect 4454 350 4786 430
rect 4902 350 5234 430
rect 5350 350 5682 430
rect 5798 350 6130 430
rect 6246 350 6578 430
rect 6694 350 7026 430
rect 7142 350 7474 430
rect 7590 350 7922 430
rect 8038 350 8370 430
rect 8486 350 8818 430
rect 8934 350 9266 430
rect 9382 350 9714 430
rect 9830 350 10162 430
rect 10278 350 10610 430
rect 10726 350 11058 430
rect 11174 350 11506 430
rect 11622 350 11954 430
rect 12070 350 12402 430
rect 12518 350 12850 430
rect 12966 350 13298 430
rect 13414 350 13746 430
rect 13862 350 14194 430
rect 14310 350 14642 430
rect 14758 350 15090 430
rect 15206 350 15538 430
rect 15654 350 15986 430
rect 16102 350 16434 430
rect 16550 350 16882 430
rect 16998 350 17330 430
rect 17446 350 17778 430
rect 17894 350 18226 430
rect 18342 350 18674 430
rect 18790 350 19122 430
rect 19238 350 19570 430
rect 19686 350 20018 430
rect 20134 350 20466 430
rect 20582 350 20914 430
rect 21030 350 21362 430
rect 21478 350 21810 430
rect 21926 350 22258 430
rect 22374 350 22706 430
rect 22822 350 23154 430
rect 23270 350 23602 430
rect 23718 350 24050 430
rect 24166 350 24498 430
rect 24614 350 24946 430
rect 25062 350 25394 430
rect 25510 350 25842 430
rect 25958 350 26290 430
rect 26406 350 26738 430
rect 26854 350 27186 430
rect 27302 350 27634 430
rect 27750 350 28082 430
rect 28198 350 28530 430
rect 28646 350 28978 430
rect 29094 350 29426 430
rect 29542 350 29874 430
rect 29990 350 30322 430
rect 30438 350 30770 430
rect 30886 350 31218 430
rect 31334 350 31666 430
rect 31782 350 32114 430
rect 32230 350 32562 430
rect 32678 350 33010 430
rect 33126 350 33458 430
rect 33574 350 33906 430
rect 34022 350 34354 430
rect 34470 350 34802 430
rect 34918 350 35250 430
rect 35366 350 35698 430
rect 35814 350 36146 430
rect 36262 350 36594 430
rect 36710 350 37042 430
rect 37158 350 37490 430
rect 37606 350 37938 430
rect 38054 350 38386 430
rect 38502 350 38834 430
rect 38950 350 39282 430
rect 39398 350 39730 430
rect 39846 350 40178 430
rect 40294 350 40626 430
rect 40742 350 41074 430
rect 41190 350 41522 430
rect 41638 350 41970 430
rect 42086 350 42418 430
rect 42534 350 42866 430
rect 42982 350 43314 430
rect 43430 350 43762 430
rect 43878 350 44210 430
rect 44326 350 44658 430
rect 44774 350 45106 430
rect 45222 350 45554 430
rect 45670 350 46002 430
rect 46118 350 46450 430
rect 46566 350 46898 430
rect 47014 350 47346 430
rect 47462 350 47794 430
rect 47910 350 48242 430
rect 48358 350 48690 430
rect 48806 350 49138 430
rect 49254 350 49586 430
rect 49702 350 50034 430
rect 50150 350 50482 430
rect 50598 350 50930 430
rect 51046 350 51378 430
rect 51494 350 51826 430
rect 51942 350 52274 430
rect 52390 350 52722 430
rect 52838 350 53170 430
rect 53286 350 53618 430
rect 53734 350 54066 430
rect 54182 350 54514 430
rect 54630 350 54962 430
rect 55078 350 55410 430
rect 55526 350 55858 430
rect 55974 350 56306 430
rect 56422 350 56754 430
rect 56870 350 57202 430
rect 57318 350 57650 430
rect 57766 350 58098 430
rect 58214 350 58546 430
rect 58662 350 58994 430
rect 59110 350 59442 430
rect 59558 350 59890 430
rect 60006 350 60338 430
rect 60454 350 60786 430
rect 60902 350 61234 430
rect 61350 350 61682 430
rect 61798 350 62130 430
rect 62246 350 64610 430
<< metal3 >>
rect 0 60704 400 60760
rect 0 60144 400 60200
rect 0 59584 400 59640
rect 0 59024 400 59080
rect 64600 58576 65000 58632
rect 0 58464 400 58520
rect 64600 58128 65000 58184
rect 0 57904 400 57960
rect 64600 57680 65000 57736
rect 0 57344 400 57400
rect 64600 57232 65000 57288
rect 0 56784 400 56840
rect 64600 56784 65000 56840
rect 64600 56336 65000 56392
rect 0 56224 400 56280
rect 64600 55888 65000 55944
rect 0 55664 400 55720
rect 64600 55440 65000 55496
rect 0 55104 400 55160
rect 64600 54992 65000 55048
rect 0 54544 400 54600
rect 64600 54544 65000 54600
rect 64600 54096 65000 54152
rect 0 53984 400 54040
rect 64600 53648 65000 53704
rect 0 53424 400 53480
rect 64600 53200 65000 53256
rect 0 52864 400 52920
rect 64600 52752 65000 52808
rect 0 52304 400 52360
rect 64600 52304 65000 52360
rect 64600 51856 65000 51912
rect 0 51744 400 51800
rect 64600 51408 65000 51464
rect 0 51184 400 51240
rect 64600 50960 65000 51016
rect 0 50624 400 50680
rect 64600 50512 65000 50568
rect 0 50064 400 50120
rect 64600 50064 65000 50120
rect 64600 49616 65000 49672
rect 0 49504 400 49560
rect 64600 49168 65000 49224
rect 0 48944 400 49000
rect 64600 48720 65000 48776
rect 0 48384 400 48440
rect 64600 48272 65000 48328
rect 0 47824 400 47880
rect 64600 47824 65000 47880
rect 64600 47376 65000 47432
rect 0 47264 400 47320
rect 64600 46928 65000 46984
rect 0 46704 400 46760
rect 64600 46480 65000 46536
rect 0 46144 400 46200
rect 64600 46032 65000 46088
rect 0 45584 400 45640
rect 64600 45584 65000 45640
rect 64600 45136 65000 45192
rect 0 45024 400 45080
rect 64600 44688 65000 44744
rect 0 44464 400 44520
rect 64600 44240 65000 44296
rect 0 43904 400 43960
rect 64600 43792 65000 43848
rect 0 43344 400 43400
rect 64600 43344 65000 43400
rect 64600 42896 65000 42952
rect 0 42784 400 42840
rect 64600 42448 65000 42504
rect 0 42224 400 42280
rect 64600 42000 65000 42056
rect 0 41664 400 41720
rect 64600 41552 65000 41608
rect 0 41104 400 41160
rect 64600 41104 65000 41160
rect 64600 40656 65000 40712
rect 0 40544 400 40600
rect 64600 40208 65000 40264
rect 0 39984 400 40040
rect 64600 39760 65000 39816
rect 0 39424 400 39480
rect 64600 39312 65000 39368
rect 0 38864 400 38920
rect 64600 38864 65000 38920
rect 64600 38416 65000 38472
rect 0 38304 400 38360
rect 64600 37968 65000 38024
rect 0 37744 400 37800
rect 64600 37520 65000 37576
rect 0 37184 400 37240
rect 64600 37072 65000 37128
rect 0 36624 400 36680
rect 64600 36624 65000 36680
rect 64600 36176 65000 36232
rect 0 36064 400 36120
rect 64600 35728 65000 35784
rect 0 35504 400 35560
rect 64600 35280 65000 35336
rect 0 34944 400 35000
rect 64600 34832 65000 34888
rect 0 34384 400 34440
rect 64600 34384 65000 34440
rect 64600 33936 65000 33992
rect 0 33824 400 33880
rect 64600 33488 65000 33544
rect 0 33264 400 33320
rect 64600 33040 65000 33096
rect 0 32704 400 32760
rect 64600 32592 65000 32648
rect 0 32144 400 32200
rect 64600 32144 65000 32200
rect 64600 31696 65000 31752
rect 0 31584 400 31640
rect 64600 31248 65000 31304
rect 0 31024 400 31080
rect 64600 30800 65000 30856
rect 0 30464 400 30520
rect 64600 30352 65000 30408
rect 0 29904 400 29960
rect 64600 29904 65000 29960
rect 64600 29456 65000 29512
rect 0 29344 400 29400
rect 64600 29008 65000 29064
rect 0 28784 400 28840
rect 64600 28560 65000 28616
rect 0 28224 400 28280
rect 64600 28112 65000 28168
rect 0 27664 400 27720
rect 64600 27664 65000 27720
rect 64600 27216 65000 27272
rect 0 27104 400 27160
rect 64600 26768 65000 26824
rect 0 26544 400 26600
rect 64600 26320 65000 26376
rect 0 25984 400 26040
rect 64600 25872 65000 25928
rect 0 25424 400 25480
rect 64600 25424 65000 25480
rect 64600 24976 65000 25032
rect 0 24864 400 24920
rect 64600 24528 65000 24584
rect 0 24304 400 24360
rect 64600 24080 65000 24136
rect 0 23744 400 23800
rect 64600 23632 65000 23688
rect 0 23184 400 23240
rect 64600 23184 65000 23240
rect 64600 22736 65000 22792
rect 0 22624 400 22680
rect 64600 22288 65000 22344
rect 0 22064 400 22120
rect 64600 21840 65000 21896
rect 0 21504 400 21560
rect 64600 21392 65000 21448
rect 0 20944 400 21000
rect 64600 20944 65000 21000
rect 64600 20496 65000 20552
rect 0 20384 400 20440
rect 64600 20048 65000 20104
rect 0 19824 400 19880
rect 64600 19600 65000 19656
rect 0 19264 400 19320
rect 64600 19152 65000 19208
rect 0 18704 400 18760
rect 64600 18704 65000 18760
rect 64600 18256 65000 18312
rect 0 18144 400 18200
rect 64600 17808 65000 17864
rect 0 17584 400 17640
rect 64600 17360 65000 17416
rect 0 17024 400 17080
rect 64600 16912 65000 16968
rect 0 16464 400 16520
rect 64600 16464 65000 16520
rect 64600 16016 65000 16072
rect 0 15904 400 15960
rect 64600 15568 65000 15624
rect 0 15344 400 15400
rect 64600 15120 65000 15176
rect 0 14784 400 14840
rect 64600 14672 65000 14728
rect 0 14224 400 14280
rect 64600 14224 65000 14280
rect 64600 13776 65000 13832
rect 0 13664 400 13720
rect 64600 13328 65000 13384
rect 0 13104 400 13160
rect 64600 12880 65000 12936
rect 0 12544 400 12600
rect 64600 12432 65000 12488
rect 0 11984 400 12040
rect 64600 11984 65000 12040
rect 64600 11536 65000 11592
rect 0 11424 400 11480
rect 64600 11088 65000 11144
rect 0 10864 400 10920
rect 64600 10640 65000 10696
rect 0 10304 400 10360
rect 64600 10192 65000 10248
rect 0 9744 400 9800
rect 64600 9744 65000 9800
rect 64600 9296 65000 9352
rect 0 9184 400 9240
rect 64600 8848 65000 8904
rect 0 8624 400 8680
rect 64600 8400 65000 8456
rect 0 8064 400 8120
rect 64600 7952 65000 8008
rect 0 7504 400 7560
rect 64600 7504 65000 7560
rect 64600 7056 65000 7112
rect 0 6944 400 7000
rect 64600 6608 65000 6664
rect 0 6384 400 6440
rect 64600 6160 65000 6216
rect 0 5824 400 5880
rect 0 5264 400 5320
rect 0 4704 400 4760
rect 0 4144 400 4200
<< obsm3 >>
rect 400 60790 64666 64106
rect 430 60674 64666 60790
rect 400 60230 64666 60674
rect 430 60114 64666 60230
rect 400 59670 64666 60114
rect 430 59554 64666 59670
rect 400 59110 64666 59554
rect 430 58994 64666 59110
rect 400 58662 64666 58994
rect 400 58550 64570 58662
rect 430 58546 64570 58550
rect 430 58434 64666 58546
rect 400 58214 64666 58434
rect 400 58098 64570 58214
rect 400 57990 64666 58098
rect 430 57874 64666 57990
rect 400 57766 64666 57874
rect 400 57650 64570 57766
rect 400 57430 64666 57650
rect 430 57318 64666 57430
rect 430 57314 64570 57318
rect 400 57202 64570 57314
rect 400 56870 64666 57202
rect 430 56754 64570 56870
rect 400 56422 64666 56754
rect 400 56310 64570 56422
rect 430 56306 64570 56310
rect 430 56194 64666 56306
rect 400 55974 64666 56194
rect 400 55858 64570 55974
rect 400 55750 64666 55858
rect 430 55634 64666 55750
rect 400 55526 64666 55634
rect 400 55410 64570 55526
rect 400 55190 64666 55410
rect 430 55078 64666 55190
rect 430 55074 64570 55078
rect 400 54962 64570 55074
rect 400 54630 64666 54962
rect 430 54514 64570 54630
rect 400 54182 64666 54514
rect 400 54070 64570 54182
rect 430 54066 64570 54070
rect 430 53954 64666 54066
rect 400 53734 64666 53954
rect 400 53618 64570 53734
rect 400 53510 64666 53618
rect 430 53394 64666 53510
rect 400 53286 64666 53394
rect 400 53170 64570 53286
rect 400 52950 64666 53170
rect 430 52838 64666 52950
rect 430 52834 64570 52838
rect 400 52722 64570 52834
rect 400 52390 64666 52722
rect 430 52274 64570 52390
rect 400 51942 64666 52274
rect 400 51830 64570 51942
rect 430 51826 64570 51830
rect 430 51714 64666 51826
rect 400 51494 64666 51714
rect 400 51378 64570 51494
rect 400 51270 64666 51378
rect 430 51154 64666 51270
rect 400 51046 64666 51154
rect 400 50930 64570 51046
rect 400 50710 64666 50930
rect 430 50598 64666 50710
rect 430 50594 64570 50598
rect 400 50482 64570 50594
rect 400 50150 64666 50482
rect 430 50034 64570 50150
rect 400 49702 64666 50034
rect 400 49590 64570 49702
rect 430 49586 64570 49590
rect 430 49474 64666 49586
rect 400 49254 64666 49474
rect 400 49138 64570 49254
rect 400 49030 64666 49138
rect 430 48914 64666 49030
rect 400 48806 64666 48914
rect 400 48690 64570 48806
rect 400 48470 64666 48690
rect 430 48358 64666 48470
rect 430 48354 64570 48358
rect 400 48242 64570 48354
rect 400 47910 64666 48242
rect 430 47794 64570 47910
rect 400 47462 64666 47794
rect 400 47350 64570 47462
rect 430 47346 64570 47350
rect 430 47234 64666 47346
rect 400 47014 64666 47234
rect 400 46898 64570 47014
rect 400 46790 64666 46898
rect 430 46674 64666 46790
rect 400 46566 64666 46674
rect 400 46450 64570 46566
rect 400 46230 64666 46450
rect 430 46118 64666 46230
rect 430 46114 64570 46118
rect 400 46002 64570 46114
rect 400 45670 64666 46002
rect 430 45554 64570 45670
rect 400 45222 64666 45554
rect 400 45110 64570 45222
rect 430 45106 64570 45110
rect 430 44994 64666 45106
rect 400 44774 64666 44994
rect 400 44658 64570 44774
rect 400 44550 64666 44658
rect 430 44434 64666 44550
rect 400 44326 64666 44434
rect 400 44210 64570 44326
rect 400 43990 64666 44210
rect 430 43878 64666 43990
rect 430 43874 64570 43878
rect 400 43762 64570 43874
rect 400 43430 64666 43762
rect 430 43314 64570 43430
rect 400 42982 64666 43314
rect 400 42870 64570 42982
rect 430 42866 64570 42870
rect 430 42754 64666 42866
rect 400 42534 64666 42754
rect 400 42418 64570 42534
rect 400 42310 64666 42418
rect 430 42194 64666 42310
rect 400 42086 64666 42194
rect 400 41970 64570 42086
rect 400 41750 64666 41970
rect 430 41638 64666 41750
rect 430 41634 64570 41638
rect 400 41522 64570 41634
rect 400 41190 64666 41522
rect 430 41074 64570 41190
rect 400 40742 64666 41074
rect 400 40630 64570 40742
rect 430 40626 64570 40630
rect 430 40514 64666 40626
rect 400 40294 64666 40514
rect 400 40178 64570 40294
rect 400 40070 64666 40178
rect 430 39954 64666 40070
rect 400 39846 64666 39954
rect 400 39730 64570 39846
rect 400 39510 64666 39730
rect 430 39398 64666 39510
rect 430 39394 64570 39398
rect 400 39282 64570 39394
rect 400 38950 64666 39282
rect 430 38834 64570 38950
rect 400 38502 64666 38834
rect 400 38390 64570 38502
rect 430 38386 64570 38390
rect 430 38274 64666 38386
rect 400 38054 64666 38274
rect 400 37938 64570 38054
rect 400 37830 64666 37938
rect 430 37714 64666 37830
rect 400 37606 64666 37714
rect 400 37490 64570 37606
rect 400 37270 64666 37490
rect 430 37158 64666 37270
rect 430 37154 64570 37158
rect 400 37042 64570 37154
rect 400 36710 64666 37042
rect 430 36594 64570 36710
rect 400 36262 64666 36594
rect 400 36150 64570 36262
rect 430 36146 64570 36150
rect 430 36034 64666 36146
rect 400 35814 64666 36034
rect 400 35698 64570 35814
rect 400 35590 64666 35698
rect 430 35474 64666 35590
rect 400 35366 64666 35474
rect 400 35250 64570 35366
rect 400 35030 64666 35250
rect 430 34918 64666 35030
rect 430 34914 64570 34918
rect 400 34802 64570 34914
rect 400 34470 64666 34802
rect 430 34354 64570 34470
rect 400 34022 64666 34354
rect 400 33910 64570 34022
rect 430 33906 64570 33910
rect 430 33794 64666 33906
rect 400 33574 64666 33794
rect 400 33458 64570 33574
rect 400 33350 64666 33458
rect 430 33234 64666 33350
rect 400 33126 64666 33234
rect 400 33010 64570 33126
rect 400 32790 64666 33010
rect 430 32678 64666 32790
rect 430 32674 64570 32678
rect 400 32562 64570 32674
rect 400 32230 64666 32562
rect 430 32114 64570 32230
rect 400 31782 64666 32114
rect 400 31670 64570 31782
rect 430 31666 64570 31670
rect 430 31554 64666 31666
rect 400 31334 64666 31554
rect 400 31218 64570 31334
rect 400 31110 64666 31218
rect 430 30994 64666 31110
rect 400 30886 64666 30994
rect 400 30770 64570 30886
rect 400 30550 64666 30770
rect 430 30438 64666 30550
rect 430 30434 64570 30438
rect 400 30322 64570 30434
rect 400 29990 64666 30322
rect 430 29874 64570 29990
rect 400 29542 64666 29874
rect 400 29430 64570 29542
rect 430 29426 64570 29430
rect 430 29314 64666 29426
rect 400 29094 64666 29314
rect 400 28978 64570 29094
rect 400 28870 64666 28978
rect 430 28754 64666 28870
rect 400 28646 64666 28754
rect 400 28530 64570 28646
rect 400 28310 64666 28530
rect 430 28198 64666 28310
rect 430 28194 64570 28198
rect 400 28082 64570 28194
rect 400 27750 64666 28082
rect 430 27634 64570 27750
rect 400 27302 64666 27634
rect 400 27190 64570 27302
rect 430 27186 64570 27190
rect 430 27074 64666 27186
rect 400 26854 64666 27074
rect 400 26738 64570 26854
rect 400 26630 64666 26738
rect 430 26514 64666 26630
rect 400 26406 64666 26514
rect 400 26290 64570 26406
rect 400 26070 64666 26290
rect 430 25958 64666 26070
rect 430 25954 64570 25958
rect 400 25842 64570 25954
rect 400 25510 64666 25842
rect 430 25394 64570 25510
rect 400 25062 64666 25394
rect 400 24950 64570 25062
rect 430 24946 64570 24950
rect 430 24834 64666 24946
rect 400 24614 64666 24834
rect 400 24498 64570 24614
rect 400 24390 64666 24498
rect 430 24274 64666 24390
rect 400 24166 64666 24274
rect 400 24050 64570 24166
rect 400 23830 64666 24050
rect 430 23718 64666 23830
rect 430 23714 64570 23718
rect 400 23602 64570 23714
rect 400 23270 64666 23602
rect 430 23154 64570 23270
rect 400 22822 64666 23154
rect 400 22710 64570 22822
rect 430 22706 64570 22710
rect 430 22594 64666 22706
rect 400 22374 64666 22594
rect 400 22258 64570 22374
rect 400 22150 64666 22258
rect 430 22034 64666 22150
rect 400 21926 64666 22034
rect 400 21810 64570 21926
rect 400 21590 64666 21810
rect 430 21478 64666 21590
rect 430 21474 64570 21478
rect 400 21362 64570 21474
rect 400 21030 64666 21362
rect 430 20914 64570 21030
rect 400 20582 64666 20914
rect 400 20470 64570 20582
rect 430 20466 64570 20470
rect 430 20354 64666 20466
rect 400 20134 64666 20354
rect 400 20018 64570 20134
rect 400 19910 64666 20018
rect 430 19794 64666 19910
rect 400 19686 64666 19794
rect 400 19570 64570 19686
rect 400 19350 64666 19570
rect 430 19238 64666 19350
rect 430 19234 64570 19238
rect 400 19122 64570 19234
rect 400 18790 64666 19122
rect 430 18674 64570 18790
rect 400 18342 64666 18674
rect 400 18230 64570 18342
rect 430 18226 64570 18230
rect 430 18114 64666 18226
rect 400 17894 64666 18114
rect 400 17778 64570 17894
rect 400 17670 64666 17778
rect 430 17554 64666 17670
rect 400 17446 64666 17554
rect 400 17330 64570 17446
rect 400 17110 64666 17330
rect 430 16998 64666 17110
rect 430 16994 64570 16998
rect 400 16882 64570 16994
rect 400 16550 64666 16882
rect 430 16434 64570 16550
rect 400 16102 64666 16434
rect 400 15990 64570 16102
rect 430 15986 64570 15990
rect 430 15874 64666 15986
rect 400 15654 64666 15874
rect 400 15538 64570 15654
rect 400 15430 64666 15538
rect 430 15314 64666 15430
rect 400 15206 64666 15314
rect 400 15090 64570 15206
rect 400 14870 64666 15090
rect 430 14758 64666 14870
rect 430 14754 64570 14758
rect 400 14642 64570 14754
rect 400 14310 64666 14642
rect 430 14194 64570 14310
rect 400 13862 64666 14194
rect 400 13750 64570 13862
rect 430 13746 64570 13750
rect 430 13634 64666 13746
rect 400 13414 64666 13634
rect 400 13298 64570 13414
rect 400 13190 64666 13298
rect 430 13074 64666 13190
rect 400 12966 64666 13074
rect 400 12850 64570 12966
rect 400 12630 64666 12850
rect 430 12518 64666 12630
rect 430 12514 64570 12518
rect 400 12402 64570 12514
rect 400 12070 64666 12402
rect 430 11954 64570 12070
rect 400 11622 64666 11954
rect 400 11510 64570 11622
rect 430 11506 64570 11510
rect 430 11394 64666 11506
rect 400 11174 64666 11394
rect 400 11058 64570 11174
rect 400 10950 64666 11058
rect 430 10834 64666 10950
rect 400 10726 64666 10834
rect 400 10610 64570 10726
rect 400 10390 64666 10610
rect 430 10278 64666 10390
rect 430 10274 64570 10278
rect 400 10162 64570 10274
rect 400 9830 64666 10162
rect 430 9714 64570 9830
rect 400 9382 64666 9714
rect 400 9270 64570 9382
rect 430 9266 64570 9270
rect 430 9154 64666 9266
rect 400 8934 64666 9154
rect 400 8818 64570 8934
rect 400 8710 64666 8818
rect 430 8594 64666 8710
rect 400 8486 64666 8594
rect 400 8370 64570 8486
rect 400 8150 64666 8370
rect 430 8038 64666 8150
rect 430 8034 64570 8038
rect 400 7922 64570 8034
rect 400 7590 64666 7922
rect 430 7474 64570 7590
rect 400 7142 64666 7474
rect 400 7030 64570 7142
rect 430 7026 64570 7030
rect 430 6914 64666 7026
rect 400 6694 64666 6914
rect 400 6578 64570 6694
rect 400 6470 64666 6578
rect 430 6354 64666 6470
rect 400 6246 64666 6354
rect 400 6130 64570 6246
rect 400 5910 64666 6130
rect 430 5794 64666 5910
rect 400 5350 64666 5794
rect 430 5234 64666 5350
rect 400 4790 64666 5234
rect 430 4674 64666 4790
rect 400 4230 64666 4674
rect 430 4114 64666 4230
rect 400 1470 64666 4114
<< metal4 >>
rect 2224 1538 2384 63142
rect 9904 1538 10064 63142
rect 17584 1538 17744 63142
rect 25264 1538 25424 63142
rect 32944 1538 33104 63142
rect 40624 1538 40784 63142
rect 48304 1538 48464 63142
rect 55984 1538 56144 63142
rect 63664 1538 63824 63142
<< obsm4 >>
rect 10150 1633 17554 62879
rect 17774 1633 25234 62879
rect 25454 1633 32914 62879
rect 33134 1633 40594 62879
rect 40814 1633 48274 62879
rect 48494 1633 55954 62879
rect 56174 1633 63154 62879
<< labels >>
rlabel metal2 s 48496 64600 48552 65000 6 ay8913_do[0]
port 1 nsew signal input
rlabel metal2 s 52976 64600 53032 65000 6 ay8913_do[10]
port 2 nsew signal input
rlabel metal2 s 53424 64600 53480 65000 6 ay8913_do[11]
port 3 nsew signal input
rlabel metal2 s 53872 64600 53928 65000 6 ay8913_do[12]
port 4 nsew signal input
rlabel metal2 s 54320 64600 54376 65000 6 ay8913_do[13]
port 5 nsew signal input
rlabel metal2 s 54768 64600 54824 65000 6 ay8913_do[14]
port 6 nsew signal input
rlabel metal2 s 55216 64600 55272 65000 6 ay8913_do[15]
port 7 nsew signal input
rlabel metal2 s 55664 64600 55720 65000 6 ay8913_do[16]
port 8 nsew signal input
rlabel metal2 s 56112 64600 56168 65000 6 ay8913_do[17]
port 9 nsew signal input
rlabel metal2 s 56560 64600 56616 65000 6 ay8913_do[18]
port 10 nsew signal input
rlabel metal2 s 57008 64600 57064 65000 6 ay8913_do[19]
port 11 nsew signal input
rlabel metal2 s 48944 64600 49000 65000 6 ay8913_do[1]
port 12 nsew signal input
rlabel metal2 s 57456 64600 57512 65000 6 ay8913_do[20]
port 13 nsew signal input
rlabel metal2 s 57904 64600 57960 65000 6 ay8913_do[21]
port 14 nsew signal input
rlabel metal2 s 58352 64600 58408 65000 6 ay8913_do[22]
port 15 nsew signal input
rlabel metal2 s 58800 64600 58856 65000 6 ay8913_do[23]
port 16 nsew signal input
rlabel metal2 s 59248 64600 59304 65000 6 ay8913_do[24]
port 17 nsew signal input
rlabel metal2 s 59696 64600 59752 65000 6 ay8913_do[25]
port 18 nsew signal input
rlabel metal2 s 60144 64600 60200 65000 6 ay8913_do[26]
port 19 nsew signal input
rlabel metal2 s 60592 64600 60648 65000 6 ay8913_do[27]
port 20 nsew signal input
rlabel metal2 s 49392 64600 49448 65000 6 ay8913_do[2]
port 21 nsew signal input
rlabel metal2 s 49840 64600 49896 65000 6 ay8913_do[3]
port 22 nsew signal input
rlabel metal2 s 50288 64600 50344 65000 6 ay8913_do[4]
port 23 nsew signal input
rlabel metal2 s 50736 64600 50792 65000 6 ay8913_do[5]
port 24 nsew signal input
rlabel metal2 s 51184 64600 51240 65000 6 ay8913_do[6]
port 25 nsew signal input
rlabel metal2 s 51632 64600 51688 65000 6 ay8913_do[7]
port 26 nsew signal input
rlabel metal2 s 52080 64600 52136 65000 6 ay8913_do[8]
port 27 nsew signal input
rlabel metal2 s 52528 64600 52584 65000 6 ay8913_do[9]
port 28 nsew signal input
rlabel metal2 s 39984 64600 40040 65000 6 blinker_do[0]
port 29 nsew signal input
rlabel metal2 s 40432 64600 40488 65000 6 blinker_do[1]
port 30 nsew signal input
rlabel metal2 s 40880 64600 40936 65000 6 blinker_do[2]
port 31 nsew signal input
rlabel metal3 s 64600 22288 65000 22344 6 custom_settings[0]
port 32 nsew signal output
rlabel metal3 s 64600 26768 65000 26824 6 custom_settings[10]
port 33 nsew signal output
rlabel metal3 s 64600 27216 65000 27272 6 custom_settings[11]
port 34 nsew signal output
rlabel metal3 s 64600 27664 65000 27720 6 custom_settings[12]
port 35 nsew signal output
rlabel metal3 s 64600 28112 65000 28168 6 custom_settings[13]
port 36 nsew signal output
rlabel metal3 s 64600 28560 65000 28616 6 custom_settings[14]
port 37 nsew signal output
rlabel metal3 s 64600 29008 65000 29064 6 custom_settings[15]
port 38 nsew signal output
rlabel metal3 s 64600 29456 65000 29512 6 custom_settings[16]
port 39 nsew signal output
rlabel metal3 s 64600 29904 65000 29960 6 custom_settings[17]
port 40 nsew signal output
rlabel metal3 s 64600 30352 65000 30408 6 custom_settings[18]
port 41 nsew signal output
rlabel metal3 s 64600 30800 65000 30856 6 custom_settings[19]
port 42 nsew signal output
rlabel metal3 s 64600 22736 65000 22792 6 custom_settings[1]
port 43 nsew signal output
rlabel metal3 s 64600 31248 65000 31304 6 custom_settings[20]
port 44 nsew signal output
rlabel metal3 s 64600 31696 65000 31752 6 custom_settings[21]
port 45 nsew signal output
rlabel metal3 s 64600 32144 65000 32200 6 custom_settings[22]
port 46 nsew signal output
rlabel metal3 s 64600 32592 65000 32648 6 custom_settings[23]
port 47 nsew signal output
rlabel metal3 s 64600 33040 65000 33096 6 custom_settings[24]
port 48 nsew signal output
rlabel metal3 s 64600 33488 65000 33544 6 custom_settings[25]
port 49 nsew signal output
rlabel metal3 s 64600 33936 65000 33992 6 custom_settings[26]
port 50 nsew signal output
rlabel metal3 s 64600 34384 65000 34440 6 custom_settings[27]
port 51 nsew signal output
rlabel metal3 s 64600 34832 65000 34888 6 custom_settings[28]
port 52 nsew signal output
rlabel metal3 s 64600 35280 65000 35336 6 custom_settings[29]
port 53 nsew signal output
rlabel metal3 s 64600 23184 65000 23240 6 custom_settings[2]
port 54 nsew signal output
rlabel metal3 s 64600 35728 65000 35784 6 custom_settings[30]
port 55 nsew signal output
rlabel metal3 s 64600 36176 65000 36232 6 custom_settings[31]
port 56 nsew signal output
rlabel metal3 s 64600 23632 65000 23688 6 custom_settings[3]
port 57 nsew signal output
rlabel metal3 s 64600 24080 65000 24136 6 custom_settings[4]
port 58 nsew signal output
rlabel metal3 s 64600 24528 65000 24584 6 custom_settings[5]
port 59 nsew signal output
rlabel metal3 s 64600 24976 65000 25032 6 custom_settings[6]
port 60 nsew signal output
rlabel metal3 s 64600 25424 65000 25480 6 custom_settings[7]
port 61 nsew signal output
rlabel metal3 s 64600 25872 65000 25928 6 custom_settings[8]
port 62 nsew signal output
rlabel metal3 s 64600 26320 65000 26376 6 custom_settings[9]
port 63 nsew signal output
rlabel metal3 s 0 57344 400 57400 6 hellorld_do
port 64 nsew signal input
rlabel metal2 s 4144 64600 4200 65000 6 io_in[0]
port 65 nsew signal input
rlabel metal2 s 8624 64600 8680 65000 6 io_in[10]
port 66 nsew signal input
rlabel metal2 s 9072 64600 9128 65000 6 io_in[11]
port 67 nsew signal input
rlabel metal2 s 9520 64600 9576 65000 6 io_in[12]
port 68 nsew signal input
rlabel metal2 s 9968 64600 10024 65000 6 io_in[13]
port 69 nsew signal input
rlabel metal2 s 10416 64600 10472 65000 6 io_in[14]
port 70 nsew signal input
rlabel metal2 s 10864 64600 10920 65000 6 io_in[15]
port 71 nsew signal input
rlabel metal2 s 11312 64600 11368 65000 6 io_in[16]
port 72 nsew signal input
rlabel metal2 s 11760 64600 11816 65000 6 io_in[17]
port 73 nsew signal input
rlabel metal2 s 12208 64600 12264 65000 6 io_in[18]
port 74 nsew signal input
rlabel metal2 s 12656 64600 12712 65000 6 io_in[19]
port 75 nsew signal input
rlabel metal2 s 4592 64600 4648 65000 6 io_in[1]
port 76 nsew signal input
rlabel metal2 s 13104 64600 13160 65000 6 io_in[20]
port 77 nsew signal input
rlabel metal2 s 13552 64600 13608 65000 6 io_in[21]
port 78 nsew signal input
rlabel metal2 s 14000 64600 14056 65000 6 io_in[22]
port 79 nsew signal input
rlabel metal2 s 14448 64600 14504 65000 6 io_in[23]
port 80 nsew signal input
rlabel metal2 s 14896 64600 14952 65000 6 io_in[24]
port 81 nsew signal input
rlabel metal2 s 15344 64600 15400 65000 6 io_in[25]
port 82 nsew signal input
rlabel metal2 s 15792 64600 15848 65000 6 io_in[26]
port 83 nsew signal input
rlabel metal2 s 16240 64600 16296 65000 6 io_in[27]
port 84 nsew signal input
rlabel metal2 s 16688 64600 16744 65000 6 io_in[28]
port 85 nsew signal input
rlabel metal2 s 17136 64600 17192 65000 6 io_in[29]
port 86 nsew signal input
rlabel metal2 s 5040 64600 5096 65000 6 io_in[2]
port 87 nsew signal input
rlabel metal2 s 17584 64600 17640 65000 6 io_in[30]
port 88 nsew signal input
rlabel metal2 s 18032 64600 18088 65000 6 io_in[31]
port 89 nsew signal input
rlabel metal2 s 18480 64600 18536 65000 6 io_in[32]
port 90 nsew signal input
rlabel metal2 s 18928 64600 18984 65000 6 io_in[33]
port 91 nsew signal input
rlabel metal2 s 19376 64600 19432 65000 6 io_in[34]
port 92 nsew signal input
rlabel metal2 s 19824 64600 19880 65000 6 io_in[35]
port 93 nsew signal input
rlabel metal2 s 20272 64600 20328 65000 6 io_in[36]
port 94 nsew signal input
rlabel metal2 s 20720 64600 20776 65000 6 io_in[37]
port 95 nsew signal input
rlabel metal2 s 5488 64600 5544 65000 6 io_in[3]
port 96 nsew signal input
rlabel metal2 s 5936 64600 5992 65000 6 io_in[4]
port 97 nsew signal input
rlabel metal2 s 6384 64600 6440 65000 6 io_in[5]
port 98 nsew signal input
rlabel metal2 s 6832 64600 6888 65000 6 io_in[6]
port 99 nsew signal input
rlabel metal2 s 7280 64600 7336 65000 6 io_in[7]
port 100 nsew signal input
rlabel metal2 s 7728 64600 7784 65000 6 io_in[8]
port 101 nsew signal input
rlabel metal2 s 8176 64600 8232 65000 6 io_in[9]
port 102 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 io_oeb[0]
port 103 nsew signal output
rlabel metal3 s 0 9744 400 9800 6 io_oeb[10]
port 104 nsew signal output
rlabel metal3 s 0 10304 400 10360 6 io_oeb[11]
port 105 nsew signal output
rlabel metal3 s 0 10864 400 10920 6 io_oeb[12]
port 106 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 io_oeb[13]
port 107 nsew signal output
rlabel metal3 s 0 11984 400 12040 6 io_oeb[14]
port 108 nsew signal output
rlabel metal3 s 0 12544 400 12600 6 io_oeb[15]
port 109 nsew signal output
rlabel metal3 s 0 13104 400 13160 6 io_oeb[16]
port 110 nsew signal output
rlabel metal3 s 0 13664 400 13720 6 io_oeb[17]
port 111 nsew signal output
rlabel metal3 s 0 14224 400 14280 6 io_oeb[18]
port 112 nsew signal output
rlabel metal3 s 0 14784 400 14840 6 io_oeb[19]
port 113 nsew signal output
rlabel metal3 s 0 4704 400 4760 6 io_oeb[1]
port 114 nsew signal output
rlabel metal3 s 0 15344 400 15400 6 io_oeb[20]
port 115 nsew signal output
rlabel metal3 s 0 15904 400 15960 6 io_oeb[21]
port 116 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 io_oeb[22]
port 117 nsew signal output
rlabel metal3 s 0 17024 400 17080 6 io_oeb[23]
port 118 nsew signal output
rlabel metal3 s 0 17584 400 17640 6 io_oeb[24]
port 119 nsew signal output
rlabel metal3 s 0 18144 400 18200 6 io_oeb[25]
port 120 nsew signal output
rlabel metal3 s 0 18704 400 18760 6 io_oeb[26]
port 121 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 io_oeb[27]
port 122 nsew signal output
rlabel metal3 s 0 19824 400 19880 6 io_oeb[28]
port 123 nsew signal output
rlabel metal3 s 0 20384 400 20440 6 io_oeb[29]
port 124 nsew signal output
rlabel metal3 s 0 5264 400 5320 6 io_oeb[2]
port 125 nsew signal output
rlabel metal3 s 0 20944 400 21000 6 io_oeb[30]
port 126 nsew signal output
rlabel metal3 s 0 21504 400 21560 6 io_oeb[31]
port 127 nsew signal output
rlabel metal3 s 0 22064 400 22120 6 io_oeb[32]
port 128 nsew signal output
rlabel metal3 s 0 22624 400 22680 6 io_oeb[33]
port 129 nsew signal output
rlabel metal3 s 0 23184 400 23240 6 io_oeb[34]
port 130 nsew signal output
rlabel metal3 s 0 23744 400 23800 6 io_oeb[35]
port 131 nsew signal output
rlabel metal3 s 0 24304 400 24360 6 io_oeb[36]
port 132 nsew signal output
rlabel metal3 s 0 24864 400 24920 6 io_oeb[37]
port 133 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 io_oeb[3]
port 134 nsew signal output
rlabel metal3 s 0 6384 400 6440 6 io_oeb[4]
port 135 nsew signal output
rlabel metal3 s 0 6944 400 7000 6 io_oeb[5]
port 136 nsew signal output
rlabel metal3 s 0 7504 400 7560 6 io_oeb[6]
port 137 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 io_oeb[7]
port 138 nsew signal output
rlabel metal3 s 0 8624 400 8680 6 io_oeb[8]
port 139 nsew signal output
rlabel metal3 s 0 9184 400 9240 6 io_oeb[9]
port 140 nsew signal output
rlabel metal2 s 21168 64600 21224 65000 6 io_out[0]
port 141 nsew signal output
rlabel metal2 s 25648 64600 25704 65000 6 io_out[10]
port 142 nsew signal output
rlabel metal2 s 26096 64600 26152 65000 6 io_out[11]
port 143 nsew signal output
rlabel metal2 s 26544 64600 26600 65000 6 io_out[12]
port 144 nsew signal output
rlabel metal2 s 26992 64600 27048 65000 6 io_out[13]
port 145 nsew signal output
rlabel metal2 s 27440 64600 27496 65000 6 io_out[14]
port 146 nsew signal output
rlabel metal2 s 27888 64600 27944 65000 6 io_out[15]
port 147 nsew signal output
rlabel metal2 s 28336 64600 28392 65000 6 io_out[16]
port 148 nsew signal output
rlabel metal2 s 28784 64600 28840 65000 6 io_out[17]
port 149 nsew signal output
rlabel metal2 s 29232 64600 29288 65000 6 io_out[18]
port 150 nsew signal output
rlabel metal2 s 29680 64600 29736 65000 6 io_out[19]
port 151 nsew signal output
rlabel metal2 s 21616 64600 21672 65000 6 io_out[1]
port 152 nsew signal output
rlabel metal2 s 30128 64600 30184 65000 6 io_out[20]
port 153 nsew signal output
rlabel metal2 s 30576 64600 30632 65000 6 io_out[21]
port 154 nsew signal output
rlabel metal2 s 31024 64600 31080 65000 6 io_out[22]
port 155 nsew signal output
rlabel metal2 s 31472 64600 31528 65000 6 io_out[23]
port 156 nsew signal output
rlabel metal2 s 31920 64600 31976 65000 6 io_out[24]
port 157 nsew signal output
rlabel metal2 s 32368 64600 32424 65000 6 io_out[25]
port 158 nsew signal output
rlabel metal2 s 32816 64600 32872 65000 6 io_out[26]
port 159 nsew signal output
rlabel metal2 s 33264 64600 33320 65000 6 io_out[27]
port 160 nsew signal output
rlabel metal2 s 33712 64600 33768 65000 6 io_out[28]
port 161 nsew signal output
rlabel metal2 s 34160 64600 34216 65000 6 io_out[29]
port 162 nsew signal output
rlabel metal2 s 22064 64600 22120 65000 6 io_out[2]
port 163 nsew signal output
rlabel metal2 s 34608 64600 34664 65000 6 io_out[30]
port 164 nsew signal output
rlabel metal2 s 35056 64600 35112 65000 6 io_out[31]
port 165 nsew signal output
rlabel metal2 s 35504 64600 35560 65000 6 io_out[32]
port 166 nsew signal output
rlabel metal2 s 35952 64600 36008 65000 6 io_out[33]
port 167 nsew signal output
rlabel metal2 s 36400 64600 36456 65000 6 io_out[34]
port 168 nsew signal output
rlabel metal2 s 36848 64600 36904 65000 6 io_out[35]
port 169 nsew signal output
rlabel metal2 s 37296 64600 37352 65000 6 io_out[36]
port 170 nsew signal output
rlabel metal2 s 37744 64600 37800 65000 6 io_out[37]
port 171 nsew signal output
rlabel metal2 s 22512 64600 22568 65000 6 io_out[3]
port 172 nsew signal output
rlabel metal2 s 22960 64600 23016 65000 6 io_out[4]
port 173 nsew signal output
rlabel metal2 s 23408 64600 23464 65000 6 io_out[5]
port 174 nsew signal output
rlabel metal2 s 23856 64600 23912 65000 6 io_out[6]
port 175 nsew signal output
rlabel metal2 s 24304 64600 24360 65000 6 io_out[7]
port 176 nsew signal output
rlabel metal2 s 24752 64600 24808 65000 6 io_out[8]
port 177 nsew signal output
rlabel metal2 s 25200 64600 25256 65000 6 io_out[9]
port 178 nsew signal output
rlabel metal2 s 38192 64600 38248 65000 6 irq[0]
port 179 nsew signal output
rlabel metal2 s 38640 64600 38696 65000 6 irq[1]
port 180 nsew signal output
rlabel metal2 s 39088 64600 39144 65000 6 irq[2]
port 181 nsew signal output
rlabel metal3 s 0 39424 400 39480 6 mc14500_do[0]
port 182 nsew signal input
rlabel metal3 s 0 45024 400 45080 6 mc14500_do[10]
port 183 nsew signal input
rlabel metal3 s 0 45584 400 45640 6 mc14500_do[11]
port 184 nsew signal input
rlabel metal3 s 0 46144 400 46200 6 mc14500_do[12]
port 185 nsew signal input
rlabel metal3 s 0 46704 400 46760 6 mc14500_do[13]
port 186 nsew signal input
rlabel metal3 s 0 47264 400 47320 6 mc14500_do[14]
port 187 nsew signal input
rlabel metal3 s 0 47824 400 47880 6 mc14500_do[15]
port 188 nsew signal input
rlabel metal3 s 0 48384 400 48440 6 mc14500_do[16]
port 189 nsew signal input
rlabel metal3 s 0 48944 400 49000 6 mc14500_do[17]
port 190 nsew signal input
rlabel metal3 s 0 49504 400 49560 6 mc14500_do[18]
port 191 nsew signal input
rlabel metal3 s 0 50064 400 50120 6 mc14500_do[19]
port 192 nsew signal input
rlabel metal3 s 0 39984 400 40040 6 mc14500_do[1]
port 193 nsew signal input
rlabel metal3 s 0 50624 400 50680 6 mc14500_do[20]
port 194 nsew signal input
rlabel metal3 s 0 51184 400 51240 6 mc14500_do[21]
port 195 nsew signal input
rlabel metal3 s 0 51744 400 51800 6 mc14500_do[22]
port 196 nsew signal input
rlabel metal3 s 0 52304 400 52360 6 mc14500_do[23]
port 197 nsew signal input
rlabel metal3 s 0 52864 400 52920 6 mc14500_do[24]
port 198 nsew signal input
rlabel metal3 s 0 53424 400 53480 6 mc14500_do[25]
port 199 nsew signal input
rlabel metal3 s 0 53984 400 54040 6 mc14500_do[26]
port 200 nsew signal input
rlabel metal3 s 0 54544 400 54600 6 mc14500_do[27]
port 201 nsew signal input
rlabel metal3 s 0 55104 400 55160 6 mc14500_do[28]
port 202 nsew signal input
rlabel metal3 s 0 55664 400 55720 6 mc14500_do[29]
port 203 nsew signal input
rlabel metal3 s 0 40544 400 40600 6 mc14500_do[2]
port 204 nsew signal input
rlabel metal3 s 0 56224 400 56280 6 mc14500_do[30]
port 205 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 mc14500_do[3]
port 206 nsew signal input
rlabel metal3 s 0 41664 400 41720 6 mc14500_do[4]
port 207 nsew signal input
rlabel metal3 s 0 42224 400 42280 6 mc14500_do[5]
port 208 nsew signal input
rlabel metal3 s 0 42784 400 42840 6 mc14500_do[6]
port 209 nsew signal input
rlabel metal3 s 0 43344 400 43400 6 mc14500_do[7]
port 210 nsew signal input
rlabel metal3 s 0 43904 400 43960 6 mc14500_do[8]
port 211 nsew signal input
rlabel metal3 s 0 44464 400 44520 6 mc14500_do[9]
port 212 nsew signal input
rlabel metal2 s 41776 64600 41832 65000 6 mc14500_sram_addr[0]
port 213 nsew signal input
rlabel metal2 s 42224 64600 42280 65000 6 mc14500_sram_addr[1]
port 214 nsew signal input
rlabel metal2 s 42672 64600 42728 65000 6 mc14500_sram_addr[2]
port 215 nsew signal input
rlabel metal2 s 43120 64600 43176 65000 6 mc14500_sram_addr[3]
port 216 nsew signal input
rlabel metal2 s 43568 64600 43624 65000 6 mc14500_sram_addr[4]
port 217 nsew signal input
rlabel metal2 s 44016 64600 44072 65000 6 mc14500_sram_addr[5]
port 218 nsew signal input
rlabel metal2 s 48048 64600 48104 65000 6 mc14500_sram_gwe
port 219 nsew signal input
rlabel metal2 s 44464 64600 44520 65000 6 mc14500_sram_in[0]
port 220 nsew signal input
rlabel metal2 s 44912 64600 44968 65000 6 mc14500_sram_in[1]
port 221 nsew signal input
rlabel metal2 s 45360 64600 45416 65000 6 mc14500_sram_in[2]
port 222 nsew signal input
rlabel metal2 s 45808 64600 45864 65000 6 mc14500_sram_in[3]
port 223 nsew signal input
rlabel metal2 s 46256 64600 46312 65000 6 mc14500_sram_in[4]
port 224 nsew signal input
rlabel metal2 s 46704 64600 46760 65000 6 mc14500_sram_in[5]
port 225 nsew signal input
rlabel metal2 s 47152 64600 47208 65000 6 mc14500_sram_in[6]
port 226 nsew signal input
rlabel metal2 s 47600 64600 47656 65000 6 mc14500_sram_in[7]
port 227 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 qcpu_do[0]
port 228 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 qcpu_do[10]
port 229 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 qcpu_do[11]
port 230 nsew signal input
rlabel metal2 s 50064 0 50120 400 6 qcpu_do[12]
port 231 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 qcpu_do[13]
port 232 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 qcpu_do[14]
port 233 nsew signal input
rlabel metal2 s 51408 0 51464 400 6 qcpu_do[15]
port 234 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 qcpu_do[16]
port 235 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 qcpu_do[17]
port 236 nsew signal input
rlabel metal2 s 52752 0 52808 400 6 qcpu_do[18]
port 237 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 qcpu_do[19]
port 238 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 qcpu_do[1]
port 239 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 qcpu_do[20]
port 240 nsew signal input
rlabel metal2 s 54096 0 54152 400 6 qcpu_do[21]
port 241 nsew signal input
rlabel metal2 s 54544 0 54600 400 6 qcpu_do[22]
port 242 nsew signal input
rlabel metal2 s 54992 0 55048 400 6 qcpu_do[23]
port 243 nsew signal input
rlabel metal2 s 55440 0 55496 400 6 qcpu_do[24]
port 244 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 qcpu_do[25]
port 245 nsew signal input
rlabel metal2 s 56336 0 56392 400 6 qcpu_do[26]
port 246 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 qcpu_do[27]
port 247 nsew signal input
rlabel metal2 s 57232 0 57288 400 6 qcpu_do[28]
port 248 nsew signal input
rlabel metal2 s 57680 0 57736 400 6 qcpu_do[29]
port 249 nsew signal input
rlabel metal2 s 45584 0 45640 400 6 qcpu_do[2]
port 250 nsew signal input
rlabel metal2 s 58128 0 58184 400 6 qcpu_do[30]
port 251 nsew signal input
rlabel metal2 s 58576 0 58632 400 6 qcpu_do[31]
port 252 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 qcpu_do[32]
port 253 nsew signal input
rlabel metal2 s 46032 0 46088 400 6 qcpu_do[3]
port 254 nsew signal input
rlabel metal2 s 46480 0 46536 400 6 qcpu_do[4]
port 255 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 qcpu_do[5]
port 256 nsew signal input
rlabel metal2 s 47376 0 47432 400 6 qcpu_do[6]
port 257 nsew signal input
rlabel metal2 s 47824 0 47880 400 6 qcpu_do[7]
port 258 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 qcpu_do[8]
port 259 nsew signal input
rlabel metal2 s 48720 0 48776 400 6 qcpu_do[9]
port 260 nsew signal input
rlabel metal3 s 64600 36624 65000 36680 6 qcpu_oeb[0]
port 261 nsew signal input
rlabel metal3 s 64600 41104 65000 41160 6 qcpu_oeb[10]
port 262 nsew signal input
rlabel metal3 s 64600 41552 65000 41608 6 qcpu_oeb[11]
port 263 nsew signal input
rlabel metal3 s 64600 42000 65000 42056 6 qcpu_oeb[12]
port 264 nsew signal input
rlabel metal3 s 64600 42448 65000 42504 6 qcpu_oeb[13]
port 265 nsew signal input
rlabel metal3 s 64600 42896 65000 42952 6 qcpu_oeb[14]
port 266 nsew signal input
rlabel metal3 s 64600 43344 65000 43400 6 qcpu_oeb[15]
port 267 nsew signal input
rlabel metal3 s 64600 43792 65000 43848 6 qcpu_oeb[16]
port 268 nsew signal input
rlabel metal3 s 64600 44240 65000 44296 6 qcpu_oeb[17]
port 269 nsew signal input
rlabel metal3 s 64600 44688 65000 44744 6 qcpu_oeb[18]
port 270 nsew signal input
rlabel metal3 s 64600 45136 65000 45192 6 qcpu_oeb[19]
port 271 nsew signal input
rlabel metal3 s 64600 37072 65000 37128 6 qcpu_oeb[1]
port 272 nsew signal input
rlabel metal3 s 64600 45584 65000 45640 6 qcpu_oeb[20]
port 273 nsew signal input
rlabel metal3 s 64600 46032 65000 46088 6 qcpu_oeb[21]
port 274 nsew signal input
rlabel metal3 s 64600 46480 65000 46536 6 qcpu_oeb[22]
port 275 nsew signal input
rlabel metal3 s 64600 46928 65000 46984 6 qcpu_oeb[23]
port 276 nsew signal input
rlabel metal3 s 64600 47376 65000 47432 6 qcpu_oeb[24]
port 277 nsew signal input
rlabel metal3 s 64600 47824 65000 47880 6 qcpu_oeb[25]
port 278 nsew signal input
rlabel metal3 s 64600 48272 65000 48328 6 qcpu_oeb[26]
port 279 nsew signal input
rlabel metal3 s 64600 48720 65000 48776 6 qcpu_oeb[27]
port 280 nsew signal input
rlabel metal3 s 64600 49168 65000 49224 6 qcpu_oeb[28]
port 281 nsew signal input
rlabel metal3 s 64600 49616 65000 49672 6 qcpu_oeb[29]
port 282 nsew signal input
rlabel metal3 s 64600 37520 65000 37576 6 qcpu_oeb[2]
port 283 nsew signal input
rlabel metal3 s 64600 50064 65000 50120 6 qcpu_oeb[30]
port 284 nsew signal input
rlabel metal3 s 64600 50512 65000 50568 6 qcpu_oeb[31]
port 285 nsew signal input
rlabel metal3 s 64600 50960 65000 51016 6 qcpu_oeb[32]
port 286 nsew signal input
rlabel metal3 s 64600 37968 65000 38024 6 qcpu_oeb[3]
port 287 nsew signal input
rlabel metal3 s 64600 38416 65000 38472 6 qcpu_oeb[4]
port 288 nsew signal input
rlabel metal3 s 64600 38864 65000 38920 6 qcpu_oeb[5]
port 289 nsew signal input
rlabel metal3 s 64600 39312 65000 39368 6 qcpu_oeb[6]
port 290 nsew signal input
rlabel metal3 s 64600 39760 65000 39816 6 qcpu_oeb[7]
port 291 nsew signal input
rlabel metal3 s 64600 40208 65000 40264 6 qcpu_oeb[8]
port 292 nsew signal input
rlabel metal3 s 64600 40656 65000 40712 6 qcpu_oeb[9]
port 293 nsew signal input
rlabel metal2 s 59472 0 59528 400 6 qcpu_sram_addr[0]
port 294 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 qcpu_sram_addr[1]
port 295 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 qcpu_sram_addr[2]
port 296 nsew signal input
rlabel metal2 s 60816 0 60872 400 6 qcpu_sram_addr[3]
port 297 nsew signal input
rlabel metal2 s 61264 0 61320 400 6 qcpu_sram_addr[4]
port 298 nsew signal input
rlabel metal2 s 61712 0 61768 400 6 qcpu_sram_addr[5]
port 299 nsew signal input
rlabel metal2 s 62160 0 62216 400 6 qcpu_sram_gwe
port 300 nsew signal input
rlabel metal3 s 64600 51408 65000 51464 6 qcpu_sram_in[0]
port 301 nsew signal input
rlabel metal3 s 64600 51856 65000 51912 6 qcpu_sram_in[1]
port 302 nsew signal input
rlabel metal3 s 64600 52304 65000 52360 6 qcpu_sram_in[2]
port 303 nsew signal input
rlabel metal3 s 64600 52752 65000 52808 6 qcpu_sram_in[3]
port 304 nsew signal input
rlabel metal3 s 64600 53200 65000 53256 6 qcpu_sram_in[4]
port 305 nsew signal input
rlabel metal3 s 64600 53648 65000 53704 6 qcpu_sram_in[5]
port 306 nsew signal input
rlabel metal3 s 64600 54096 65000 54152 6 qcpu_sram_in[6]
port 307 nsew signal input
rlabel metal3 s 64600 54544 65000 54600 6 qcpu_sram_in[7]
port 308 nsew signal input
rlabel metal3 s 64600 54992 65000 55048 6 qcpu_sram_out[0]
port 309 nsew signal output
rlabel metal3 s 64600 55440 65000 55496 6 qcpu_sram_out[1]
port 310 nsew signal output
rlabel metal3 s 64600 55888 65000 55944 6 qcpu_sram_out[2]
port 311 nsew signal output
rlabel metal3 s 64600 56336 65000 56392 6 qcpu_sram_out[3]
port 312 nsew signal output
rlabel metal3 s 64600 56784 65000 56840 6 qcpu_sram_out[4]
port 313 nsew signal output
rlabel metal3 s 64600 57232 65000 57288 6 qcpu_sram_out[5]
port 314 nsew signal output
rlabel metal3 s 64600 57680 65000 57736 6 qcpu_sram_out[6]
port 315 nsew signal output
rlabel metal3 s 64600 58128 65000 58184 6 qcpu_sram_out[7]
port 316 nsew signal output
rlabel metal3 s 64600 58576 65000 58632 6 rst_ay8913
port 317 nsew signal output
rlabel metal2 s 39536 64600 39592 65000 6 rst_blinker
port 318 nsew signal output
rlabel metal3 s 0 56784 400 56840 6 rst_hellorld
port 319 nsew signal output
rlabel metal3 s 0 38864 400 38920 6 rst_mc14500
port 320 nsew signal output
rlabel metal3 s 0 38304 400 38360 6 rst_qcpu
port 321 nsew signal output
rlabel metal3 s 0 25424 400 25480 6 rst_sid
port 322 nsew signal output
rlabel metal2 s 41328 64600 41384 65000 6 rst_sn76489
port 323 nsew signal output
rlabel metal3 s 0 57904 400 57960 6 rst_tbb1143
port 324 nsew signal output
rlabel metal3 s 0 25984 400 26040 6 sid_do[0]
port 325 nsew signal input
rlabel metal3 s 0 31584 400 31640 6 sid_do[10]
port 326 nsew signal input
rlabel metal3 s 0 32144 400 32200 6 sid_do[11]
port 327 nsew signal input
rlabel metal3 s 0 32704 400 32760 6 sid_do[12]
port 328 nsew signal input
rlabel metal3 s 0 33264 400 33320 6 sid_do[13]
port 329 nsew signal input
rlabel metal3 s 0 33824 400 33880 6 sid_do[14]
port 330 nsew signal input
rlabel metal3 s 0 34384 400 34440 6 sid_do[15]
port 331 nsew signal input
rlabel metal3 s 0 34944 400 35000 6 sid_do[16]
port 332 nsew signal input
rlabel metal3 s 0 35504 400 35560 6 sid_do[17]
port 333 nsew signal input
rlabel metal3 s 0 36064 400 36120 6 sid_do[18]
port 334 nsew signal input
rlabel metal3 s 0 36624 400 36680 6 sid_do[19]
port 335 nsew signal input
rlabel metal3 s 0 26544 400 26600 6 sid_do[1]
port 336 nsew signal input
rlabel metal3 s 0 37184 400 37240 6 sid_do[20]
port 337 nsew signal input
rlabel metal3 s 0 27104 400 27160 6 sid_do[2]
port 338 nsew signal input
rlabel metal3 s 0 27664 400 27720 6 sid_do[3]
port 339 nsew signal input
rlabel metal3 s 0 28224 400 28280 6 sid_do[4]
port 340 nsew signal input
rlabel metal3 s 0 28784 400 28840 6 sid_do[5]
port 341 nsew signal input
rlabel metal3 s 0 29344 400 29400 6 sid_do[6]
port 342 nsew signal input
rlabel metal3 s 0 29904 400 29960 6 sid_do[7]
port 343 nsew signal input
rlabel metal3 s 0 30464 400 30520 6 sid_do[8]
port 344 nsew signal input
rlabel metal3 s 0 31024 400 31080 6 sid_do[9]
port 345 nsew signal input
rlabel metal3 s 0 37744 400 37800 6 sid_oeb
port 346 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 sn76489_do[0]
port 347 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 sn76489_do[10]
port 348 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 sn76489_do[11]
port 349 nsew signal input
rlabel metal2 s 37520 0 37576 400 6 sn76489_do[12]
port 350 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 sn76489_do[13]
port 351 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 sn76489_do[14]
port 352 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 sn76489_do[15]
port 353 nsew signal input
rlabel metal2 s 39312 0 39368 400 6 sn76489_do[16]
port 354 nsew signal input
rlabel metal2 s 39760 0 39816 400 6 sn76489_do[17]
port 355 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 sn76489_do[18]
port 356 nsew signal input
rlabel metal2 s 40656 0 40712 400 6 sn76489_do[19]
port 357 nsew signal input
rlabel metal2 s 32592 0 32648 400 6 sn76489_do[1]
port 358 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 sn76489_do[20]
port 359 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 sn76489_do[21]
port 360 nsew signal input
rlabel metal2 s 42000 0 42056 400 6 sn76489_do[22]
port 361 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 sn76489_do[23]
port 362 nsew signal input
rlabel metal2 s 42896 0 42952 400 6 sn76489_do[24]
port 363 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 sn76489_do[25]
port 364 nsew signal input
rlabel metal2 s 43792 0 43848 400 6 sn76489_do[26]
port 365 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 sn76489_do[27]
port 366 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 sn76489_do[2]
port 367 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 sn76489_do[3]
port 368 nsew signal input
rlabel metal2 s 33936 0 33992 400 6 sn76489_do[4]
port 369 nsew signal input
rlabel metal2 s 34384 0 34440 400 6 sn76489_do[5]
port 370 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 sn76489_do[6]
port 371 nsew signal input
rlabel metal2 s 35280 0 35336 400 6 sn76489_do[7]
port 372 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 sn76489_do[8]
port 373 nsew signal input
rlabel metal2 s 36176 0 36232 400 6 sn76489_do[9]
port 374 nsew signal input
rlabel metal3 s 0 58464 400 58520 6 tbb1143_do[0]
port 375 nsew signal input
rlabel metal3 s 0 59024 400 59080 6 tbb1143_do[1]
port 376 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 tbb1143_do[2]
port 377 nsew signal input
rlabel metal3 s 0 60144 400 60200 6 tbb1143_do[3]
port 378 nsew signal input
rlabel metal3 s 0 60704 400 60760 6 tbb1143_do[4]
port 379 nsew signal input
rlabel metal4 s 2224 1538 2384 63142 6 vdd
port 380 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 63142 6 vdd
port 380 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 63142 6 vdd
port 380 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 63142 6 vdd
port 380 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 63142 6 vdd
port 380 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 63142 6 vss
port 381 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 63142 6 vss
port 381 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 63142 6 vss
port 381 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 63142 6 vss
port 381 nsew ground bidirectional
rlabel metal2 s 2576 0 2632 400 6 wb_clk_i
port 382 nsew signal input
rlabel metal2 s 3024 0 3080 400 6 wb_rst_i
port 383 nsew signal input
rlabel metal3 s 64600 21840 65000 21896 6 wbs_ack_o
port 384 nsew signal output
rlabel metal2 s 3472 0 3528 400 6 wbs_adr_i[0]
port 385 nsew signal input
rlabel metal2 s 7952 0 8008 400 6 wbs_adr_i[10]
port 386 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 wbs_adr_i[11]
port 387 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_adr_i[12]
port 388 nsew signal input
rlabel metal2 s 9296 0 9352 400 6 wbs_adr_i[13]
port 389 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_adr_i[14]
port 390 nsew signal input
rlabel metal2 s 10192 0 10248 400 6 wbs_adr_i[15]
port 391 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_adr_i[16]
port 392 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_adr_i[17]
port 393 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 wbs_adr_i[18]
port 394 nsew signal input
rlabel metal2 s 11984 0 12040 400 6 wbs_adr_i[19]
port 395 nsew signal input
rlabel metal2 s 3920 0 3976 400 6 wbs_adr_i[1]
port 396 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 wbs_adr_i[20]
port 397 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_adr_i[21]
port 398 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[22]
port 399 nsew signal input
rlabel metal2 s 13776 0 13832 400 6 wbs_adr_i[23]
port 400 nsew signal input
rlabel metal2 s 14224 0 14280 400 6 wbs_adr_i[24]
port 401 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_adr_i[25]
port 402 nsew signal input
rlabel metal2 s 15120 0 15176 400 6 wbs_adr_i[26]
port 403 nsew signal input
rlabel metal2 s 15568 0 15624 400 6 wbs_adr_i[27]
port 404 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 wbs_adr_i[28]
port 405 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 wbs_adr_i[29]
port 406 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_adr_i[2]
port 407 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_adr_i[30]
port 408 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 wbs_adr_i[31]
port 409 nsew signal input
rlabel metal2 s 4816 0 4872 400 6 wbs_adr_i[3]
port 410 nsew signal input
rlabel metal2 s 5264 0 5320 400 6 wbs_adr_i[4]
port 411 nsew signal input
rlabel metal2 s 5712 0 5768 400 6 wbs_adr_i[5]
port 412 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 wbs_adr_i[6]
port 413 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_adr_i[7]
port 414 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 wbs_adr_i[8]
port 415 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 wbs_adr_i[9]
port 416 nsew signal input
rlabel metal3 s 64600 20944 65000 21000 6 wbs_cyc_i
port 417 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[0]
port 418 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[10]
port 419 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 wbs_dat_i[11]
port 420 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 wbs_dat_i[12]
port 421 nsew signal input
rlabel metal2 s 23632 0 23688 400 6 wbs_dat_i[13]
port 422 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 wbs_dat_i[14]
port 423 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 wbs_dat_i[15]
port 424 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 wbs_dat_i[16]
port 425 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 wbs_dat_i[17]
port 426 nsew signal input
rlabel metal2 s 25872 0 25928 400 6 wbs_dat_i[18]
port 427 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 wbs_dat_i[19]
port 428 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 wbs_dat_i[1]
port 429 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_dat_i[20]
port 430 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 wbs_dat_i[21]
port 431 nsew signal input
rlabel metal2 s 27664 0 27720 400 6 wbs_dat_i[22]
port 432 nsew signal input
rlabel metal2 s 28112 0 28168 400 6 wbs_dat_i[23]
port 433 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 wbs_dat_i[24]
port 434 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 wbs_dat_i[25]
port 435 nsew signal input
rlabel metal2 s 29456 0 29512 400 6 wbs_dat_i[26]
port 436 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 wbs_dat_i[27]
port 437 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 wbs_dat_i[28]
port 438 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 wbs_dat_i[29]
port 439 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 wbs_dat_i[2]
port 440 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 wbs_dat_i[30]
port 441 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 wbs_dat_i[31]
port 442 nsew signal input
rlabel metal2 s 19152 0 19208 400 6 wbs_dat_i[3]
port 443 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_i[4]
port 444 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_dat_i[5]
port 445 nsew signal input
rlabel metal2 s 20496 0 20552 400 6 wbs_dat_i[6]
port 446 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_dat_i[7]
port 447 nsew signal input
rlabel metal2 s 21392 0 21448 400 6 wbs_dat_i[8]
port 448 nsew signal input
rlabel metal2 s 21840 0 21896 400 6 wbs_dat_i[9]
port 449 nsew signal input
rlabel metal3 s 64600 6160 65000 6216 6 wbs_dat_o[0]
port 450 nsew signal output
rlabel metal3 s 64600 10640 65000 10696 6 wbs_dat_o[10]
port 451 nsew signal output
rlabel metal3 s 64600 11088 65000 11144 6 wbs_dat_o[11]
port 452 nsew signal output
rlabel metal3 s 64600 11536 65000 11592 6 wbs_dat_o[12]
port 453 nsew signal output
rlabel metal3 s 64600 11984 65000 12040 6 wbs_dat_o[13]
port 454 nsew signal output
rlabel metal3 s 64600 12432 65000 12488 6 wbs_dat_o[14]
port 455 nsew signal output
rlabel metal3 s 64600 12880 65000 12936 6 wbs_dat_o[15]
port 456 nsew signal output
rlabel metal3 s 64600 13328 65000 13384 6 wbs_dat_o[16]
port 457 nsew signal output
rlabel metal3 s 64600 13776 65000 13832 6 wbs_dat_o[17]
port 458 nsew signal output
rlabel metal3 s 64600 14224 65000 14280 6 wbs_dat_o[18]
port 459 nsew signal output
rlabel metal3 s 64600 14672 65000 14728 6 wbs_dat_o[19]
port 460 nsew signal output
rlabel metal3 s 64600 6608 65000 6664 6 wbs_dat_o[1]
port 461 nsew signal output
rlabel metal3 s 64600 15120 65000 15176 6 wbs_dat_o[20]
port 462 nsew signal output
rlabel metal3 s 64600 15568 65000 15624 6 wbs_dat_o[21]
port 463 nsew signal output
rlabel metal3 s 64600 16016 65000 16072 6 wbs_dat_o[22]
port 464 nsew signal output
rlabel metal3 s 64600 16464 65000 16520 6 wbs_dat_o[23]
port 465 nsew signal output
rlabel metal3 s 64600 16912 65000 16968 6 wbs_dat_o[24]
port 466 nsew signal output
rlabel metal3 s 64600 17360 65000 17416 6 wbs_dat_o[25]
port 467 nsew signal output
rlabel metal3 s 64600 17808 65000 17864 6 wbs_dat_o[26]
port 468 nsew signal output
rlabel metal3 s 64600 18256 65000 18312 6 wbs_dat_o[27]
port 469 nsew signal output
rlabel metal3 s 64600 18704 65000 18760 6 wbs_dat_o[28]
port 470 nsew signal output
rlabel metal3 s 64600 19152 65000 19208 6 wbs_dat_o[29]
port 471 nsew signal output
rlabel metal3 s 64600 7056 65000 7112 6 wbs_dat_o[2]
port 472 nsew signal output
rlabel metal3 s 64600 19600 65000 19656 6 wbs_dat_o[30]
port 473 nsew signal output
rlabel metal3 s 64600 20048 65000 20104 6 wbs_dat_o[31]
port 474 nsew signal output
rlabel metal3 s 64600 7504 65000 7560 6 wbs_dat_o[3]
port 475 nsew signal output
rlabel metal3 s 64600 7952 65000 8008 6 wbs_dat_o[4]
port 476 nsew signal output
rlabel metal3 s 64600 8400 65000 8456 6 wbs_dat_o[5]
port 477 nsew signal output
rlabel metal3 s 64600 8848 65000 8904 6 wbs_dat_o[6]
port 478 nsew signal output
rlabel metal3 s 64600 9296 65000 9352 6 wbs_dat_o[7]
port 479 nsew signal output
rlabel metal3 s 64600 9744 65000 9800 6 wbs_dat_o[8]
port 480 nsew signal output
rlabel metal3 s 64600 10192 65000 10248 6 wbs_dat_o[9]
port 481 nsew signal output
rlabel metal3 s 64600 21392 65000 21448 6 wbs_stb_i
port 482 nsew signal input
rlabel metal3 s 64600 20496 65000 20552 6 wbs_we_i
port 483 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 65000 65000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8777358
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/Multiplexer/runs/23_11_15_15_44/results/signoff/multiplexer.magic.gds
string GDS_START 387912
<< end >>

