VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ay8913
  CLASS BLOCK ;
  FOREIGN wrapped_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 255.000 BY 255.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 180.320 255.000 180.880 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 201.600 255.000 202.160 ;
    END
  END custom_settings[1]
  PIN custom_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 222.880 255.000 223.440 ;
    END
  END custom_settings[2]
  PIN custom_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 244.160 255.000 244.720 ;
    END
  END custom_settings[3]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 10.080 255.000 10.640 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 31.360 255.000 31.920 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 52.640 255.000 53.200 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 73.920 255.000 74.480 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 95.200 255.000 95.760 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 116.480 255.000 117.040 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 137.760 255.000 138.320 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 251.000 159.040 255.000 159.600 ;
    END
  END io_in_1[7]
  PIN io_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 251.000 159.600 255.000 ;
    END
  END io_in_2[0]
  PIN io_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 222.880 251.000 223.440 255.000 ;
    END
  END io_in_2[1]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 0.000 15.120 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 251.000 95.760 255.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 239.420 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 239.420 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 239.420 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 251.000 31.920 255.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 248.080 240.090 ;
      LAYER Metal2 ;
        RECT 5.740 250.700 31.060 251.000 ;
        RECT 32.220 250.700 94.900 251.000 ;
        RECT 96.060 250.700 158.740 251.000 ;
        RECT 159.900 250.700 222.580 251.000 ;
        RECT 223.740 250.700 248.500 251.000 ;
        RECT 5.740 4.300 248.500 250.700 ;
        RECT 6.460 3.500 14.260 4.300 ;
        RECT 15.420 3.500 23.220 4.300 ;
        RECT 24.380 3.500 32.180 4.300 ;
        RECT 33.340 3.500 41.140 4.300 ;
        RECT 42.300 3.500 50.100 4.300 ;
        RECT 51.260 3.500 59.060 4.300 ;
        RECT 60.220 3.500 68.020 4.300 ;
        RECT 69.180 3.500 76.980 4.300 ;
        RECT 78.140 3.500 85.940 4.300 ;
        RECT 87.100 3.500 94.900 4.300 ;
        RECT 96.060 3.500 103.860 4.300 ;
        RECT 105.020 3.500 112.820 4.300 ;
        RECT 113.980 3.500 121.780 4.300 ;
        RECT 122.940 3.500 130.740 4.300 ;
        RECT 131.900 3.500 139.700 4.300 ;
        RECT 140.860 3.500 148.660 4.300 ;
        RECT 149.820 3.500 157.620 4.300 ;
        RECT 158.780 3.500 166.580 4.300 ;
        RECT 167.740 3.500 175.540 4.300 ;
        RECT 176.700 3.500 184.500 4.300 ;
        RECT 185.660 3.500 193.460 4.300 ;
        RECT 194.620 3.500 202.420 4.300 ;
        RECT 203.580 3.500 211.380 4.300 ;
        RECT 212.540 3.500 220.340 4.300 ;
        RECT 221.500 3.500 229.300 4.300 ;
        RECT 230.460 3.500 238.260 4.300 ;
        RECT 239.420 3.500 247.220 4.300 ;
        RECT 248.380 3.500 248.500 4.300 ;
      LAYER Metal3 ;
        RECT 8.490 243.860 250.700 244.580 ;
        RECT 8.490 223.740 251.000 243.860 ;
        RECT 8.490 222.580 250.700 223.740 ;
        RECT 8.490 202.460 251.000 222.580 ;
        RECT 8.490 201.300 250.700 202.460 ;
        RECT 8.490 181.180 251.000 201.300 ;
        RECT 8.490 180.020 250.700 181.180 ;
        RECT 8.490 159.900 251.000 180.020 ;
        RECT 8.490 158.740 250.700 159.900 ;
        RECT 8.490 138.620 251.000 158.740 ;
        RECT 8.490 137.460 250.700 138.620 ;
        RECT 8.490 117.340 251.000 137.460 ;
        RECT 8.490 116.180 250.700 117.340 ;
        RECT 8.490 96.060 251.000 116.180 ;
        RECT 8.490 94.900 250.700 96.060 ;
        RECT 8.490 74.780 251.000 94.900 ;
        RECT 8.490 73.620 250.700 74.780 ;
        RECT 8.490 53.500 251.000 73.620 ;
        RECT 8.490 52.340 250.700 53.500 ;
        RECT 8.490 32.220 251.000 52.340 ;
        RECT 8.490 31.060 250.700 32.220 ;
        RECT 8.490 10.940 251.000 31.060 ;
        RECT 8.490 10.220 250.700 10.940 ;
      LAYER Metal4 ;
        RECT 16.940 16.890 21.940 235.110 ;
        RECT 24.140 16.890 98.740 235.110 ;
        RECT 100.940 16.890 175.540 235.110 ;
        RECT 177.740 16.890 241.220 235.110 ;
  END
END wrapped_ay8913
END LIBRARY

